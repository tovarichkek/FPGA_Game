module logo_rom (
  input  wire    [16:0]     addr,
  output wire    [11:0]     word
);
  logic [11:0] rom [(400 * 320)];
  assign word = rom[addr];
  initial begin
rom[0] = 12'h444;
rom[1] = 12'h444;
rom[2] = 12'h444;
rom[3] = 12'h444;
rom[4] = 12'h444;
rom[5] = 12'h444;
rom[6] = 12'h444;
rom[7] = 12'h444;
rom[8] = 12'h444;
rom[9] = 12'h444;
rom[10] = 12'h444;
rom[11] = 12'h444;
rom[12] = 12'h444;
rom[13] = 12'h444;
rom[14] = 12'h444;
rom[15] = 12'h444;
rom[16] = 12'h444;
rom[17] = 12'h555;
rom[18] = 12'h555;
rom[19] = 12'h555;
rom[20] = 12'h555;
rom[21] = 12'h555;
rom[22] = 12'h555;
rom[23] = 12'h555;
rom[24] = 12'h555;
rom[25] = 12'h555;
rom[26] = 12'h555;
rom[27] = 12'h666;
rom[28] = 12'h666;
rom[29] = 12'h666;
rom[30] = 12'h666;
rom[31] = 12'h666;
rom[32] = 12'h666;
rom[33] = 12'h666;
rom[34] = 12'h777;
rom[35] = 12'h777;
rom[36] = 12'h777;
rom[37] = 12'h777;
rom[38] = 12'h777;
rom[39] = 12'h777;
rom[40] = 12'h777;
rom[41] = 12'h777;
rom[42] = 12'h666;
rom[43] = 12'h666;
rom[44] = 12'h666;
rom[45] = 12'h555;
rom[46] = 12'h555;
rom[47] = 12'h555;
rom[48] = 12'h555;
rom[49] = 12'h555;
rom[50] = 12'h555;
rom[51] = 12'h555;
rom[52] = 12'h555;
rom[53] = 12'h555;
rom[54] = 12'h555;
rom[55] = 12'h555;
rom[56] = 12'h555;
rom[57] = 12'h555;
rom[58] = 12'h555;
rom[59] = 12'h666;
rom[60] = 12'h666;
rom[61] = 12'h666;
rom[62] = 12'h666;
rom[63] = 12'h666;
rom[64] = 12'h666;
rom[65] = 12'h666;
rom[66] = 12'h666;
rom[67] = 12'h666;
rom[68] = 12'h777;
rom[69] = 12'h777;
rom[70] = 12'h777;
rom[71] = 12'h777;
rom[72] = 12'h777;
rom[73] = 12'h777;
rom[74] = 12'h777;
rom[75] = 12'h777;
rom[76] = 12'h777;
rom[77] = 12'h666;
rom[78] = 12'h666;
rom[79] = 12'h666;
rom[80] = 12'h666;
rom[81] = 12'h666;
rom[82] = 12'h555;
rom[83] = 12'h555;
rom[84] = 12'h555;
rom[85] = 12'h555;
rom[86] = 12'h555;
rom[87] = 12'h555;
rom[88] = 12'h555;
rom[89] = 12'h555;
rom[90] = 12'h555;
rom[91] = 12'h555;
rom[92] = 12'h555;
rom[93] = 12'h555;
rom[94] = 12'h555;
rom[95] = 12'h666;
rom[96] = 12'h666;
rom[97] = 12'h666;
rom[98] = 12'h666;
rom[99] = 12'h777;
rom[100] = 12'h888;
rom[101] = 12'h888;
rom[102] = 12'h888;
rom[103] = 12'h888;
rom[104] = 12'h999;
rom[105] = 12'h999;
rom[106] = 12'h999;
rom[107] = 12'h999;
rom[108] = 12'h999;
rom[109] = 12'h999;
rom[110] = 12'h999;
rom[111] = 12'h999;
rom[112] = 12'h999;
rom[113] = 12'h999;
rom[114] = 12'h999;
rom[115] = 12'ha99;
rom[116] = 12'haaa;
rom[117] = 12'haaa;
rom[118] = 12'hbaa;
rom[119] = 12'hbaa;
rom[120] = 12'hbab;
rom[121] = 12'hbab;
rom[122] = 12'hbaa;
rom[123] = 12'hbaa;
rom[124] = 12'hbaa;
rom[125] = 12'hbaa;
rom[126] = 12'hbaa;
rom[127] = 12'hbaa;
rom[128] = 12'haaa;
rom[129] = 12'haaa;
rom[130] = 12'haaa;
rom[131] = 12'h9aa;
rom[132] = 12'h9aa;
rom[133] = 12'h9aa;
rom[134] = 12'h9aa;
rom[135] = 12'h9aa;
rom[136] = 12'h9aa;
rom[137] = 12'h9aa;
rom[138] = 12'h9aa;
rom[139] = 12'h9a9;
rom[140] = 12'h999;
rom[141] = 12'h999;
rom[142] = 12'h888;
rom[143] = 12'h888;
rom[144] = 12'h787;
rom[145] = 12'h787;
rom[146] = 12'h787;
rom[147] = 12'h777;
rom[148] = 12'h777;
rom[149] = 12'h676;
rom[150] = 12'h676;
rom[151] = 12'h666;
rom[152] = 12'h566;
rom[153] = 12'h565;
rom[154] = 12'h565;
rom[155] = 12'h565;
rom[156] = 12'h565;
rom[157] = 12'h565;
rom[158] = 12'h565;
rom[159] = 12'h566;
rom[160] = 12'h556;
rom[161] = 12'h555;
rom[162] = 12'h555;
rom[163] = 12'h555;
rom[164] = 12'h445;
rom[165] = 12'h444;
rom[166] = 12'h444;
rom[167] = 12'h444;
rom[168] = 12'h334;
rom[169] = 12'h333;
rom[170] = 12'h333;
rom[171] = 12'h333;
rom[172] = 12'h334;
rom[173] = 12'h333;
rom[174] = 12'h333;
rom[175] = 12'h222;
rom[176] = 12'h222;
rom[177] = 12'h222;
rom[178] = 12'h222;
rom[179] = 12'h333;
rom[180] = 12'h333;
rom[181] = 12'h444;
rom[182] = 12'h444;
rom[183] = 12'h333;
rom[184] = 12'h444;
rom[185] = 12'h444;
rom[186] = 12'h444;
rom[187] = 12'h444;
rom[188] = 12'h333;
rom[189] = 12'h333;
rom[190] = 12'h333;
rom[191] = 12'h444;
rom[192] = 12'h444;
rom[193] = 12'h444;
rom[194] = 12'h555;
rom[195] = 12'h666;
rom[196] = 12'h777;
rom[197] = 12'h666;
rom[198] = 12'h666;
rom[199] = 12'h777;
rom[200] = 12'h555;
rom[201] = 12'h444;
rom[202] = 12'h333;
rom[203] = 12'h444;
rom[204] = 12'h444;
rom[205] = 12'h444;
rom[206] = 12'h444;
rom[207] = 12'h333;
rom[208] = 12'h222;
rom[209] = 12'h111;
rom[210] = 12'h  0;
rom[211] = 12'h111;
rom[212] = 12'h111;
rom[213] = 12'h  0;
rom[214] = 12'h  0;
rom[215] = 12'h  0;
rom[216] = 12'h  0;
rom[217] = 12'h  0;
rom[218] = 12'h111;
rom[219] = 12'h222;
rom[220] = 12'h222;
rom[221] = 12'h  0;
rom[222] = 12'h  0;
rom[223] = 12'h  0;
rom[224] = 12'h  0;
rom[225] = 12'h  0;
rom[226] = 12'h  0;
rom[227] = 12'h  0;
rom[228] = 12'h  0;
rom[229] = 12'h  0;
rom[230] = 12'h  0;
rom[231] = 12'h  0;
rom[232] = 12'h  0;
rom[233] = 12'h  0;
rom[234] = 12'h  0;
rom[235] = 12'h  0;
rom[236] = 12'h  0;
rom[237] = 12'h  0;
rom[238] = 12'h  0;
rom[239] = 12'h  0;
rom[240] = 12'h  0;
rom[241] = 12'h  0;
rom[242] = 12'h  0;
rom[243] = 12'h  0;
rom[244] = 12'h  0;
rom[245] = 12'h  0;
rom[246] = 12'h  0;
rom[247] = 12'h  0;
rom[248] = 12'h  0;
rom[249] = 12'h  0;
rom[250] = 12'h  0;
rom[251] = 12'h  0;
rom[252] = 12'h  0;
rom[253] = 12'h  0;
rom[254] = 12'h  0;
rom[255] = 12'h  0;
rom[256] = 12'h  0;
rom[257] = 12'h  0;
rom[258] = 12'h111;
rom[259] = 12'h  0;
rom[260] = 12'h  0;
rom[261] = 12'h222;
rom[262] = 12'h333;
rom[263] = 12'h333;
rom[264] = 12'h333;
rom[265] = 12'h222;
rom[266] = 12'h111;
rom[267] = 12'h  0;
rom[268] = 12'h  0;
rom[269] = 12'h  0;
rom[270] = 12'h  0;
rom[271] = 12'h  0;
rom[272] = 12'h  0;
rom[273] = 12'h  0;
rom[274] = 12'h  0;
rom[275] = 12'h  0;
rom[276] = 12'h  0;
rom[277] = 12'h  0;
rom[278] = 12'h  0;
rom[279] = 12'h  0;
rom[280] = 12'h  0;
rom[281] = 12'h  0;
rom[282] = 12'h  0;
rom[283] = 12'h  0;
rom[284] = 12'h  0;
rom[285] = 12'h  0;
rom[286] = 12'h  0;
rom[287] = 12'h  0;
rom[288] = 12'h  0;
rom[289] = 12'h  0;
rom[290] = 12'h  0;
rom[291] = 12'h  0;
rom[292] = 12'h  0;
rom[293] = 12'h  0;
rom[294] = 12'h  0;
rom[295] = 12'h  0;
rom[296] = 12'h  0;
rom[297] = 12'h  0;
rom[298] = 12'h  0;
rom[299] = 12'h  0;
rom[300] = 12'h111;
rom[301] = 12'h111;
rom[302] = 12'h111;
rom[303] = 12'h  0;
rom[304] = 12'h  0;
rom[305] = 12'h  0;
rom[306] = 12'h  0;
rom[307] = 12'h  0;
rom[308] = 12'h  0;
rom[309] = 12'h  0;
rom[310] = 12'h  0;
rom[311] = 12'h  0;
rom[312] = 12'h  0;
rom[313] = 12'h  0;
rom[314] = 12'h  0;
rom[315] = 12'h  0;
rom[316] = 12'h  0;
rom[317] = 12'h  0;
rom[318] = 12'h  0;
rom[319] = 12'h  0;
rom[320] = 12'h  0;
rom[321] = 12'h111;
rom[322] = 12'h222;
rom[323] = 12'h444;
rom[324] = 12'h555;
rom[325] = 12'h555;
rom[326] = 12'h444;
rom[327] = 12'h333;
rom[328] = 12'h222;
rom[329] = 12'h222;
rom[330] = 12'h111;
rom[331] = 12'h111;
rom[332] = 12'h111;
rom[333] = 12'h111;
rom[334] = 12'h111;
rom[335] = 12'h111;
rom[336] = 12'h111;
rom[337] = 12'h111;
rom[338] = 12'h111;
rom[339] = 12'h111;
rom[340] = 12'h111;
rom[341] = 12'h111;
rom[342] = 12'h222;
rom[343] = 12'h222;
rom[344] = 12'h222;
rom[345] = 12'h222;
rom[346] = 12'h222;
rom[347] = 12'h222;
rom[348] = 12'h222;
rom[349] = 12'h333;
rom[350] = 12'h333;
rom[351] = 12'h333;
rom[352] = 12'h333;
rom[353] = 12'h333;
rom[354] = 12'h333;
rom[355] = 12'h444;
rom[356] = 12'h666;
rom[357] = 12'h777;
rom[358] = 12'h666;
rom[359] = 12'h555;
rom[360] = 12'h555;
rom[361] = 12'h555;
rom[362] = 12'h555;
rom[363] = 12'h444;
rom[364] = 12'h444;
rom[365] = 12'h444;
rom[366] = 12'h444;
rom[367] = 12'h444;
rom[368] = 12'h555;
rom[369] = 12'h555;
rom[370] = 12'h555;
rom[371] = 12'h555;
rom[372] = 12'h444;
rom[373] = 12'h555;
rom[374] = 12'h555;
rom[375] = 12'h666;
rom[376] = 12'h777;
rom[377] = 12'h777;
rom[378] = 12'h777;
rom[379] = 12'h777;
rom[380] = 12'h999;
rom[381] = 12'haaa;
rom[382] = 12'hbbb;
rom[383] = 12'hccc;
rom[384] = 12'h999;
rom[385] = 12'h999;
rom[386] = 12'h999;
rom[387] = 12'h999;
rom[388] = 12'h999;
rom[389] = 12'h999;
rom[390] = 12'haaa;
rom[391] = 12'haaa;
rom[392] = 12'haaa;
rom[393] = 12'haaa;
rom[394] = 12'haaa;
rom[395] = 12'h999;
rom[396] = 12'h999;
rom[397] = 12'h999;
rom[398] = 12'h999;
rom[399] = 12'h999;
rom[400] = 12'h444;
rom[401] = 12'h444;
rom[402] = 12'h444;
rom[403] = 12'h444;
rom[404] = 12'h444;
rom[405] = 12'h444;
rom[406] = 12'h444;
rom[407] = 12'h444;
rom[408] = 12'h444;
rom[409] = 12'h444;
rom[410] = 12'h444;
rom[411] = 12'h444;
rom[412] = 12'h444;
rom[413] = 12'h444;
rom[414] = 12'h444;
rom[415] = 12'h444;
rom[416] = 12'h444;
rom[417] = 12'h444;
rom[418] = 12'h555;
rom[419] = 12'h555;
rom[420] = 12'h555;
rom[421] = 12'h555;
rom[422] = 12'h555;
rom[423] = 12'h555;
rom[424] = 12'h555;
rom[425] = 12'h555;
rom[426] = 12'h555;
rom[427] = 12'h666;
rom[428] = 12'h666;
rom[429] = 12'h666;
rom[430] = 12'h666;
rom[431] = 12'h666;
rom[432] = 12'h666;
rom[433] = 12'h666;
rom[434] = 12'h666;
rom[435] = 12'h666;
rom[436] = 12'h666;
rom[437] = 12'h666;
rom[438] = 12'h666;
rom[439] = 12'h666;
rom[440] = 12'h666;
rom[441] = 12'h666;
rom[442] = 12'h666;
rom[443] = 12'h555;
rom[444] = 12'h555;
rom[445] = 12'h555;
rom[446] = 12'h555;
rom[447] = 12'h444;
rom[448] = 12'h555;
rom[449] = 12'h555;
rom[450] = 12'h555;
rom[451] = 12'h555;
rom[452] = 12'h555;
rom[453] = 12'h555;
rom[454] = 12'h555;
rom[455] = 12'h555;
rom[456] = 12'h555;
rom[457] = 12'h555;
rom[458] = 12'h555;
rom[459] = 12'h555;
rom[460] = 12'h555;
rom[461] = 12'h555;
rom[462] = 12'h555;
rom[463] = 12'h666;
rom[464] = 12'h555;
rom[465] = 12'h555;
rom[466] = 12'h666;
rom[467] = 12'h666;
rom[468] = 12'h666;
rom[469] = 12'h666;
rom[470] = 12'h666;
rom[471] = 12'h666;
rom[472] = 12'h777;
rom[473] = 12'h777;
rom[474] = 12'h777;
rom[475] = 12'h666;
rom[476] = 12'h666;
rom[477] = 12'h666;
rom[478] = 12'h666;
rom[479] = 12'h666;
rom[480] = 12'h666;
rom[481] = 12'h666;
rom[482] = 12'h666;
rom[483] = 12'h666;
rom[484] = 12'h666;
rom[485] = 12'h666;
rom[486] = 12'h666;
rom[487] = 12'h555;
rom[488] = 12'h555;
rom[489] = 12'h666;
rom[490] = 12'h666;
rom[491] = 12'h666;
rom[492] = 12'h666;
rom[493] = 12'h666;
rom[494] = 12'h666;
rom[495] = 12'h666;
rom[496] = 12'h666;
rom[497] = 12'h666;
rom[498] = 12'h777;
rom[499] = 12'h777;
rom[500] = 12'h777;
rom[501] = 12'h888;
rom[502] = 12'h888;
rom[503] = 12'h888;
rom[504] = 12'h888;
rom[505] = 12'h888;
rom[506] = 12'h888;
rom[507] = 12'h888;
rom[508] = 12'h888;
rom[509] = 12'h999;
rom[510] = 12'h999;
rom[511] = 12'h999;
rom[512] = 12'h999;
rom[513] = 12'h999;
rom[514] = 12'h999;
rom[515] = 12'h999;
rom[516] = 12'h999;
rom[517] = 12'ha9a;
rom[518] = 12'ha9a;
rom[519] = 12'ha9a;
rom[520] = 12'ha9a;
rom[521] = 12'ha9a;
rom[522] = 12'hbaa;
rom[523] = 12'hbaa;
rom[524] = 12'hbaa;
rom[525] = 12'hbaa;
rom[526] = 12'hcaa;
rom[527] = 12'hbba;
rom[528] = 12'haaa;
rom[529] = 12'haaa;
rom[530] = 12'haaa;
rom[531] = 12'h9aa;
rom[532] = 12'h9aa;
rom[533] = 12'h9aa;
rom[534] = 12'h9aa;
rom[535] = 12'haaa;
rom[536] = 12'h9aa;
rom[537] = 12'h9aa;
rom[538] = 12'h9a9;
rom[539] = 12'h999;
rom[540] = 12'h999;
rom[541] = 12'h999;
rom[542] = 12'h888;
rom[543] = 12'h888;
rom[544] = 12'h887;
rom[545] = 12'h787;
rom[546] = 12'h777;
rom[547] = 12'h777;
rom[548] = 12'h777;
rom[549] = 12'h776;
rom[550] = 12'h676;
rom[551] = 12'h676;
rom[552] = 12'h666;
rom[553] = 12'h666;
rom[554] = 12'h566;
rom[555] = 12'h565;
rom[556] = 12'h565;
rom[557] = 12'h565;
rom[558] = 12'h565;
rom[559] = 12'h565;
rom[560] = 12'h555;
rom[561] = 12'h555;
rom[562] = 12'h555;
rom[563] = 12'h555;
rom[564] = 12'h445;
rom[565] = 12'h444;
rom[566] = 12'h444;
rom[567] = 12'h444;
rom[568] = 12'h333;
rom[569] = 12'h333;
rom[570] = 12'h333;
rom[571] = 12'h333;
rom[572] = 12'h334;
rom[573] = 12'h333;
rom[574] = 12'h333;
rom[575] = 12'h323;
rom[576] = 12'h222;
rom[577] = 12'h222;
rom[578] = 12'h222;
rom[579] = 12'h333;
rom[580] = 12'h333;
rom[581] = 12'h333;
rom[582] = 12'h444;
rom[583] = 12'h333;
rom[584] = 12'h444;
rom[585] = 12'h444;
rom[586] = 12'h444;
rom[587] = 12'h444;
rom[588] = 12'h444;
rom[589] = 12'h333;
rom[590] = 12'h333;
rom[591] = 12'h444;
rom[592] = 12'h444;
rom[593] = 12'h444;
rom[594] = 12'h555;
rom[595] = 12'h666;
rom[596] = 12'h777;
rom[597] = 12'h666;
rom[598] = 12'h666;
rom[599] = 12'h777;
rom[600] = 12'h555;
rom[601] = 12'h444;
rom[602] = 12'h444;
rom[603] = 12'h444;
rom[604] = 12'h444;
rom[605] = 12'h444;
rom[606] = 12'h444;
rom[607] = 12'h333;
rom[608] = 12'h222;
rom[609] = 12'h111;
rom[610] = 12'h  0;
rom[611] = 12'h111;
rom[612] = 12'h111;
rom[613] = 12'h  0;
rom[614] = 12'h  0;
rom[615] = 12'h  0;
rom[616] = 12'h  0;
rom[617] = 12'h  0;
rom[618] = 12'h111;
rom[619] = 12'h222;
rom[620] = 12'h222;
rom[621] = 12'h  0;
rom[622] = 12'h  0;
rom[623] = 12'h  0;
rom[624] = 12'h  0;
rom[625] = 12'h  0;
rom[626] = 12'h  0;
rom[627] = 12'h  0;
rom[628] = 12'h  0;
rom[629] = 12'h  0;
rom[630] = 12'h  0;
rom[631] = 12'h  0;
rom[632] = 12'h  0;
rom[633] = 12'h  0;
rom[634] = 12'h  0;
rom[635] = 12'h  0;
rom[636] = 12'h  0;
rom[637] = 12'h  0;
rom[638] = 12'h  0;
rom[639] = 12'h  0;
rom[640] = 12'h  0;
rom[641] = 12'h  0;
rom[642] = 12'h  0;
rom[643] = 12'h  0;
rom[644] = 12'h  0;
rom[645] = 12'h  0;
rom[646] = 12'h  0;
rom[647] = 12'h  0;
rom[648] = 12'h  0;
rom[649] = 12'h  0;
rom[650] = 12'h  0;
rom[651] = 12'h  0;
rom[652] = 12'h  0;
rom[653] = 12'h  0;
rom[654] = 12'h  0;
rom[655] = 12'h111;
rom[656] = 12'h  0;
rom[657] = 12'h111;
rom[658] = 12'h  0;
rom[659] = 12'h  0;
rom[660] = 12'h  0;
rom[661] = 12'h222;
rom[662] = 12'h333;
rom[663] = 12'h333;
rom[664] = 12'h333;
rom[665] = 12'h222;
rom[666] = 12'h111;
rom[667] = 12'h  0;
rom[668] = 12'h  0;
rom[669] = 12'h  0;
rom[670] = 12'h  0;
rom[671] = 12'h  0;
rom[672] = 12'h  0;
rom[673] = 12'h  0;
rom[674] = 12'h  0;
rom[675] = 12'h  0;
rom[676] = 12'h  0;
rom[677] = 12'h  0;
rom[678] = 12'h  0;
rom[679] = 12'h  0;
rom[680] = 12'h  0;
rom[681] = 12'h  0;
rom[682] = 12'h  0;
rom[683] = 12'h  0;
rom[684] = 12'h  0;
rom[685] = 12'h  0;
rom[686] = 12'h  0;
rom[687] = 12'h  0;
rom[688] = 12'h  0;
rom[689] = 12'h  0;
rom[690] = 12'h  0;
rom[691] = 12'h  0;
rom[692] = 12'h  0;
rom[693] = 12'h  0;
rom[694] = 12'h  0;
rom[695] = 12'h  0;
rom[696] = 12'h  0;
rom[697] = 12'h  0;
rom[698] = 12'h  0;
rom[699] = 12'h  0;
rom[700] = 12'h111;
rom[701] = 12'h111;
rom[702] = 12'h111;
rom[703] = 12'h  0;
rom[704] = 12'h  0;
rom[705] = 12'h  0;
rom[706] = 12'h  0;
rom[707] = 12'h  0;
rom[708] = 12'h  0;
rom[709] = 12'h  0;
rom[710] = 12'h  0;
rom[711] = 12'h  0;
rom[712] = 12'h  0;
rom[713] = 12'h  0;
rom[714] = 12'h  0;
rom[715] = 12'h  0;
rom[716] = 12'h  0;
rom[717] = 12'h  0;
rom[718] = 12'h  0;
rom[719] = 12'h  0;
rom[720] = 12'h111;
rom[721] = 12'h111;
rom[722] = 12'h222;
rom[723] = 12'h444;
rom[724] = 12'h555;
rom[725] = 12'h555;
rom[726] = 12'h444;
rom[727] = 12'h333;
rom[728] = 12'h222;
rom[729] = 12'h111;
rom[730] = 12'h111;
rom[731] = 12'h111;
rom[732] = 12'h111;
rom[733] = 12'h111;
rom[734] = 12'h111;
rom[735] = 12'h111;
rom[736] = 12'h111;
rom[737] = 12'h111;
rom[738] = 12'h111;
rom[739] = 12'h111;
rom[740] = 12'h111;
rom[741] = 12'h111;
rom[742] = 12'h222;
rom[743] = 12'h222;
rom[744] = 12'h222;
rom[745] = 12'h222;
rom[746] = 12'h222;
rom[747] = 12'h222;
rom[748] = 12'h333;
rom[749] = 12'h333;
rom[750] = 12'h333;
rom[751] = 12'h333;
rom[752] = 12'h333;
rom[753] = 12'h333;
rom[754] = 12'h333;
rom[755] = 12'h555;
rom[756] = 12'h666;
rom[757] = 12'h777;
rom[758] = 12'h666;
rom[759] = 12'h555;
rom[760] = 12'h555;
rom[761] = 12'h555;
rom[762] = 12'h555;
rom[763] = 12'h555;
rom[764] = 12'h555;
rom[765] = 12'h555;
rom[766] = 12'h555;
rom[767] = 12'h555;
rom[768] = 12'h555;
rom[769] = 12'h555;
rom[770] = 12'h555;
rom[771] = 12'h555;
rom[772] = 12'h666;
rom[773] = 12'h666;
rom[774] = 12'h666;
rom[775] = 12'h666;
rom[776] = 12'h666;
rom[777] = 12'h777;
rom[778] = 12'h888;
rom[779] = 12'h999;
rom[780] = 12'haaa;
rom[781] = 12'haaa;
rom[782] = 12'haaa;
rom[783] = 12'haaa;
rom[784] = 12'h999;
rom[785] = 12'h999;
rom[786] = 12'h888;
rom[787] = 12'h888;
rom[788] = 12'h999;
rom[789] = 12'h999;
rom[790] = 12'haaa;
rom[791] = 12'haaa;
rom[792] = 12'haaa;
rom[793] = 12'haaa;
rom[794] = 12'h999;
rom[795] = 12'h999;
rom[796] = 12'h999;
rom[797] = 12'h999;
rom[798] = 12'h999;
rom[799] = 12'h999;
rom[800] = 12'h444;
rom[801] = 12'h444;
rom[802] = 12'h444;
rom[803] = 12'h444;
rom[804] = 12'h444;
rom[805] = 12'h444;
rom[806] = 12'h444;
rom[807] = 12'h444;
rom[808] = 12'h444;
rom[809] = 12'h444;
rom[810] = 12'h444;
rom[811] = 12'h444;
rom[812] = 12'h444;
rom[813] = 12'h444;
rom[814] = 12'h444;
rom[815] = 12'h444;
rom[816] = 12'h444;
rom[817] = 12'h444;
rom[818] = 12'h444;
rom[819] = 12'h555;
rom[820] = 12'h555;
rom[821] = 12'h555;
rom[822] = 12'h555;
rom[823] = 12'h555;
rom[824] = 12'h555;
rom[825] = 12'h555;
rom[826] = 12'h555;
rom[827] = 12'h555;
rom[828] = 12'h666;
rom[829] = 12'h666;
rom[830] = 12'h666;
rom[831] = 12'h555;
rom[832] = 12'h666;
rom[833] = 12'h666;
rom[834] = 12'h666;
rom[835] = 12'h555;
rom[836] = 12'h555;
rom[837] = 12'h555;
rom[838] = 12'h555;
rom[839] = 12'h555;
rom[840] = 12'h555;
rom[841] = 12'h555;
rom[842] = 12'h555;
rom[843] = 12'h444;
rom[844] = 12'h444;
rom[845] = 12'h444;
rom[846] = 12'h444;
rom[847] = 12'h444;
rom[848] = 12'h444;
rom[849] = 12'h444;
rom[850] = 12'h444;
rom[851] = 12'h444;
rom[852] = 12'h444;
rom[853] = 12'h444;
rom[854] = 12'h444;
rom[855] = 12'h444;
rom[856] = 12'h444;
rom[857] = 12'h444;
rom[858] = 12'h444;
rom[859] = 12'h444;
rom[860] = 12'h444;
rom[861] = 12'h444;
rom[862] = 12'h555;
rom[863] = 12'h555;
rom[864] = 12'h444;
rom[865] = 12'h444;
rom[866] = 12'h555;
rom[867] = 12'h555;
rom[868] = 12'h555;
rom[869] = 12'h555;
rom[870] = 12'h555;
rom[871] = 12'h555;
rom[872] = 12'h666;
rom[873] = 12'h666;
rom[874] = 12'h666;
rom[875] = 12'h666;
rom[876] = 12'h666;
rom[877] = 12'h666;
rom[878] = 12'h666;
rom[879] = 12'h666;
rom[880] = 12'h666;
rom[881] = 12'h666;
rom[882] = 12'h666;
rom[883] = 12'h666;
rom[884] = 12'h666;
rom[885] = 12'h666;
rom[886] = 12'h666;
rom[887] = 12'h666;
rom[888] = 12'h666;
rom[889] = 12'h666;
rom[890] = 12'h666;
rom[891] = 12'h666;
rom[892] = 12'h666;
rom[893] = 12'h666;
rom[894] = 12'h666;
rom[895] = 12'h777;
rom[896] = 12'h777;
rom[897] = 12'h777;
rom[898] = 12'h777;
rom[899] = 12'h777;
rom[900] = 12'h777;
rom[901] = 12'h777;
rom[902] = 12'h777;
rom[903] = 12'h777;
rom[904] = 12'h888;
rom[905] = 12'h888;
rom[906] = 12'h888;
rom[907] = 12'h888;
rom[908] = 12'h888;
rom[909] = 12'h888;
rom[910] = 12'h999;
rom[911] = 12'h999;
rom[912] = 12'h999;
rom[913] = 12'h999;
rom[914] = 12'h999;
rom[915] = 12'h999;
rom[916] = 12'h999;
rom[917] = 12'h999;
rom[918] = 12'ha9a;
rom[919] = 12'ha9a;
rom[920] = 12'ha9a;
rom[921] = 12'ha9a;
rom[922] = 12'haaa;
rom[923] = 12'hbaa;
rom[924] = 12'hbaa;
rom[925] = 12'hbaa;
rom[926] = 12'hbbb;
rom[927] = 12'hbbb;
rom[928] = 12'haaa;
rom[929] = 12'haaa;
rom[930] = 12'haaa;
rom[931] = 12'haaa;
rom[932] = 12'haaa;
rom[933] = 12'haaa;
rom[934] = 12'haaa;
rom[935] = 12'haaa;
rom[936] = 12'haaa;
rom[937] = 12'haaa;
rom[938] = 12'ha9a;
rom[939] = 12'ha9a;
rom[940] = 12'h999;
rom[941] = 12'h999;
rom[942] = 12'h999;
rom[943] = 12'h988;
rom[944] = 12'h888;
rom[945] = 12'h888;
rom[946] = 12'h877;
rom[947] = 12'h777;
rom[948] = 12'h777;
rom[949] = 12'h777;
rom[950] = 12'h777;
rom[951] = 12'h776;
rom[952] = 12'h676;
rom[953] = 12'h666;
rom[954] = 12'h666;
rom[955] = 12'h666;
rom[956] = 12'h566;
rom[957] = 12'h565;
rom[958] = 12'h565;
rom[959] = 12'h565;
rom[960] = 12'h556;
rom[961] = 12'h555;
rom[962] = 12'h555;
rom[963] = 12'h555;
rom[964] = 12'h545;
rom[965] = 12'h445;
rom[966] = 12'h444;
rom[967] = 12'h444;
rom[968] = 12'h333;
rom[969] = 12'h333;
rom[970] = 12'h333;
rom[971] = 12'h333;
rom[972] = 12'h333;
rom[973] = 12'h334;
rom[974] = 12'h333;
rom[975] = 12'h333;
rom[976] = 12'h333;
rom[977] = 12'h333;
rom[978] = 12'h333;
rom[979] = 12'h333;
rom[980] = 12'h333;
rom[981] = 12'h333;
rom[982] = 12'h333;
rom[983] = 12'h333;
rom[984] = 12'h444;
rom[985] = 12'h444;
rom[986] = 12'h444;
rom[987] = 12'h444;
rom[988] = 12'h444;
rom[989] = 12'h444;
rom[990] = 12'h444;
rom[991] = 12'h333;
rom[992] = 12'h444;
rom[993] = 12'h444;
rom[994] = 12'h555;
rom[995] = 12'h666;
rom[996] = 12'h666;
rom[997] = 12'h666;
rom[998] = 12'h777;
rom[999] = 12'h777;
rom[1000] = 12'h555;
rom[1001] = 12'h444;
rom[1002] = 12'h444;
rom[1003] = 12'h444;
rom[1004] = 12'h444;
rom[1005] = 12'h444;
rom[1006] = 12'h444;
rom[1007] = 12'h333;
rom[1008] = 12'h222;
rom[1009] = 12'h111;
rom[1010] = 12'h  0;
rom[1011] = 12'h  0;
rom[1012] = 12'h111;
rom[1013] = 12'h  0;
rom[1014] = 12'h  0;
rom[1015] = 12'h  0;
rom[1016] = 12'h  0;
rom[1017] = 12'h111;
rom[1018] = 12'h222;
rom[1019] = 12'h222;
rom[1020] = 12'h111;
rom[1021] = 12'h  0;
rom[1022] = 12'h  0;
rom[1023] = 12'h  0;
rom[1024] = 12'h  0;
rom[1025] = 12'h  0;
rom[1026] = 12'h  0;
rom[1027] = 12'h  0;
rom[1028] = 12'h  0;
rom[1029] = 12'h  0;
rom[1030] = 12'h  0;
rom[1031] = 12'h  0;
rom[1032] = 12'h  0;
rom[1033] = 12'h  0;
rom[1034] = 12'h  0;
rom[1035] = 12'h  0;
rom[1036] = 12'h  0;
rom[1037] = 12'h  0;
rom[1038] = 12'h  0;
rom[1039] = 12'h  0;
rom[1040] = 12'h  0;
rom[1041] = 12'h  0;
rom[1042] = 12'h  0;
rom[1043] = 12'h  0;
rom[1044] = 12'h  0;
rom[1045] = 12'h  0;
rom[1046] = 12'h  0;
rom[1047] = 12'h  0;
rom[1048] = 12'h  0;
rom[1049] = 12'h  0;
rom[1050] = 12'h  0;
rom[1051] = 12'h  0;
rom[1052] = 12'h  0;
rom[1053] = 12'h  0;
rom[1054] = 12'h111;
rom[1055] = 12'h111;
rom[1056] = 12'h111;
rom[1057] = 12'h111;
rom[1058] = 12'h  0;
rom[1059] = 12'h  0;
rom[1060] = 12'h111;
rom[1061] = 12'h222;
rom[1062] = 12'h333;
rom[1063] = 12'h333;
rom[1064] = 12'h333;
rom[1065] = 12'h222;
rom[1066] = 12'h  0;
rom[1067] = 12'h  0;
rom[1068] = 12'h  0;
rom[1069] = 12'h  0;
rom[1070] = 12'h  0;
rom[1071] = 12'h  0;
rom[1072] = 12'h  0;
rom[1073] = 12'h  0;
rom[1074] = 12'h  0;
rom[1075] = 12'h  0;
rom[1076] = 12'h  0;
rom[1077] = 12'h  0;
rom[1078] = 12'h  0;
rom[1079] = 12'h  0;
rom[1080] = 12'h  0;
rom[1081] = 12'h  0;
rom[1082] = 12'h  0;
rom[1083] = 12'h  0;
rom[1084] = 12'h  0;
rom[1085] = 12'h  0;
rom[1086] = 12'h  0;
rom[1087] = 12'h  0;
rom[1088] = 12'h  0;
rom[1089] = 12'h  0;
rom[1090] = 12'h  0;
rom[1091] = 12'h  0;
rom[1092] = 12'h  0;
rom[1093] = 12'h  0;
rom[1094] = 12'h  0;
rom[1095] = 12'h  0;
rom[1096] = 12'h  0;
rom[1097] = 12'h  0;
rom[1098] = 12'h  0;
rom[1099] = 12'h  0;
rom[1100] = 12'h111;
rom[1101] = 12'h111;
rom[1102] = 12'h111;
rom[1103] = 12'h111;
rom[1104] = 12'h  0;
rom[1105] = 12'h  0;
rom[1106] = 12'h  0;
rom[1107] = 12'h  0;
rom[1108] = 12'h  0;
rom[1109] = 12'h  0;
rom[1110] = 12'h  0;
rom[1111] = 12'h  0;
rom[1112] = 12'h  0;
rom[1113] = 12'h  0;
rom[1114] = 12'h  0;
rom[1115] = 12'h  0;
rom[1116] = 12'h  0;
rom[1117] = 12'h  0;
rom[1118] = 12'h  0;
rom[1119] = 12'h  0;
rom[1120] = 12'h111;
rom[1121] = 12'h111;
rom[1122] = 12'h222;
rom[1123] = 12'h444;
rom[1124] = 12'h555;
rom[1125] = 12'h444;
rom[1126] = 12'h444;
rom[1127] = 12'h333;
rom[1128] = 12'h222;
rom[1129] = 12'h111;
rom[1130] = 12'h111;
rom[1131] = 12'h111;
rom[1132] = 12'h111;
rom[1133] = 12'h111;
rom[1134] = 12'h111;
rom[1135] = 12'h111;
rom[1136] = 12'h111;
rom[1137] = 12'h111;
rom[1138] = 12'h111;
rom[1139] = 12'h111;
rom[1140] = 12'h111;
rom[1141] = 12'h111;
rom[1142] = 12'h111;
rom[1143] = 12'h222;
rom[1144] = 12'h222;
rom[1145] = 12'h222;
rom[1146] = 12'h222;
rom[1147] = 12'h222;
rom[1148] = 12'h333;
rom[1149] = 12'h333;
rom[1150] = 12'h333;
rom[1151] = 12'h333;
rom[1152] = 12'h333;
rom[1153] = 12'h333;
rom[1154] = 12'h555;
rom[1155] = 12'h666;
rom[1156] = 12'h666;
rom[1157] = 12'h666;
rom[1158] = 12'h666;
rom[1159] = 12'h555;
rom[1160] = 12'h555;
rom[1161] = 12'h555;
rom[1162] = 12'h555;
rom[1163] = 12'h555;
rom[1164] = 12'h555;
rom[1165] = 12'h666;
rom[1166] = 12'h666;
rom[1167] = 12'h666;
rom[1168] = 12'h666;
rom[1169] = 12'h666;
rom[1170] = 12'h666;
rom[1171] = 12'h666;
rom[1172] = 12'h777;
rom[1173] = 12'h777;
rom[1174] = 12'h777;
rom[1175] = 12'h777;
rom[1176] = 12'h777;
rom[1177] = 12'h888;
rom[1178] = 12'h999;
rom[1179] = 12'haaa;
rom[1180] = 12'haaa;
rom[1181] = 12'haaa;
rom[1182] = 12'h999;
rom[1183] = 12'h999;
rom[1184] = 12'h888;
rom[1185] = 12'h888;
rom[1186] = 12'h888;
rom[1187] = 12'h888;
rom[1188] = 12'h888;
rom[1189] = 12'h999;
rom[1190] = 12'h999;
rom[1191] = 12'h999;
rom[1192] = 12'haaa;
rom[1193] = 12'haaa;
rom[1194] = 12'h999;
rom[1195] = 12'h999;
rom[1196] = 12'h999;
rom[1197] = 12'h999;
rom[1198] = 12'h999;
rom[1199] = 12'h999;
rom[1200] = 12'h444;
rom[1201] = 12'h444;
rom[1202] = 12'h444;
rom[1203] = 12'h444;
rom[1204] = 12'h444;
rom[1205] = 12'h444;
rom[1206] = 12'h444;
rom[1207] = 12'h444;
rom[1208] = 12'h444;
rom[1209] = 12'h444;
rom[1210] = 12'h444;
rom[1211] = 12'h444;
rom[1212] = 12'h444;
rom[1213] = 12'h444;
rom[1214] = 12'h444;
rom[1215] = 12'h444;
rom[1216] = 12'h444;
rom[1217] = 12'h444;
rom[1218] = 12'h444;
rom[1219] = 12'h444;
rom[1220] = 12'h444;
rom[1221] = 12'h444;
rom[1222] = 12'h444;
rom[1223] = 12'h444;
rom[1224] = 12'h555;
rom[1225] = 12'h555;
rom[1226] = 12'h555;
rom[1227] = 12'h555;
rom[1228] = 12'h555;
rom[1229] = 12'h555;
rom[1230] = 12'h555;
rom[1231] = 12'h555;
rom[1232] = 12'h555;
rom[1233] = 12'h555;
rom[1234] = 12'h555;
rom[1235] = 12'h555;
rom[1236] = 12'h555;
rom[1237] = 12'h444;
rom[1238] = 12'h444;
rom[1239] = 12'h444;
rom[1240] = 12'h444;
rom[1241] = 12'h444;
rom[1242] = 12'h444;
rom[1243] = 12'h333;
rom[1244] = 12'h333;
rom[1245] = 12'h333;
rom[1246] = 12'h333;
rom[1247] = 12'h333;
rom[1248] = 12'h333;
rom[1249] = 12'h333;
rom[1250] = 12'h333;
rom[1251] = 12'h333;
rom[1252] = 12'h333;
rom[1253] = 12'h333;
rom[1254] = 12'h333;
rom[1255] = 12'h333;
rom[1256] = 12'h333;
rom[1257] = 12'h333;
rom[1258] = 12'h333;
rom[1259] = 12'h333;
rom[1260] = 12'h444;
rom[1261] = 12'h444;
rom[1262] = 12'h444;
rom[1263] = 12'h444;
rom[1264] = 12'h444;
rom[1265] = 12'h444;
rom[1266] = 12'h444;
rom[1267] = 12'h444;
rom[1268] = 12'h444;
rom[1269] = 12'h444;
rom[1270] = 12'h444;
rom[1271] = 12'h444;
rom[1272] = 12'h444;
rom[1273] = 12'h444;
rom[1274] = 12'h444;
rom[1275] = 12'h555;
rom[1276] = 12'h555;
rom[1277] = 12'h555;
rom[1278] = 12'h555;
rom[1279] = 12'h555;
rom[1280] = 12'h555;
rom[1281] = 12'h555;
rom[1282] = 12'h555;
rom[1283] = 12'h666;
rom[1284] = 12'h666;
rom[1285] = 12'h666;
rom[1286] = 12'h666;
rom[1287] = 12'h666;
rom[1288] = 12'h666;
rom[1289] = 12'h666;
rom[1290] = 12'h666;
rom[1291] = 12'h666;
rom[1292] = 12'h666;
rom[1293] = 12'h666;
rom[1294] = 12'h666;
rom[1295] = 12'h666;
rom[1296] = 12'h777;
rom[1297] = 12'h777;
rom[1298] = 12'h777;
rom[1299] = 12'h777;
rom[1300] = 12'h777;
rom[1301] = 12'h777;
rom[1302] = 12'h777;
rom[1303] = 12'h777;
rom[1304] = 12'h777;
rom[1305] = 12'h888;
rom[1306] = 12'h888;
rom[1307] = 12'h888;
rom[1308] = 12'h888;
rom[1309] = 12'h999;
rom[1310] = 12'h999;
rom[1311] = 12'h999;
rom[1312] = 12'h999;
rom[1313] = 12'h999;
rom[1314] = 12'h999;
rom[1315] = 12'h999;
rom[1316] = 12'h99a;
rom[1317] = 12'haaa;
rom[1318] = 12'haaa;
rom[1319] = 12'haaa;
rom[1320] = 12'haaa;
rom[1321] = 12'haab;
rom[1322] = 12'hbab;
rom[1323] = 12'hbab;
rom[1324] = 12'hbab;
rom[1325] = 12'hbbb;
rom[1326] = 12'hbbb;
rom[1327] = 12'hbbb;
rom[1328] = 12'hbbb;
rom[1329] = 12'hbbb;
rom[1330] = 12'hbab;
rom[1331] = 12'hbaa;
rom[1332] = 12'hbaa;
rom[1333] = 12'hbaa;
rom[1334] = 12'hbaa;
rom[1335] = 12'hbaa;
rom[1336] = 12'haaa;
rom[1337] = 12'haaa;
rom[1338] = 12'haaa;
rom[1339] = 12'ha9a;
rom[1340] = 12'ha9a;
rom[1341] = 12'ha99;
rom[1342] = 12'h999;
rom[1343] = 12'h999;
rom[1344] = 12'h999;
rom[1345] = 12'h988;
rom[1346] = 12'h888;
rom[1347] = 12'h877;
rom[1348] = 12'h777;
rom[1349] = 12'h777;
rom[1350] = 12'h777;
rom[1351] = 12'h766;
rom[1352] = 12'h766;
rom[1353] = 12'h666;
rom[1354] = 12'h666;
rom[1355] = 12'h666;
rom[1356] = 12'h666;
rom[1357] = 12'h666;
rom[1358] = 12'h666;
rom[1359] = 12'h666;
rom[1360] = 12'h666;
rom[1361] = 12'h556;
rom[1362] = 12'h555;
rom[1363] = 12'h555;
rom[1364] = 12'h555;
rom[1365] = 12'h555;
rom[1366] = 12'h444;
rom[1367] = 12'h444;
rom[1368] = 12'h444;
rom[1369] = 12'h333;
rom[1370] = 12'h333;
rom[1371] = 12'h333;
rom[1372] = 12'h333;
rom[1373] = 12'h333;
rom[1374] = 12'h334;
rom[1375] = 12'h334;
rom[1376] = 12'h333;
rom[1377] = 12'h333;
rom[1378] = 12'h333;
rom[1379] = 12'h333;
rom[1380] = 12'h333;
rom[1381] = 12'h333;
rom[1382] = 12'h333;
rom[1383] = 12'h444;
rom[1384] = 12'h444;
rom[1385] = 12'h444;
rom[1386] = 12'h444;
rom[1387] = 12'h444;
rom[1388] = 12'h555;
rom[1389] = 12'h555;
rom[1390] = 12'h444;
rom[1391] = 12'h333;
rom[1392] = 12'h444;
rom[1393] = 12'h444;
rom[1394] = 12'h555;
rom[1395] = 12'h666;
rom[1396] = 12'h666;
rom[1397] = 12'h666;
rom[1398] = 12'h777;
rom[1399] = 12'h777;
rom[1400] = 12'h555;
rom[1401] = 12'h444;
rom[1402] = 12'h444;
rom[1403] = 12'h444;
rom[1404] = 12'h444;
rom[1405] = 12'h444;
rom[1406] = 12'h444;
rom[1407] = 12'h333;
rom[1408] = 12'h222;
rom[1409] = 12'h111;
rom[1410] = 12'h  0;
rom[1411] = 12'h  0;
rom[1412] = 12'h111;
rom[1413] = 12'h  0;
rom[1414] = 12'h  0;
rom[1415] = 12'h  0;
rom[1416] = 12'h  0;
rom[1417] = 12'h111;
rom[1418] = 12'h222;
rom[1419] = 12'h222;
rom[1420] = 12'h111;
rom[1421] = 12'h  0;
rom[1422] = 12'h  0;
rom[1423] = 12'h  0;
rom[1424] = 12'h  0;
rom[1425] = 12'h  0;
rom[1426] = 12'h  0;
rom[1427] = 12'h  0;
rom[1428] = 12'h  0;
rom[1429] = 12'h  0;
rom[1430] = 12'h  0;
rom[1431] = 12'h  0;
rom[1432] = 12'h  0;
rom[1433] = 12'h  0;
rom[1434] = 12'h  0;
rom[1435] = 12'h  0;
rom[1436] = 12'h  0;
rom[1437] = 12'h  0;
rom[1438] = 12'h  0;
rom[1439] = 12'h  0;
rom[1440] = 12'h  0;
rom[1441] = 12'h  0;
rom[1442] = 12'h  0;
rom[1443] = 12'h  0;
rom[1444] = 12'h  0;
rom[1445] = 12'h  0;
rom[1446] = 12'h  0;
rom[1447] = 12'h  0;
rom[1448] = 12'h  0;
rom[1449] = 12'h  0;
rom[1450] = 12'h  0;
rom[1451] = 12'h  0;
rom[1452] = 12'h111;
rom[1453] = 12'h111;
rom[1454] = 12'h111;
rom[1455] = 12'h111;
rom[1456] = 12'h111;
rom[1457] = 12'h111;
rom[1458] = 12'h111;
rom[1459] = 12'h111;
rom[1460] = 12'h222;
rom[1461] = 12'h333;
rom[1462] = 12'h333;
rom[1463] = 12'h333;
rom[1464] = 12'h333;
rom[1465] = 12'h222;
rom[1466] = 12'h  0;
rom[1467] = 12'h  0;
rom[1468] = 12'h  0;
rom[1469] = 12'h  0;
rom[1470] = 12'h  0;
rom[1471] = 12'h  0;
rom[1472] = 12'h  0;
rom[1473] = 12'h  0;
rom[1474] = 12'h  0;
rom[1475] = 12'h  0;
rom[1476] = 12'h  0;
rom[1477] = 12'h  0;
rom[1478] = 12'h  0;
rom[1479] = 12'h  0;
rom[1480] = 12'h  0;
rom[1481] = 12'h  0;
rom[1482] = 12'h  0;
rom[1483] = 12'h  0;
rom[1484] = 12'h  0;
rom[1485] = 12'h  0;
rom[1486] = 12'h  0;
rom[1487] = 12'h  0;
rom[1488] = 12'h  0;
rom[1489] = 12'h  0;
rom[1490] = 12'h  0;
rom[1491] = 12'h  0;
rom[1492] = 12'h  0;
rom[1493] = 12'h  0;
rom[1494] = 12'h  0;
rom[1495] = 12'h  0;
rom[1496] = 12'h  0;
rom[1497] = 12'h  0;
rom[1498] = 12'h  0;
rom[1499] = 12'h  0;
rom[1500] = 12'h111;
rom[1501] = 12'h111;
rom[1502] = 12'h111;
rom[1503] = 12'h111;
rom[1504] = 12'h  0;
rom[1505] = 12'h  0;
rom[1506] = 12'h  0;
rom[1507] = 12'h  0;
rom[1508] = 12'h  0;
rom[1509] = 12'h  0;
rom[1510] = 12'h  0;
rom[1511] = 12'h  0;
rom[1512] = 12'h  0;
rom[1513] = 12'h  0;
rom[1514] = 12'h  0;
rom[1515] = 12'h  0;
rom[1516] = 12'h  0;
rom[1517] = 12'h  0;
rom[1518] = 12'h  0;
rom[1519] = 12'h  0;
rom[1520] = 12'h111;
rom[1521] = 12'h111;
rom[1522] = 12'h333;
rom[1523] = 12'h444;
rom[1524] = 12'h555;
rom[1525] = 12'h444;
rom[1526] = 12'h444;
rom[1527] = 12'h333;
rom[1528] = 12'h222;
rom[1529] = 12'h222;
rom[1530] = 12'h111;
rom[1531] = 12'h111;
rom[1532] = 12'h222;
rom[1533] = 12'h111;
rom[1534] = 12'h111;
rom[1535] = 12'h111;
rom[1536] = 12'h111;
rom[1537] = 12'h111;
rom[1538] = 12'h111;
rom[1539] = 12'h111;
rom[1540] = 12'h111;
rom[1541] = 12'h111;
rom[1542] = 12'h111;
rom[1543] = 12'h111;
rom[1544] = 12'h222;
rom[1545] = 12'h222;
rom[1546] = 12'h222;
rom[1547] = 12'h333;
rom[1548] = 12'h333;
rom[1549] = 12'h333;
rom[1550] = 12'h333;
rom[1551] = 12'h333;
rom[1552] = 12'h333;
rom[1553] = 12'h444;
rom[1554] = 12'h666;
rom[1555] = 12'h666;
rom[1556] = 12'h666;
rom[1557] = 12'h555;
rom[1558] = 12'h555;
rom[1559] = 12'h555;
rom[1560] = 12'h555;
rom[1561] = 12'h555;
rom[1562] = 12'h555;
rom[1563] = 12'h555;
rom[1564] = 12'h555;
rom[1565] = 12'h666;
rom[1566] = 12'h666;
rom[1567] = 12'h666;
rom[1568] = 12'h666;
rom[1569] = 12'h777;
rom[1570] = 12'h777;
rom[1571] = 12'h777;
rom[1572] = 12'h666;
rom[1573] = 12'h666;
rom[1574] = 12'h777;
rom[1575] = 12'h888;
rom[1576] = 12'h999;
rom[1577] = 12'haaa;
rom[1578] = 12'haaa;
rom[1579] = 12'haaa;
rom[1580] = 12'haaa;
rom[1581] = 12'h999;
rom[1582] = 12'h888;
rom[1583] = 12'h888;
rom[1584] = 12'h888;
rom[1585] = 12'h888;
rom[1586] = 12'h888;
rom[1587] = 12'h888;
rom[1588] = 12'h888;
rom[1589] = 12'h888;
rom[1590] = 12'h999;
rom[1591] = 12'h999;
rom[1592] = 12'haaa;
rom[1593] = 12'h999;
rom[1594] = 12'h999;
rom[1595] = 12'h999;
rom[1596] = 12'h999;
rom[1597] = 12'h999;
rom[1598] = 12'h999;
rom[1599] = 12'h999;
rom[1600] = 12'h444;
rom[1601] = 12'h444;
rom[1602] = 12'h444;
rom[1603] = 12'h444;
rom[1604] = 12'h444;
rom[1605] = 12'h444;
rom[1606] = 12'h444;
rom[1607] = 12'h444;
rom[1608] = 12'h444;
rom[1609] = 12'h444;
rom[1610] = 12'h444;
rom[1611] = 12'h444;
rom[1612] = 12'h444;
rom[1613] = 12'h444;
rom[1614] = 12'h444;
rom[1615] = 12'h444;
rom[1616] = 12'h444;
rom[1617] = 12'h444;
rom[1618] = 12'h444;
rom[1619] = 12'h444;
rom[1620] = 12'h444;
rom[1621] = 12'h444;
rom[1622] = 12'h444;
rom[1623] = 12'h444;
rom[1624] = 12'h555;
rom[1625] = 12'h555;
rom[1626] = 12'h555;
rom[1627] = 12'h555;
rom[1628] = 12'h555;
rom[1629] = 12'h555;
rom[1630] = 12'h555;
rom[1631] = 12'h555;
rom[1632] = 12'h444;
rom[1633] = 12'h444;
rom[1634] = 12'h444;
rom[1635] = 12'h444;
rom[1636] = 12'h444;
rom[1637] = 12'h444;
rom[1638] = 12'h333;
rom[1639] = 12'h333;
rom[1640] = 12'h333;
rom[1641] = 12'h333;
rom[1642] = 12'h333;
rom[1643] = 12'h333;
rom[1644] = 12'h333;
rom[1645] = 12'h333;
rom[1646] = 12'h333;
rom[1647] = 12'h333;
rom[1648] = 12'h333;
rom[1649] = 12'h333;
rom[1650] = 12'h333;
rom[1651] = 12'h333;
rom[1652] = 12'h333;
rom[1653] = 12'h333;
rom[1654] = 12'h333;
rom[1655] = 12'h333;
rom[1656] = 12'h333;
rom[1657] = 12'h333;
rom[1658] = 12'h333;
rom[1659] = 12'h333;
rom[1660] = 12'h333;
rom[1661] = 12'h333;
rom[1662] = 12'h333;
rom[1663] = 12'h333;
rom[1664] = 12'h333;
rom[1665] = 12'h333;
rom[1666] = 12'h333;
rom[1667] = 12'h333;
rom[1668] = 12'h333;
rom[1669] = 12'h333;
rom[1670] = 12'h333;
rom[1671] = 12'h333;
rom[1672] = 12'h333;
rom[1673] = 12'h333;
rom[1674] = 12'h444;
rom[1675] = 12'h444;
rom[1676] = 12'h444;
rom[1677] = 12'h444;
rom[1678] = 12'h444;
rom[1679] = 12'h444;
rom[1680] = 12'h444;
rom[1681] = 12'h444;
rom[1682] = 12'h555;
rom[1683] = 12'h555;
rom[1684] = 12'h555;
rom[1685] = 12'h555;
rom[1686] = 12'h555;
rom[1687] = 12'h555;
rom[1688] = 12'h666;
rom[1689] = 12'h666;
rom[1690] = 12'h666;
rom[1691] = 12'h666;
rom[1692] = 12'h666;
rom[1693] = 12'h666;
rom[1694] = 12'h777;
rom[1695] = 12'h777;
rom[1696] = 12'h777;
rom[1697] = 12'h777;
rom[1698] = 12'h777;
rom[1699] = 12'h777;
rom[1700] = 12'h777;
rom[1701] = 12'h777;
rom[1702] = 12'h777;
rom[1703] = 12'h777;
rom[1704] = 12'h777;
rom[1705] = 12'h888;
rom[1706] = 12'h888;
rom[1707] = 12'h888;
rom[1708] = 12'h888;
rom[1709] = 12'h999;
rom[1710] = 12'h999;
rom[1711] = 12'h999;
rom[1712] = 12'h999;
rom[1713] = 12'h999;
rom[1714] = 12'h99a;
rom[1715] = 12'h9aa;
rom[1716] = 12'haaa;
rom[1717] = 12'haab;
rom[1718] = 12'haab;
rom[1719] = 12'haab;
rom[1720] = 12'hbab;
rom[1721] = 12'hbbb;
rom[1722] = 12'hbbb;
rom[1723] = 12'hbbb;
rom[1724] = 12'hbbb;
rom[1725] = 12'hbbb;
rom[1726] = 12'hbbb;
rom[1727] = 12'hbbb;
rom[1728] = 12'hcbb;
rom[1729] = 12'hcbb;
rom[1730] = 12'hbbb;
rom[1731] = 12'hbbb;
rom[1732] = 12'hbab;
rom[1733] = 12'hbab;
rom[1734] = 12'hbab;
rom[1735] = 12'hbab;
rom[1736] = 12'haaa;
rom[1737] = 12'haaa;
rom[1738] = 12'ha9a;
rom[1739] = 12'ha9a;
rom[1740] = 12'ha9a;
rom[1741] = 12'ha9a;
rom[1742] = 12'ha99;
rom[1743] = 12'h999;
rom[1744] = 12'h999;
rom[1745] = 12'h999;
rom[1746] = 12'h988;
rom[1747] = 12'h888;
rom[1748] = 12'h888;
rom[1749] = 12'h877;
rom[1750] = 12'h777;
rom[1751] = 12'h777;
rom[1752] = 12'h777;
rom[1753] = 12'h777;
rom[1754] = 12'h777;
rom[1755] = 12'h767;
rom[1756] = 12'h766;
rom[1757] = 12'h666;
rom[1758] = 12'h666;
rom[1759] = 12'h666;
rom[1760] = 12'h666;
rom[1761] = 12'h666;
rom[1762] = 12'h555;
rom[1763] = 12'h555;
rom[1764] = 12'h555;
rom[1765] = 12'h555;
rom[1766] = 12'h555;
rom[1767] = 12'h545;
rom[1768] = 12'h444;
rom[1769] = 12'h444;
rom[1770] = 12'h334;
rom[1771] = 12'h333;
rom[1772] = 12'h333;
rom[1773] = 12'h333;
rom[1774] = 12'h333;
rom[1775] = 12'h334;
rom[1776] = 12'h444;
rom[1777] = 12'h444;
rom[1778] = 12'h333;
rom[1779] = 12'h333;
rom[1780] = 12'h333;
rom[1781] = 12'h333;
rom[1782] = 12'h444;
rom[1783] = 12'h444;
rom[1784] = 12'h444;
rom[1785] = 12'h444;
rom[1786] = 12'h444;
rom[1787] = 12'h444;
rom[1788] = 12'h555;
rom[1789] = 12'h555;
rom[1790] = 12'h444;
rom[1791] = 12'h444;
rom[1792] = 12'h444;
rom[1793] = 12'h444;
rom[1794] = 12'h555;
rom[1795] = 12'h555;
rom[1796] = 12'h666;
rom[1797] = 12'h777;
rom[1798] = 12'h777;
rom[1799] = 12'h777;
rom[1800] = 12'h666;
rom[1801] = 12'h555;
rom[1802] = 12'h444;
rom[1803] = 12'h555;
rom[1804] = 12'h444;
rom[1805] = 12'h444;
rom[1806] = 12'h444;
rom[1807] = 12'h333;
rom[1808] = 12'h222;
rom[1809] = 12'h111;
rom[1810] = 12'h  0;
rom[1811] = 12'h111;
rom[1812] = 12'h111;
rom[1813] = 12'h  0;
rom[1814] = 12'h  0;
rom[1815] = 12'h  0;
rom[1816] = 12'h  0;
rom[1817] = 12'h222;
rom[1818] = 12'h222;
rom[1819] = 12'h222;
rom[1820] = 12'h  0;
rom[1821] = 12'h  0;
rom[1822] = 12'h  0;
rom[1823] = 12'h  0;
rom[1824] = 12'h  0;
rom[1825] = 12'h  0;
rom[1826] = 12'h  0;
rom[1827] = 12'h  0;
rom[1828] = 12'h  0;
rom[1829] = 12'h  0;
rom[1830] = 12'h  0;
rom[1831] = 12'h  0;
rom[1832] = 12'h  0;
rom[1833] = 12'h  0;
rom[1834] = 12'h  0;
rom[1835] = 12'h  0;
rom[1836] = 12'h  0;
rom[1837] = 12'h  0;
rom[1838] = 12'h  0;
rom[1839] = 12'h  0;
rom[1840] = 12'h  0;
rom[1841] = 12'h  0;
rom[1842] = 12'h  0;
rom[1843] = 12'h  0;
rom[1844] = 12'h  0;
rom[1845] = 12'h  0;
rom[1846] = 12'h  0;
rom[1847] = 12'h  0;
rom[1848] = 12'h  0;
rom[1849] = 12'h  0;
rom[1850] = 12'h111;
rom[1851] = 12'h111;
rom[1852] = 12'h111;
rom[1853] = 12'h111;
rom[1854] = 12'h111;
rom[1855] = 12'h111;
rom[1856] = 12'h  0;
rom[1857] = 12'h  0;
rom[1858] = 12'h111;
rom[1859] = 12'h222;
rom[1860] = 12'h222;
rom[1861] = 12'h333;
rom[1862] = 12'h333;
rom[1863] = 12'h222;
rom[1864] = 12'h222;
rom[1865] = 12'h111;
rom[1866] = 12'h  0;
rom[1867] = 12'h  0;
rom[1868] = 12'h  0;
rom[1869] = 12'h  0;
rom[1870] = 12'h  0;
rom[1871] = 12'h  0;
rom[1872] = 12'h  0;
rom[1873] = 12'h  0;
rom[1874] = 12'h  0;
rom[1875] = 12'h  0;
rom[1876] = 12'h  0;
rom[1877] = 12'h  0;
rom[1878] = 12'h  0;
rom[1879] = 12'h  0;
rom[1880] = 12'h  0;
rom[1881] = 12'h  0;
rom[1882] = 12'h  0;
rom[1883] = 12'h  0;
rom[1884] = 12'h  0;
rom[1885] = 12'h  0;
rom[1886] = 12'h  0;
rom[1887] = 12'h  0;
rom[1888] = 12'h  0;
rom[1889] = 12'h  0;
rom[1890] = 12'h  0;
rom[1891] = 12'h  0;
rom[1892] = 12'h  0;
rom[1893] = 12'h  0;
rom[1894] = 12'h  0;
rom[1895] = 12'h  0;
rom[1896] = 12'h  0;
rom[1897] = 12'h  0;
rom[1898] = 12'h  0;
rom[1899] = 12'h  0;
rom[1900] = 12'h111;
rom[1901] = 12'h111;
rom[1902] = 12'h111;
rom[1903] = 12'h111;
rom[1904] = 12'h  0;
rom[1905] = 12'h  0;
rom[1906] = 12'h  0;
rom[1907] = 12'h  0;
rom[1908] = 12'h  0;
rom[1909] = 12'h  0;
rom[1910] = 12'h  0;
rom[1911] = 12'h  0;
rom[1912] = 12'h  0;
rom[1913] = 12'h  0;
rom[1914] = 12'h  0;
rom[1915] = 12'h  0;
rom[1916] = 12'h  0;
rom[1917] = 12'h  0;
rom[1918] = 12'h  0;
rom[1919] = 12'h  0;
rom[1920] = 12'h111;
rom[1921] = 12'h222;
rom[1922] = 12'h333;
rom[1923] = 12'h444;
rom[1924] = 12'h555;
rom[1925] = 12'h444;
rom[1926] = 12'h444;
rom[1927] = 12'h333;
rom[1928] = 12'h222;
rom[1929] = 12'h222;
rom[1930] = 12'h222;
rom[1931] = 12'h222;
rom[1932] = 12'h222;
rom[1933] = 12'h111;
rom[1934] = 12'h111;
rom[1935] = 12'h111;
rom[1936] = 12'h111;
rom[1937] = 12'h111;
rom[1938] = 12'h111;
rom[1939] = 12'h111;
rom[1940] = 12'h111;
rom[1941] = 12'h111;
rom[1942] = 12'h111;
rom[1943] = 12'h111;
rom[1944] = 12'h111;
rom[1945] = 12'h222;
rom[1946] = 12'h222;
rom[1947] = 12'h333;
rom[1948] = 12'h333;
rom[1949] = 12'h333;
rom[1950] = 12'h333;
rom[1951] = 12'h333;
rom[1952] = 12'h444;
rom[1953] = 12'h555;
rom[1954] = 12'h666;
rom[1955] = 12'h666;
rom[1956] = 12'h555;
rom[1957] = 12'h555;
rom[1958] = 12'h555;
rom[1959] = 12'h555;
rom[1960] = 12'h555;
rom[1961] = 12'h555;
rom[1962] = 12'h444;
rom[1963] = 12'h444;
rom[1964] = 12'h555;
rom[1965] = 12'h555;
rom[1966] = 12'h555;
rom[1967] = 12'h666;
rom[1968] = 12'h555;
rom[1969] = 12'h666;
rom[1970] = 12'h666;
rom[1971] = 12'h666;
rom[1972] = 12'h666;
rom[1973] = 12'h777;
rom[1974] = 12'h888;
rom[1975] = 12'h999;
rom[1976] = 12'haaa;
rom[1977] = 12'haaa;
rom[1978] = 12'haaa;
rom[1979] = 12'h999;
rom[1980] = 12'h888;
rom[1981] = 12'h777;
rom[1982] = 12'h777;
rom[1983] = 12'h777;
rom[1984] = 12'h777;
rom[1985] = 12'h777;
rom[1986] = 12'h777;
rom[1987] = 12'h777;
rom[1988] = 12'h777;
rom[1989] = 12'h888;
rom[1990] = 12'h999;
rom[1991] = 12'h999;
rom[1992] = 12'haaa;
rom[1993] = 12'h999;
rom[1994] = 12'h999;
rom[1995] = 12'h999;
rom[1996] = 12'h999;
rom[1997] = 12'h999;
rom[1998] = 12'h999;
rom[1999] = 12'h999;
rom[2000] = 12'h555;
rom[2001] = 12'h444;
rom[2002] = 12'h444;
rom[2003] = 12'h444;
rom[2004] = 12'h444;
rom[2005] = 12'h444;
rom[2006] = 12'h444;
rom[2007] = 12'h444;
rom[2008] = 12'h444;
rom[2009] = 12'h444;
rom[2010] = 12'h444;
rom[2011] = 12'h444;
rom[2012] = 12'h444;
rom[2013] = 12'h444;
rom[2014] = 12'h444;
rom[2015] = 12'h444;
rom[2016] = 12'h444;
rom[2017] = 12'h444;
rom[2018] = 12'h444;
rom[2019] = 12'h444;
rom[2020] = 12'h444;
rom[2021] = 12'h444;
rom[2022] = 12'h444;
rom[2023] = 12'h444;
rom[2024] = 12'h555;
rom[2025] = 12'h555;
rom[2026] = 12'h555;
rom[2027] = 12'h555;
rom[2028] = 12'h555;
rom[2029] = 12'h555;
rom[2030] = 12'h444;
rom[2031] = 12'h444;
rom[2032] = 12'h444;
rom[2033] = 12'h444;
rom[2034] = 12'h444;
rom[2035] = 12'h333;
rom[2036] = 12'h333;
rom[2037] = 12'h333;
rom[2038] = 12'h333;
rom[2039] = 12'h333;
rom[2040] = 12'h222;
rom[2041] = 12'h222;
rom[2042] = 12'h222;
rom[2043] = 12'h222;
rom[2044] = 12'h222;
rom[2045] = 12'h222;
rom[2046] = 12'h222;
rom[2047] = 12'h222;
rom[2048] = 12'h222;
rom[2049] = 12'h222;
rom[2050] = 12'h222;
rom[2051] = 12'h222;
rom[2052] = 12'h222;
rom[2053] = 12'h222;
rom[2054] = 12'h222;
rom[2055] = 12'h222;
rom[2056] = 12'h222;
rom[2057] = 12'h222;
rom[2058] = 12'h222;
rom[2059] = 12'h222;
rom[2060] = 12'h222;
rom[2061] = 12'h333;
rom[2062] = 12'h333;
rom[2063] = 12'h333;
rom[2064] = 12'h333;
rom[2065] = 12'h333;
rom[2066] = 12'h222;
rom[2067] = 12'h222;
rom[2068] = 12'h222;
rom[2069] = 12'h333;
rom[2070] = 12'h333;
rom[2071] = 12'h333;
rom[2072] = 12'h333;
rom[2073] = 12'h333;
rom[2074] = 12'h333;
rom[2075] = 12'h333;
rom[2076] = 12'h333;
rom[2077] = 12'h333;
rom[2078] = 12'h333;
rom[2079] = 12'h333;
rom[2080] = 12'h333;
rom[2081] = 12'h444;
rom[2082] = 12'h444;
rom[2083] = 12'h444;
rom[2084] = 12'h444;
rom[2085] = 12'h444;
rom[2086] = 12'h555;
rom[2087] = 12'h555;
rom[2088] = 12'h666;
rom[2089] = 12'h666;
rom[2090] = 12'h666;
rom[2091] = 12'h666;
rom[2092] = 12'h777;
rom[2093] = 12'h777;
rom[2094] = 12'h777;
rom[2095] = 12'h777;
rom[2096] = 12'h777;
rom[2097] = 12'h777;
rom[2098] = 12'h777;
rom[2099] = 12'h777;
rom[2100] = 12'h777;
rom[2101] = 12'h777;
rom[2102] = 12'h888;
rom[2103] = 12'h888;
rom[2104] = 12'h888;
rom[2105] = 12'h888;
rom[2106] = 12'h888;
rom[2107] = 12'h888;
rom[2108] = 12'h888;
rom[2109] = 12'h999;
rom[2110] = 12'h999;
rom[2111] = 12'h999;
rom[2112] = 12'h9aa;
rom[2113] = 12'h9aa;
rom[2114] = 12'haaa;
rom[2115] = 12'haaa;
rom[2116] = 12'haab;
rom[2117] = 12'haab;
rom[2118] = 12'haab;
rom[2119] = 12'haab;
rom[2120] = 12'hbbb;
rom[2121] = 12'hbbb;
rom[2122] = 12'hbbc;
rom[2123] = 12'hbbc;
rom[2124] = 12'hbbc;
rom[2125] = 12'hbbc;
rom[2126] = 12'hbbc;
rom[2127] = 12'hbbc;
rom[2128] = 12'hcbc;
rom[2129] = 12'hcbb;
rom[2130] = 12'hcbb;
rom[2131] = 12'hbbb;
rom[2132] = 12'hbab;
rom[2133] = 12'hbab;
rom[2134] = 12'hbab;
rom[2135] = 12'hbab;
rom[2136] = 12'haaa;
rom[2137] = 12'haaa;
rom[2138] = 12'haaa;
rom[2139] = 12'haaa;
rom[2140] = 12'ha9a;
rom[2141] = 12'ha9a;
rom[2142] = 12'ha99;
rom[2143] = 12'h999;
rom[2144] = 12'h999;
rom[2145] = 12'h989;
rom[2146] = 12'h989;
rom[2147] = 12'h989;
rom[2148] = 12'h989;
rom[2149] = 12'h888;
rom[2150] = 12'h888;
rom[2151] = 12'h878;
rom[2152] = 12'h877;
rom[2153] = 12'h777;
rom[2154] = 12'h777;
rom[2155] = 12'h777;
rom[2156] = 12'h767;
rom[2157] = 12'h666;
rom[2158] = 12'h666;
rom[2159] = 12'h666;
rom[2160] = 12'h666;
rom[2161] = 12'h666;
rom[2162] = 12'h666;
rom[2163] = 12'h666;
rom[2164] = 12'h656;
rom[2165] = 12'h555;
rom[2166] = 12'h555;
rom[2167] = 12'h555;
rom[2168] = 12'h555;
rom[2169] = 12'h555;
rom[2170] = 12'h444;
rom[2171] = 12'h444;
rom[2172] = 12'h334;
rom[2173] = 12'h333;
rom[2174] = 12'h333;
rom[2175] = 12'h333;
rom[2176] = 12'h444;
rom[2177] = 12'h444;
rom[2178] = 12'h444;
rom[2179] = 12'h444;
rom[2180] = 12'h444;
rom[2181] = 12'h444;
rom[2182] = 12'h444;
rom[2183] = 12'h444;
rom[2184] = 12'h444;
rom[2185] = 12'h444;
rom[2186] = 12'h444;
rom[2187] = 12'h444;
rom[2188] = 12'h555;
rom[2189] = 12'h555;
rom[2190] = 12'h555;
rom[2191] = 12'h444;
rom[2192] = 12'h444;
rom[2193] = 12'h555;
rom[2194] = 12'h555;
rom[2195] = 12'h555;
rom[2196] = 12'h666;
rom[2197] = 12'h777;
rom[2198] = 12'h777;
rom[2199] = 12'h777;
rom[2200] = 12'h666;
rom[2201] = 12'h555;
rom[2202] = 12'h555;
rom[2203] = 12'h555;
rom[2204] = 12'h444;
rom[2205] = 12'h444;
rom[2206] = 12'h444;
rom[2207] = 12'h333;
rom[2208] = 12'h222;
rom[2209] = 12'h111;
rom[2210] = 12'h111;
rom[2211] = 12'h111;
rom[2212] = 12'h111;
rom[2213] = 12'h  0;
rom[2214] = 12'h  0;
rom[2215] = 12'h111;
rom[2216] = 12'h111;
rom[2217] = 12'h222;
rom[2218] = 12'h222;
rom[2219] = 12'h111;
rom[2220] = 12'h  0;
rom[2221] = 12'h  0;
rom[2222] = 12'h  0;
rom[2223] = 12'h  0;
rom[2224] = 12'h  0;
rom[2225] = 12'h  0;
rom[2226] = 12'h  0;
rom[2227] = 12'h  0;
rom[2228] = 12'h  0;
rom[2229] = 12'h  0;
rom[2230] = 12'h  0;
rom[2231] = 12'h  0;
rom[2232] = 12'h  0;
rom[2233] = 12'h  0;
rom[2234] = 12'h  0;
rom[2235] = 12'h  0;
rom[2236] = 12'h  0;
rom[2237] = 12'h  0;
rom[2238] = 12'h  0;
rom[2239] = 12'h  0;
rom[2240] = 12'h  0;
rom[2241] = 12'h  0;
rom[2242] = 12'h  0;
rom[2243] = 12'h  0;
rom[2244] = 12'h  0;
rom[2245] = 12'h  0;
rom[2246] = 12'h  0;
rom[2247] = 12'h  0;
rom[2248] = 12'h  0;
rom[2249] = 12'h111;
rom[2250] = 12'h111;
rom[2251] = 12'h111;
rom[2252] = 12'h111;
rom[2253] = 12'h111;
rom[2254] = 12'h111;
rom[2255] = 12'h111;
rom[2256] = 12'h  0;
rom[2257] = 12'h111;
rom[2258] = 12'h111;
rom[2259] = 12'h222;
rom[2260] = 12'h333;
rom[2261] = 12'h333;
rom[2262] = 12'h333;
rom[2263] = 12'h222;
rom[2264] = 12'h222;
rom[2265] = 12'h111;
rom[2266] = 12'h  0;
rom[2267] = 12'h  0;
rom[2268] = 12'h  0;
rom[2269] = 12'h  0;
rom[2270] = 12'h  0;
rom[2271] = 12'h  0;
rom[2272] = 12'h  0;
rom[2273] = 12'h  0;
rom[2274] = 12'h  0;
rom[2275] = 12'h  0;
rom[2276] = 12'h  0;
rom[2277] = 12'h  0;
rom[2278] = 12'h  0;
rom[2279] = 12'h  0;
rom[2280] = 12'h  0;
rom[2281] = 12'h  0;
rom[2282] = 12'h  0;
rom[2283] = 12'h  0;
rom[2284] = 12'h  0;
rom[2285] = 12'h  0;
rom[2286] = 12'h  0;
rom[2287] = 12'h  0;
rom[2288] = 12'h  0;
rom[2289] = 12'h  0;
rom[2290] = 12'h  0;
rom[2291] = 12'h  0;
rom[2292] = 12'h  0;
rom[2293] = 12'h  0;
rom[2294] = 12'h  0;
rom[2295] = 12'h  0;
rom[2296] = 12'h  0;
rom[2297] = 12'h  0;
rom[2298] = 12'h  0;
rom[2299] = 12'h  0;
rom[2300] = 12'h111;
rom[2301] = 12'h111;
rom[2302] = 12'h111;
rom[2303] = 12'h111;
rom[2304] = 12'h111;
rom[2305] = 12'h  0;
rom[2306] = 12'h  0;
rom[2307] = 12'h  0;
rom[2308] = 12'h  0;
rom[2309] = 12'h  0;
rom[2310] = 12'h  0;
rom[2311] = 12'h  0;
rom[2312] = 12'h  0;
rom[2313] = 12'h  0;
rom[2314] = 12'h  0;
rom[2315] = 12'h  0;
rom[2316] = 12'h  0;
rom[2317] = 12'h  0;
rom[2318] = 12'h  0;
rom[2319] = 12'h  0;
rom[2320] = 12'h111;
rom[2321] = 12'h222;
rom[2322] = 12'h333;
rom[2323] = 12'h555;
rom[2324] = 12'h555;
rom[2325] = 12'h444;
rom[2326] = 12'h333;
rom[2327] = 12'h333;
rom[2328] = 12'h333;
rom[2329] = 12'h222;
rom[2330] = 12'h222;
rom[2331] = 12'h222;
rom[2332] = 12'h222;
rom[2333] = 12'h111;
rom[2334] = 12'h111;
rom[2335] = 12'h111;
rom[2336] = 12'h111;
rom[2337] = 12'h111;
rom[2338] = 12'h111;
rom[2339] = 12'h111;
rom[2340] = 12'h111;
rom[2341] = 12'h111;
rom[2342] = 12'h111;
rom[2343] = 12'h111;
rom[2344] = 12'h111;
rom[2345] = 12'h111;
rom[2346] = 12'h222;
rom[2347] = 12'h222;
rom[2348] = 12'h333;
rom[2349] = 12'h333;
rom[2350] = 12'h333;
rom[2351] = 12'h333;
rom[2352] = 12'h555;
rom[2353] = 12'h666;
rom[2354] = 12'h666;
rom[2355] = 12'h555;
rom[2356] = 12'h444;
rom[2357] = 12'h555;
rom[2358] = 12'h555;
rom[2359] = 12'h555;
rom[2360] = 12'h555;
rom[2361] = 12'h444;
rom[2362] = 12'h444;
rom[2363] = 12'h444;
rom[2364] = 12'h444;
rom[2365] = 12'h555;
rom[2366] = 12'h555;
rom[2367] = 12'h555;
rom[2368] = 12'h555;
rom[2369] = 12'h555;
rom[2370] = 12'h555;
rom[2371] = 12'h666;
rom[2372] = 12'h777;
rom[2373] = 12'h999;
rom[2374] = 12'h999;
rom[2375] = 12'h999;
rom[2376] = 12'h999;
rom[2377] = 12'h999;
rom[2378] = 12'h888;
rom[2379] = 12'h777;
rom[2380] = 12'h666;
rom[2381] = 12'h777;
rom[2382] = 12'h777;
rom[2383] = 12'h777;
rom[2384] = 12'h777;
rom[2385] = 12'h777;
rom[2386] = 12'h777;
rom[2387] = 12'h777;
rom[2388] = 12'h777;
rom[2389] = 12'h888;
rom[2390] = 12'h999;
rom[2391] = 12'h999;
rom[2392] = 12'haaa;
rom[2393] = 12'haaa;
rom[2394] = 12'h999;
rom[2395] = 12'h999;
rom[2396] = 12'h999;
rom[2397] = 12'h999;
rom[2398] = 12'h999;
rom[2399] = 12'h999;
rom[2400] = 12'h555;
rom[2401] = 12'h444;
rom[2402] = 12'h444;
rom[2403] = 12'h444;
rom[2404] = 12'h444;
rom[2405] = 12'h444;
rom[2406] = 12'h444;
rom[2407] = 12'h444;
rom[2408] = 12'h444;
rom[2409] = 12'h444;
rom[2410] = 12'h444;
rom[2411] = 12'h444;
rom[2412] = 12'h444;
rom[2413] = 12'h444;
rom[2414] = 12'h444;
rom[2415] = 12'h444;
rom[2416] = 12'h444;
rom[2417] = 12'h444;
rom[2418] = 12'h444;
rom[2419] = 12'h444;
rom[2420] = 12'h444;
rom[2421] = 12'h444;
rom[2422] = 12'h444;
rom[2423] = 12'h444;
rom[2424] = 12'h444;
rom[2425] = 12'h444;
rom[2426] = 12'h444;
rom[2427] = 12'h444;
rom[2428] = 12'h444;
rom[2429] = 12'h444;
rom[2430] = 12'h333;
rom[2431] = 12'h333;
rom[2432] = 12'h333;
rom[2433] = 12'h333;
rom[2434] = 12'h333;
rom[2435] = 12'h333;
rom[2436] = 12'h333;
rom[2437] = 12'h333;
rom[2438] = 12'h333;
rom[2439] = 12'h333;
rom[2440] = 12'h222;
rom[2441] = 12'h222;
rom[2442] = 12'h222;
rom[2443] = 12'h222;
rom[2444] = 12'h222;
rom[2445] = 12'h222;
rom[2446] = 12'h222;
rom[2447] = 12'h222;
rom[2448] = 12'h222;
rom[2449] = 12'h222;
rom[2450] = 12'h222;
rom[2451] = 12'h222;
rom[2452] = 12'h222;
rom[2453] = 12'h222;
rom[2454] = 12'h222;
rom[2455] = 12'h222;
rom[2456] = 12'h222;
rom[2457] = 12'h222;
rom[2458] = 12'h222;
rom[2459] = 12'h222;
rom[2460] = 12'h222;
rom[2461] = 12'h222;
rom[2462] = 12'h222;
rom[2463] = 12'h222;
rom[2464] = 12'h222;
rom[2465] = 12'h222;
rom[2466] = 12'h222;
rom[2467] = 12'h222;
rom[2468] = 12'h222;
rom[2469] = 12'h222;
rom[2470] = 12'h222;
rom[2471] = 12'h222;
rom[2472] = 12'h222;
rom[2473] = 12'h222;
rom[2474] = 12'h222;
rom[2475] = 12'h222;
rom[2476] = 12'h222;
rom[2477] = 12'h222;
rom[2478] = 12'h222;
rom[2479] = 12'h222;
rom[2480] = 12'h333;
rom[2481] = 12'h333;
rom[2482] = 12'h333;
rom[2483] = 12'h333;
rom[2484] = 12'h333;
rom[2485] = 12'h333;
rom[2486] = 12'h444;
rom[2487] = 12'h444;
rom[2488] = 12'h555;
rom[2489] = 12'h555;
rom[2490] = 12'h555;
rom[2491] = 12'h666;
rom[2492] = 12'h666;
rom[2493] = 12'h666;
rom[2494] = 12'h777;
rom[2495] = 12'h777;
rom[2496] = 12'h777;
rom[2497] = 12'h777;
rom[2498] = 12'h777;
rom[2499] = 12'h888;
rom[2500] = 12'h888;
rom[2501] = 12'h888;
rom[2502] = 12'h888;
rom[2503] = 12'h888;
rom[2504] = 12'h888;
rom[2505] = 12'h888;
rom[2506] = 12'h888;
rom[2507] = 12'h999;
rom[2508] = 12'h999;
rom[2509] = 12'h999;
rom[2510] = 12'h999;
rom[2511] = 12'h999;
rom[2512] = 12'haaa;
rom[2513] = 12'haaa;
rom[2514] = 12'haaa;
rom[2515] = 12'haaa;
rom[2516] = 12'haab;
rom[2517] = 12'haab;
rom[2518] = 12'habb;
rom[2519] = 12'habb;
rom[2520] = 12'hbbc;
rom[2521] = 12'hbbc;
rom[2522] = 12'hbcc;
rom[2523] = 12'hbcc;
rom[2524] = 12'hbcc;
rom[2525] = 12'hbcc;
rom[2526] = 12'hbcc;
rom[2527] = 12'hbcc;
rom[2528] = 12'hcbc;
rom[2529] = 12'hcbc;
rom[2530] = 12'hcbb;
rom[2531] = 12'hbbb;
rom[2532] = 12'hbbb;
rom[2533] = 12'hbbb;
rom[2534] = 12'hbbb;
rom[2535] = 12'hbbb;
rom[2536] = 12'hbab;
rom[2537] = 12'hbab;
rom[2538] = 12'hbab;
rom[2539] = 12'hbab;
rom[2540] = 12'hbaa;
rom[2541] = 12'haaa;
rom[2542] = 12'ha9a;
rom[2543] = 12'h999;
rom[2544] = 12'h999;
rom[2545] = 12'h999;
rom[2546] = 12'h989;
rom[2547] = 12'h989;
rom[2548] = 12'h989;
rom[2549] = 12'h989;
rom[2550] = 12'h989;
rom[2551] = 12'h888;
rom[2552] = 12'h878;
rom[2553] = 12'h888;
rom[2554] = 12'h878;
rom[2555] = 12'h778;
rom[2556] = 12'h777;
rom[2557] = 12'h777;
rom[2558] = 12'h667;
rom[2559] = 12'h667;
rom[2560] = 12'h667;
rom[2561] = 12'h666;
rom[2562] = 12'h666;
rom[2563] = 12'h666;
rom[2564] = 12'h666;
rom[2565] = 12'h666;
rom[2566] = 12'h666;
rom[2567] = 12'h555;
rom[2568] = 12'h555;
rom[2569] = 12'h555;
rom[2570] = 12'h555;
rom[2571] = 12'h444;
rom[2572] = 12'h444;
rom[2573] = 12'h444;
rom[2574] = 12'h333;
rom[2575] = 12'h333;
rom[2576] = 12'h444;
rom[2577] = 12'h444;
rom[2578] = 12'h444;
rom[2579] = 12'h444;
rom[2580] = 12'h444;
rom[2581] = 12'h444;
rom[2582] = 12'h444;
rom[2583] = 12'h444;
rom[2584] = 12'h444;
rom[2585] = 12'h444;
rom[2586] = 12'h444;
rom[2587] = 12'h444;
rom[2588] = 12'h444;
rom[2589] = 12'h555;
rom[2590] = 12'h555;
rom[2591] = 12'h555;
rom[2592] = 12'h555;
rom[2593] = 12'h555;
rom[2594] = 12'h555;
rom[2595] = 12'h555;
rom[2596] = 12'h666;
rom[2597] = 12'h777;
rom[2598] = 12'h777;
rom[2599] = 12'h777;
rom[2600] = 12'h777;
rom[2601] = 12'h555;
rom[2602] = 12'h555;
rom[2603] = 12'h555;
rom[2604] = 12'h555;
rom[2605] = 12'h444;
rom[2606] = 12'h444;
rom[2607] = 12'h333;
rom[2608] = 12'h222;
rom[2609] = 12'h111;
rom[2610] = 12'h111;
rom[2611] = 12'h111;
rom[2612] = 12'h111;
rom[2613] = 12'h111;
rom[2614] = 12'h111;
rom[2615] = 12'h111;
rom[2616] = 12'h111;
rom[2617] = 12'h222;
rom[2618] = 12'h222;
rom[2619] = 12'h111;
rom[2620] = 12'h  0;
rom[2621] = 12'h  0;
rom[2622] = 12'h  0;
rom[2623] = 12'h  0;
rom[2624] = 12'h  0;
rom[2625] = 12'h  0;
rom[2626] = 12'h  0;
rom[2627] = 12'h  0;
rom[2628] = 12'h  0;
rom[2629] = 12'h  0;
rom[2630] = 12'h  0;
rom[2631] = 12'h  0;
rom[2632] = 12'h  0;
rom[2633] = 12'h  0;
rom[2634] = 12'h  0;
rom[2635] = 12'h  0;
rom[2636] = 12'h  0;
rom[2637] = 12'h  0;
rom[2638] = 12'h  0;
rom[2639] = 12'h  0;
rom[2640] = 12'h  0;
rom[2641] = 12'h  0;
rom[2642] = 12'h  0;
rom[2643] = 12'h  0;
rom[2644] = 12'h  0;
rom[2645] = 12'h  0;
rom[2646] = 12'h  0;
rom[2647] = 12'h  0;
rom[2648] = 12'h111;
rom[2649] = 12'h111;
rom[2650] = 12'h111;
rom[2651] = 12'h111;
rom[2652] = 12'h111;
rom[2653] = 12'h111;
rom[2654] = 12'h111;
rom[2655] = 12'h111;
rom[2656] = 12'h111;
rom[2657] = 12'h111;
rom[2658] = 12'h222;
rom[2659] = 12'h333;
rom[2660] = 12'h333;
rom[2661] = 12'h333;
rom[2662] = 12'h222;
rom[2663] = 12'h222;
rom[2664] = 12'h222;
rom[2665] = 12'h111;
rom[2666] = 12'h  0;
rom[2667] = 12'h  0;
rom[2668] = 12'h  0;
rom[2669] = 12'h  0;
rom[2670] = 12'h  0;
rom[2671] = 12'h  0;
rom[2672] = 12'h111;
rom[2673] = 12'h  0;
rom[2674] = 12'h  0;
rom[2675] = 12'h  0;
rom[2676] = 12'h  0;
rom[2677] = 12'h  0;
rom[2678] = 12'h  0;
rom[2679] = 12'h  0;
rom[2680] = 12'h  0;
rom[2681] = 12'h  0;
rom[2682] = 12'h  0;
rom[2683] = 12'h  0;
rom[2684] = 12'h  0;
rom[2685] = 12'h  0;
rom[2686] = 12'h  0;
rom[2687] = 12'h  0;
rom[2688] = 12'h  0;
rom[2689] = 12'h  0;
rom[2690] = 12'h  0;
rom[2691] = 12'h  0;
rom[2692] = 12'h  0;
rom[2693] = 12'h  0;
rom[2694] = 12'h  0;
rom[2695] = 12'h  0;
rom[2696] = 12'h  0;
rom[2697] = 12'h  0;
rom[2698] = 12'h  0;
rom[2699] = 12'h  0;
rom[2700] = 12'h111;
rom[2701] = 12'h111;
rom[2702] = 12'h111;
rom[2703] = 12'h111;
rom[2704] = 12'h111;
rom[2705] = 12'h  0;
rom[2706] = 12'h  0;
rom[2707] = 12'h  0;
rom[2708] = 12'h  0;
rom[2709] = 12'h  0;
rom[2710] = 12'h  0;
rom[2711] = 12'h  0;
rom[2712] = 12'h  0;
rom[2713] = 12'h  0;
rom[2714] = 12'h  0;
rom[2715] = 12'h  0;
rom[2716] = 12'h  0;
rom[2717] = 12'h  0;
rom[2718] = 12'h111;
rom[2719] = 12'h111;
rom[2720] = 12'h111;
rom[2721] = 12'h222;
rom[2722] = 12'h444;
rom[2723] = 12'h555;
rom[2724] = 12'h555;
rom[2725] = 12'h444;
rom[2726] = 12'h333;
rom[2727] = 12'h333;
rom[2728] = 12'h333;
rom[2729] = 12'h222;
rom[2730] = 12'h222;
rom[2731] = 12'h222;
rom[2732] = 12'h222;
rom[2733] = 12'h111;
rom[2734] = 12'h111;
rom[2735] = 12'h111;
rom[2736] = 12'h111;
rom[2737] = 12'h111;
rom[2738] = 12'h111;
rom[2739] = 12'h111;
rom[2740] = 12'h111;
rom[2741] = 12'h111;
rom[2742] = 12'h111;
rom[2743] = 12'h111;
rom[2744] = 12'h111;
rom[2745] = 12'h111;
rom[2746] = 12'h222;
rom[2747] = 12'h222;
rom[2748] = 12'h222;
rom[2749] = 12'h333;
rom[2750] = 12'h333;
rom[2751] = 12'h444;
rom[2752] = 12'h666;
rom[2753] = 12'h666;
rom[2754] = 12'h555;
rom[2755] = 12'h444;
rom[2756] = 12'h444;
rom[2757] = 12'h555;
rom[2758] = 12'h555;
rom[2759] = 12'h555;
rom[2760] = 12'h555;
rom[2761] = 12'h444;
rom[2762] = 12'h444;
rom[2763] = 12'h444;
rom[2764] = 12'h444;
rom[2765] = 12'h555;
rom[2766] = 12'h555;
rom[2767] = 12'h555;
rom[2768] = 12'h666;
rom[2769] = 12'h555;
rom[2770] = 12'h666;
rom[2771] = 12'h777;
rom[2772] = 12'h999;
rom[2773] = 12'h999;
rom[2774] = 12'h999;
rom[2775] = 12'h999;
rom[2776] = 12'h888;
rom[2777] = 12'h777;
rom[2778] = 12'h666;
rom[2779] = 12'h666;
rom[2780] = 12'h666;
rom[2781] = 12'h666;
rom[2782] = 12'h777;
rom[2783] = 12'h777;
rom[2784] = 12'h777;
rom[2785] = 12'h777;
rom[2786] = 12'h777;
rom[2787] = 12'h777;
rom[2788] = 12'h777;
rom[2789] = 12'h888;
rom[2790] = 12'h888;
rom[2791] = 12'h999;
rom[2792] = 12'haaa;
rom[2793] = 12'haaa;
rom[2794] = 12'h999;
rom[2795] = 12'h999;
rom[2796] = 12'h999;
rom[2797] = 12'h999;
rom[2798] = 12'h999;
rom[2799] = 12'h999;
rom[2800] = 12'h444;
rom[2801] = 12'h444;
rom[2802] = 12'h444;
rom[2803] = 12'h444;
rom[2804] = 12'h444;
rom[2805] = 12'h444;
rom[2806] = 12'h444;
rom[2807] = 12'h444;
rom[2808] = 12'h444;
rom[2809] = 12'h444;
rom[2810] = 12'h444;
rom[2811] = 12'h444;
rom[2812] = 12'h444;
rom[2813] = 12'h444;
rom[2814] = 12'h444;
rom[2815] = 12'h444;
rom[2816] = 12'h444;
rom[2817] = 12'h444;
rom[2818] = 12'h444;
rom[2819] = 12'h444;
rom[2820] = 12'h444;
rom[2821] = 12'h444;
rom[2822] = 12'h444;
rom[2823] = 12'h444;
rom[2824] = 12'h444;
rom[2825] = 12'h444;
rom[2826] = 12'h444;
rom[2827] = 12'h333;
rom[2828] = 12'h333;
rom[2829] = 12'h333;
rom[2830] = 12'h333;
rom[2831] = 12'h222;
rom[2832] = 12'h222;
rom[2833] = 12'h333;
rom[2834] = 12'h333;
rom[2835] = 12'h333;
rom[2836] = 12'h333;
rom[2837] = 12'h333;
rom[2838] = 12'h333;
rom[2839] = 12'h222;
rom[2840] = 12'h222;
rom[2841] = 12'h222;
rom[2842] = 12'h222;
rom[2843] = 12'h222;
rom[2844] = 12'h222;
rom[2845] = 12'h222;
rom[2846] = 12'h222;
rom[2847] = 12'h222;
rom[2848] = 12'h222;
rom[2849] = 12'h222;
rom[2850] = 12'h222;
rom[2851] = 12'h222;
rom[2852] = 12'h222;
rom[2853] = 12'h222;
rom[2854] = 12'h222;
rom[2855] = 12'h222;
rom[2856] = 12'h222;
rom[2857] = 12'h222;
rom[2858] = 12'h222;
rom[2859] = 12'h222;
rom[2860] = 12'h222;
rom[2861] = 12'h222;
rom[2862] = 12'h222;
rom[2863] = 12'h222;
rom[2864] = 12'h222;
rom[2865] = 12'h222;
rom[2866] = 12'h222;
rom[2867] = 12'h111;
rom[2868] = 12'h111;
rom[2869] = 12'h111;
rom[2870] = 12'h111;
rom[2871] = 12'h222;
rom[2872] = 12'h111;
rom[2873] = 12'h111;
rom[2874] = 12'h222;
rom[2875] = 12'h222;
rom[2876] = 12'h222;
rom[2877] = 12'h222;
rom[2878] = 12'h222;
rom[2879] = 12'h222;
rom[2880] = 12'h222;
rom[2881] = 12'h222;
rom[2882] = 12'h333;
rom[2883] = 12'h333;
rom[2884] = 12'h333;
rom[2885] = 12'h333;
rom[2886] = 12'h333;
rom[2887] = 12'h333;
rom[2888] = 12'h444;
rom[2889] = 12'h444;
rom[2890] = 12'h444;
rom[2891] = 12'h555;
rom[2892] = 12'h555;
rom[2893] = 12'h666;
rom[2894] = 12'h666;
rom[2895] = 12'h666;
rom[2896] = 12'h777;
rom[2897] = 12'h777;
rom[2898] = 12'h777;
rom[2899] = 12'h888;
rom[2900] = 12'h888;
rom[2901] = 12'h888;
rom[2902] = 12'h999;
rom[2903] = 12'h999;
rom[2904] = 12'h999;
rom[2905] = 12'h999;
rom[2906] = 12'h999;
rom[2907] = 12'h999;
rom[2908] = 12'h999;
rom[2909] = 12'h999;
rom[2910] = 12'h999;
rom[2911] = 12'h99a;
rom[2912] = 12'h9aa;
rom[2913] = 12'haaa;
rom[2914] = 12'haaa;
rom[2915] = 12'haab;
rom[2916] = 12'habb;
rom[2917] = 12'hbbb;
rom[2918] = 12'hbbb;
rom[2919] = 12'hbbb;
rom[2920] = 12'hbbc;
rom[2921] = 12'hbcc;
rom[2922] = 12'hbcc;
rom[2923] = 12'hbcc;
rom[2924] = 12'hbcc;
rom[2925] = 12'hbcc;
rom[2926] = 12'hbcc;
rom[2927] = 12'hbbc;
rom[2928] = 12'hbbc;
rom[2929] = 12'hcbb;
rom[2930] = 12'hbbc;
rom[2931] = 12'hbbb;
rom[2932] = 12'hbbb;
rom[2933] = 12'hbbb;
rom[2934] = 12'hbbb;
rom[2935] = 12'hbbb;
rom[2936] = 12'hbbb;
rom[2937] = 12'hbbb;
rom[2938] = 12'hbbb;
rom[2939] = 12'hbbb;
rom[2940] = 12'hbbb;
rom[2941] = 12'hbab;
rom[2942] = 12'haaa;
rom[2943] = 12'ha9a;
rom[2944] = 12'ha9a;
rom[2945] = 12'ha9a;
rom[2946] = 12'h999;
rom[2947] = 12'h989;
rom[2948] = 12'h989;
rom[2949] = 12'h989;
rom[2950] = 12'h889;
rom[2951] = 12'h889;
rom[2952] = 12'h888;
rom[2953] = 12'h888;
rom[2954] = 12'h888;
rom[2955] = 12'h888;
rom[2956] = 12'h788;
rom[2957] = 12'h778;
rom[2958] = 12'h778;
rom[2959] = 12'h777;
rom[2960] = 12'h777;
rom[2961] = 12'h777;
rom[2962] = 12'h666;
rom[2963] = 12'h666;
rom[2964] = 12'h666;
rom[2965] = 12'h666;
rom[2966] = 12'h666;
rom[2967] = 12'h666;
rom[2968] = 12'h555;
rom[2969] = 12'h555;
rom[2970] = 12'h555;
rom[2971] = 12'h555;
rom[2972] = 12'h444;
rom[2973] = 12'h444;
rom[2974] = 12'h333;
rom[2975] = 12'h333;
rom[2976] = 12'h444;
rom[2977] = 12'h444;
rom[2978] = 12'h444;
rom[2979] = 12'h444;
rom[2980] = 12'h444;
rom[2981] = 12'h444;
rom[2982] = 12'h444;
rom[2983] = 12'h444;
rom[2984] = 12'h444;
rom[2985] = 12'h444;
rom[2986] = 12'h333;
rom[2987] = 12'h444;
rom[2988] = 12'h444;
rom[2989] = 12'h555;
rom[2990] = 12'h555;
rom[2991] = 12'h666;
rom[2992] = 12'h555;
rom[2993] = 12'h555;
rom[2994] = 12'h555;
rom[2995] = 12'h555;
rom[2996] = 12'h666;
rom[2997] = 12'h777;
rom[2998] = 12'h777;
rom[2999] = 12'h777;
rom[3000] = 12'h777;
rom[3001] = 12'h666;
rom[3002] = 12'h555;
rom[3003] = 12'h555;
rom[3004] = 12'h555;
rom[3005] = 12'h444;
rom[3006] = 12'h444;
rom[3007] = 12'h333;
rom[3008] = 12'h222;
rom[3009] = 12'h111;
rom[3010] = 12'h111;
rom[3011] = 12'h111;
rom[3012] = 12'h111;
rom[3013] = 12'h111;
rom[3014] = 12'h111;
rom[3015] = 12'h111;
rom[3016] = 12'h222;
rom[3017] = 12'h222;
rom[3018] = 12'h222;
rom[3019] = 12'h  0;
rom[3020] = 12'h  0;
rom[3021] = 12'h  0;
rom[3022] = 12'h  0;
rom[3023] = 12'h  0;
rom[3024] = 12'h  0;
rom[3025] = 12'h  0;
rom[3026] = 12'h  0;
rom[3027] = 12'h  0;
rom[3028] = 12'h  0;
rom[3029] = 12'h  0;
rom[3030] = 12'h  0;
rom[3031] = 12'h  0;
rom[3032] = 12'h  0;
rom[3033] = 12'h  0;
rom[3034] = 12'h  0;
rom[3035] = 12'h  0;
rom[3036] = 12'h  0;
rom[3037] = 12'h  0;
rom[3038] = 12'h  0;
rom[3039] = 12'h  0;
rom[3040] = 12'h  0;
rom[3041] = 12'h  0;
rom[3042] = 12'h  0;
rom[3043] = 12'h  0;
rom[3044] = 12'h  0;
rom[3045] = 12'h  0;
rom[3046] = 12'h  0;
rom[3047] = 12'h  0;
rom[3048] = 12'h111;
rom[3049] = 12'h111;
rom[3050] = 12'h111;
rom[3051] = 12'h111;
rom[3052] = 12'h111;
rom[3053] = 12'h111;
rom[3054] = 12'h111;
rom[3055] = 12'h111;
rom[3056] = 12'h111;
rom[3057] = 12'h222;
rom[3058] = 12'h222;
rom[3059] = 12'h333;
rom[3060] = 12'h333;
rom[3061] = 12'h333;
rom[3062] = 12'h222;
rom[3063] = 12'h111;
rom[3064] = 12'h111;
rom[3065] = 12'h111;
rom[3066] = 12'h  0;
rom[3067] = 12'h  0;
rom[3068] = 12'h  0;
rom[3069] = 12'h  0;
rom[3070] = 12'h  0;
rom[3071] = 12'h  0;
rom[3072] = 12'h111;
rom[3073] = 12'h111;
rom[3074] = 12'h  0;
rom[3075] = 12'h  0;
rom[3076] = 12'h  0;
rom[3077] = 12'h  0;
rom[3078] = 12'h  0;
rom[3079] = 12'h  0;
rom[3080] = 12'h  0;
rom[3081] = 12'h  0;
rom[3082] = 12'h  0;
rom[3083] = 12'h  0;
rom[3084] = 12'h  0;
rom[3085] = 12'h  0;
rom[3086] = 12'h  0;
rom[3087] = 12'h  0;
rom[3088] = 12'h  0;
rom[3089] = 12'h  0;
rom[3090] = 12'h  0;
rom[3091] = 12'h  0;
rom[3092] = 12'h  0;
rom[3093] = 12'h  0;
rom[3094] = 12'h  0;
rom[3095] = 12'h  0;
rom[3096] = 12'h  0;
rom[3097] = 12'h  0;
rom[3098] = 12'h  0;
rom[3099] = 12'h  0;
rom[3100] = 12'h111;
rom[3101] = 12'h111;
rom[3102] = 12'h111;
rom[3103] = 12'h111;
rom[3104] = 12'h111;
rom[3105] = 12'h  0;
rom[3106] = 12'h  0;
rom[3107] = 12'h  0;
rom[3108] = 12'h  0;
rom[3109] = 12'h  0;
rom[3110] = 12'h  0;
rom[3111] = 12'h  0;
rom[3112] = 12'h  0;
rom[3113] = 12'h  0;
rom[3114] = 12'h  0;
rom[3115] = 12'h  0;
rom[3116] = 12'h  0;
rom[3117] = 12'h  0;
rom[3118] = 12'h111;
rom[3119] = 12'h111;
rom[3120] = 12'h111;
rom[3121] = 12'h222;
rom[3122] = 12'h444;
rom[3123] = 12'h555;
rom[3124] = 12'h555;
rom[3125] = 12'h444;
rom[3126] = 12'h333;
rom[3127] = 12'h333;
rom[3128] = 12'h333;
rom[3129] = 12'h222;
rom[3130] = 12'h222;
rom[3131] = 12'h222;
rom[3132] = 12'h111;
rom[3133] = 12'h111;
rom[3134] = 12'h111;
rom[3135] = 12'h111;
rom[3136] = 12'h111;
rom[3137] = 12'h111;
rom[3138] = 12'h111;
rom[3139] = 12'h111;
rom[3140] = 12'h111;
rom[3141] = 12'h111;
rom[3142] = 12'h111;
rom[3143] = 12'h111;
rom[3144] = 12'h111;
rom[3145] = 12'h222;
rom[3146] = 12'h222;
rom[3147] = 12'h222;
rom[3148] = 12'h222;
rom[3149] = 12'h333;
rom[3150] = 12'h444;
rom[3151] = 12'h444;
rom[3152] = 12'h666;
rom[3153] = 12'h666;
rom[3154] = 12'h555;
rom[3155] = 12'h333;
rom[3156] = 12'h444;
rom[3157] = 12'h555;
rom[3158] = 12'h555;
rom[3159] = 12'h444;
rom[3160] = 12'h444;
rom[3161] = 12'h444;
rom[3162] = 12'h555;
rom[3163] = 12'h555;
rom[3164] = 12'h555;
rom[3165] = 12'h555;
rom[3166] = 12'h555;
rom[3167] = 12'h666;
rom[3168] = 12'h777;
rom[3169] = 12'h777;
rom[3170] = 12'h888;
rom[3171] = 12'h999;
rom[3172] = 12'h999;
rom[3173] = 12'h999;
rom[3174] = 12'h888;
rom[3175] = 12'h777;
rom[3176] = 12'h666;
rom[3177] = 12'h666;
rom[3178] = 12'h666;
rom[3179] = 12'h666;
rom[3180] = 12'h666;
rom[3181] = 12'h777;
rom[3182] = 12'h666;
rom[3183] = 12'h666;
rom[3184] = 12'h777;
rom[3185] = 12'h777;
rom[3186] = 12'h777;
rom[3187] = 12'h777;
rom[3188] = 12'h777;
rom[3189] = 12'h777;
rom[3190] = 12'h888;
rom[3191] = 12'h999;
rom[3192] = 12'haaa;
rom[3193] = 12'haaa;
rom[3194] = 12'haaa;
rom[3195] = 12'h999;
rom[3196] = 12'h999;
rom[3197] = 12'h999;
rom[3198] = 12'h999;
rom[3199] = 12'h999;
rom[3200] = 12'h555;
rom[3201] = 12'h444;
rom[3202] = 12'h444;
rom[3203] = 12'h444;
rom[3204] = 12'h333;
rom[3205] = 12'h444;
rom[3206] = 12'h444;
rom[3207] = 12'h444;
rom[3208] = 12'h444;
rom[3209] = 12'h444;
rom[3210] = 12'h444;
rom[3211] = 12'h444;
rom[3212] = 12'h444;
rom[3213] = 12'h444;
rom[3214] = 12'h444;
rom[3215] = 12'h444;
rom[3216] = 12'h444;
rom[3217] = 12'h444;
rom[3218] = 12'h444;
rom[3219] = 12'h444;
rom[3220] = 12'h444;
rom[3221] = 12'h444;
rom[3222] = 12'h444;
rom[3223] = 12'h444;
rom[3224] = 12'h333;
rom[3225] = 12'h333;
rom[3226] = 12'h333;
rom[3227] = 12'h222;
rom[3228] = 12'h222;
rom[3229] = 12'h222;
rom[3230] = 12'h222;
rom[3231] = 12'h222;
rom[3232] = 12'h222;
rom[3233] = 12'h222;
rom[3234] = 12'h222;
rom[3235] = 12'h222;
rom[3236] = 12'h222;
rom[3237] = 12'h222;
rom[3238] = 12'h222;
rom[3239] = 12'h222;
rom[3240] = 12'h222;
rom[3241] = 12'h222;
rom[3242] = 12'h222;
rom[3243] = 12'h222;
rom[3244] = 12'h111;
rom[3245] = 12'h111;
rom[3246] = 12'h111;
rom[3247] = 12'h111;
rom[3248] = 12'h111;
rom[3249] = 12'h111;
rom[3250] = 12'h111;
rom[3251] = 12'h111;
rom[3252] = 12'h111;
rom[3253] = 12'h111;
rom[3254] = 12'h111;
rom[3255] = 12'h111;
rom[3256] = 12'h111;
rom[3257] = 12'h111;
rom[3258] = 12'h111;
rom[3259] = 12'h111;
rom[3260] = 12'h111;
rom[3261] = 12'h111;
rom[3262] = 12'h222;
rom[3263] = 12'h222;
rom[3264] = 12'h111;
rom[3265] = 12'h111;
rom[3266] = 12'h111;
rom[3267] = 12'h111;
rom[3268] = 12'h111;
rom[3269] = 12'h111;
rom[3270] = 12'h111;
rom[3271] = 12'h111;
rom[3272] = 12'h111;
rom[3273] = 12'h111;
rom[3274] = 12'h111;
rom[3275] = 12'h111;
rom[3276] = 12'h111;
rom[3277] = 12'h111;
rom[3278] = 12'h111;
rom[3279] = 12'h111;
rom[3280] = 12'h222;
rom[3281] = 12'h222;
rom[3282] = 12'h222;
rom[3283] = 12'h222;
rom[3284] = 12'h222;
rom[3285] = 12'h333;
rom[3286] = 12'h333;
rom[3287] = 12'h333;
rom[3288] = 12'h333;
rom[3289] = 12'h444;
rom[3290] = 12'h444;
rom[3291] = 12'h444;
rom[3292] = 12'h555;
rom[3293] = 12'h555;
rom[3294] = 12'h555;
rom[3295] = 12'h555;
rom[3296] = 12'h666;
rom[3297] = 12'h666;
rom[3298] = 12'h666;
rom[3299] = 12'h777;
rom[3300] = 12'h888;
rom[3301] = 12'h888;
rom[3302] = 12'h999;
rom[3303] = 12'h999;
rom[3304] = 12'h999;
rom[3305] = 12'h999;
rom[3306] = 12'h999;
rom[3307] = 12'h999;
rom[3308] = 12'haaa;
rom[3309] = 12'haaa;
rom[3310] = 12'haaa;
rom[3311] = 12'haaa;
rom[3312] = 12'haaa;
rom[3313] = 12'haaa;
rom[3314] = 12'haaa;
rom[3315] = 12'habb;
rom[3316] = 12'hbbb;
rom[3317] = 12'hccc;
rom[3318] = 12'hccc;
rom[3319] = 12'hbcc;
rom[3320] = 12'hccc;
rom[3321] = 12'hccc;
rom[3322] = 12'hccc;
rom[3323] = 12'hccc;
rom[3324] = 12'hccc;
rom[3325] = 12'hccc;
rom[3326] = 12'hccc;
rom[3327] = 12'hccc;
rom[3328] = 12'hccc;
rom[3329] = 12'hccc;
rom[3330] = 12'hccc;
rom[3331] = 12'hccc;
rom[3332] = 12'hccc;
rom[3333] = 12'hccc;
rom[3334] = 12'hccc;
rom[3335] = 12'hccc;
rom[3336] = 12'hccc;
rom[3337] = 12'hccc;
rom[3338] = 12'hbcc;
rom[3339] = 12'hbbb;
rom[3340] = 12'hbbb;
rom[3341] = 12'hbbb;
rom[3342] = 12'hbbb;
rom[3343] = 12'habb;
rom[3344] = 12'haab;
rom[3345] = 12'haaa;
rom[3346] = 12'haaa;
rom[3347] = 12'h99a;
rom[3348] = 12'h99a;
rom[3349] = 12'h999;
rom[3350] = 12'h899;
rom[3351] = 12'h889;
rom[3352] = 12'h889;
rom[3353] = 12'h889;
rom[3354] = 12'h889;
rom[3355] = 12'h888;
rom[3356] = 12'h888;
rom[3357] = 12'h888;
rom[3358] = 12'h888;
rom[3359] = 12'h888;
rom[3360] = 12'h788;
rom[3361] = 12'h777;
rom[3362] = 12'h777;
rom[3363] = 12'h777;
rom[3364] = 12'h666;
rom[3365] = 12'h666;
rom[3366] = 12'h666;
rom[3367] = 12'h666;
rom[3368] = 12'h555;
rom[3369] = 12'h555;
rom[3370] = 12'h555;
rom[3371] = 12'h666;
rom[3372] = 12'h555;
rom[3373] = 12'h555;
rom[3374] = 12'h444;
rom[3375] = 12'h444;
rom[3376] = 12'h444;
rom[3377] = 12'h444;
rom[3378] = 12'h444;
rom[3379] = 12'h444;
rom[3380] = 12'h444;
rom[3381] = 12'h444;
rom[3382] = 12'h444;
rom[3383] = 12'h444;
rom[3384] = 12'h444;
rom[3385] = 12'h444;
rom[3386] = 12'h444;
rom[3387] = 12'h444;
rom[3388] = 12'h444;
rom[3389] = 12'h444;
rom[3390] = 12'h555;
rom[3391] = 12'h666;
rom[3392] = 12'h666;
rom[3393] = 12'h666;
rom[3394] = 12'h555;
rom[3395] = 12'h555;
rom[3396] = 12'h666;
rom[3397] = 12'h777;
rom[3398] = 12'h777;
rom[3399] = 12'h777;
rom[3400] = 12'h888;
rom[3401] = 12'h666;
rom[3402] = 12'h666;
rom[3403] = 12'h555;
rom[3404] = 12'h555;
rom[3405] = 12'h444;
rom[3406] = 12'h444;
rom[3407] = 12'h333;
rom[3408] = 12'h222;
rom[3409] = 12'h111;
rom[3410] = 12'h111;
rom[3411] = 12'h111;
rom[3412] = 12'h111;
rom[3413] = 12'h111;
rom[3414] = 12'h111;
rom[3415] = 12'h111;
rom[3416] = 12'h333;
rom[3417] = 12'h222;
rom[3418] = 12'h111;
rom[3419] = 12'h  0;
rom[3420] = 12'h  0;
rom[3421] = 12'h  0;
rom[3422] = 12'h  0;
rom[3423] = 12'h  0;
rom[3424] = 12'h  0;
rom[3425] = 12'h  0;
rom[3426] = 12'h  0;
rom[3427] = 12'h  0;
rom[3428] = 12'h  0;
rom[3429] = 12'h  0;
rom[3430] = 12'h  0;
rom[3431] = 12'h  0;
rom[3432] = 12'h  0;
rom[3433] = 12'h  0;
rom[3434] = 12'h  0;
rom[3435] = 12'h  0;
rom[3436] = 12'h  0;
rom[3437] = 12'h  0;
rom[3438] = 12'h  0;
rom[3439] = 12'h  0;
rom[3440] = 12'h  0;
rom[3441] = 12'h  0;
rom[3442] = 12'h  0;
rom[3443] = 12'h  0;
rom[3444] = 12'h  0;
rom[3445] = 12'h  0;
rom[3446] = 12'h111;
rom[3447] = 12'h111;
rom[3448] = 12'h111;
rom[3449] = 12'h111;
rom[3450] = 12'h111;
rom[3451] = 12'h111;
rom[3452] = 12'h111;
rom[3453] = 12'h111;
rom[3454] = 12'h111;
rom[3455] = 12'h111;
rom[3456] = 12'h111;
rom[3457] = 12'h333;
rom[3458] = 12'h333;
rom[3459] = 12'h333;
rom[3460] = 12'h222;
rom[3461] = 12'h222;
rom[3462] = 12'h222;
rom[3463] = 12'h222;
rom[3464] = 12'h222;
rom[3465] = 12'h111;
rom[3466] = 12'h  0;
rom[3467] = 12'h  0;
rom[3468] = 12'h  0;
rom[3469] = 12'h  0;
rom[3470] = 12'h  0;
rom[3471] = 12'h  0;
rom[3472] = 12'h  0;
rom[3473] = 12'h  0;
rom[3474] = 12'h  0;
rom[3475] = 12'h  0;
rom[3476] = 12'h  0;
rom[3477] = 12'h  0;
rom[3478] = 12'h  0;
rom[3479] = 12'h  0;
rom[3480] = 12'h  0;
rom[3481] = 12'h  0;
rom[3482] = 12'h  0;
rom[3483] = 12'h  0;
rom[3484] = 12'h  0;
rom[3485] = 12'h  0;
rom[3486] = 12'h  0;
rom[3487] = 12'h  0;
rom[3488] = 12'h  0;
rom[3489] = 12'h  0;
rom[3490] = 12'h  0;
rom[3491] = 12'h  0;
rom[3492] = 12'h  0;
rom[3493] = 12'h  0;
rom[3494] = 12'h  0;
rom[3495] = 12'h  0;
rom[3496] = 12'h  0;
rom[3497] = 12'h  0;
rom[3498] = 12'h  0;
rom[3499] = 12'h  0;
rom[3500] = 12'h111;
rom[3501] = 12'h111;
rom[3502] = 12'h111;
rom[3503] = 12'h111;
rom[3504] = 12'h111;
rom[3505] = 12'h  0;
rom[3506] = 12'h  0;
rom[3507] = 12'h  0;
rom[3508] = 12'h  0;
rom[3509] = 12'h  0;
rom[3510] = 12'h  0;
rom[3511] = 12'h  0;
rom[3512] = 12'h  0;
rom[3513] = 12'h  0;
rom[3514] = 12'h  0;
rom[3515] = 12'h  0;
rom[3516] = 12'h  0;
rom[3517] = 12'h111;
rom[3518] = 12'h111;
rom[3519] = 12'h111;
rom[3520] = 12'h222;
rom[3521] = 12'h222;
rom[3522] = 12'h444;
rom[3523] = 12'h555;
rom[3524] = 12'h555;
rom[3525] = 12'h444;
rom[3526] = 12'h333;
rom[3527] = 12'h444;
rom[3528] = 12'h333;
rom[3529] = 12'h222;
rom[3530] = 12'h222;
rom[3531] = 12'h222;
rom[3532] = 12'h111;
rom[3533] = 12'h111;
rom[3534] = 12'h111;
rom[3535] = 12'h111;
rom[3536] = 12'h111;
rom[3537] = 12'h111;
rom[3538] = 12'h111;
rom[3539] = 12'h111;
rom[3540] = 12'h111;
rom[3541] = 12'h111;
rom[3542] = 12'h111;
rom[3543] = 12'h111;
rom[3544] = 12'h111;
rom[3545] = 12'h111;
rom[3546] = 12'h222;
rom[3547] = 12'h222;
rom[3548] = 12'h333;
rom[3549] = 12'h333;
rom[3550] = 12'h444;
rom[3551] = 12'h666;
rom[3552] = 12'h555;
rom[3553] = 12'h444;
rom[3554] = 12'h333;
rom[3555] = 12'h444;
rom[3556] = 12'h444;
rom[3557] = 12'h444;
rom[3558] = 12'h444;
rom[3559] = 12'h444;
rom[3560] = 12'h444;
rom[3561] = 12'h555;
rom[3562] = 12'h555;
rom[3563] = 12'h555;
rom[3564] = 12'h555;
rom[3565] = 12'h555;
rom[3566] = 12'h666;
rom[3567] = 12'h777;
rom[3568] = 12'h888;
rom[3569] = 12'h999;
rom[3570] = 12'h999;
rom[3571] = 12'h999;
rom[3572] = 12'h888;
rom[3573] = 12'h666;
rom[3574] = 12'h555;
rom[3575] = 12'h555;
rom[3576] = 12'h666;
rom[3577] = 12'h666;
rom[3578] = 12'h666;
rom[3579] = 12'h666;
rom[3580] = 12'h666;
rom[3581] = 12'h666;
rom[3582] = 12'h666;
rom[3583] = 12'h666;
rom[3584] = 12'h666;
rom[3585] = 12'h777;
rom[3586] = 12'h777;
rom[3587] = 12'h666;
rom[3588] = 12'h777;
rom[3589] = 12'h777;
rom[3590] = 12'h888;
rom[3591] = 12'h999;
rom[3592] = 12'h999;
rom[3593] = 12'h999;
rom[3594] = 12'haaa;
rom[3595] = 12'h999;
rom[3596] = 12'h999;
rom[3597] = 12'h999;
rom[3598] = 12'h999;
rom[3599] = 12'h999;
rom[3600] = 12'h444;
rom[3601] = 12'h444;
rom[3602] = 12'h444;
rom[3603] = 12'h444;
rom[3604] = 12'h444;
rom[3605] = 12'h444;
rom[3606] = 12'h444;
rom[3607] = 12'h444;
rom[3608] = 12'h444;
rom[3609] = 12'h444;
rom[3610] = 12'h444;
rom[3611] = 12'h444;
rom[3612] = 12'h444;
rom[3613] = 12'h444;
rom[3614] = 12'h444;
rom[3615] = 12'h444;
rom[3616] = 12'h444;
rom[3617] = 12'h444;
rom[3618] = 12'h444;
rom[3619] = 12'h444;
rom[3620] = 12'h444;
rom[3621] = 12'h444;
rom[3622] = 12'h333;
rom[3623] = 12'h333;
rom[3624] = 12'h333;
rom[3625] = 12'h333;
rom[3626] = 12'h222;
rom[3627] = 12'h222;
rom[3628] = 12'h222;
rom[3629] = 12'h222;
rom[3630] = 12'h222;
rom[3631] = 12'h222;
rom[3632] = 12'h222;
rom[3633] = 12'h222;
rom[3634] = 12'h222;
rom[3635] = 12'h222;
rom[3636] = 12'h222;
rom[3637] = 12'h222;
rom[3638] = 12'h222;
rom[3639] = 12'h222;
rom[3640] = 12'h222;
rom[3641] = 12'h111;
rom[3642] = 12'h111;
rom[3643] = 12'h111;
rom[3644] = 12'h111;
rom[3645] = 12'h111;
rom[3646] = 12'h111;
rom[3647] = 12'h111;
rom[3648] = 12'h111;
rom[3649] = 12'h111;
rom[3650] = 12'h111;
rom[3651] = 12'h111;
rom[3652] = 12'h111;
rom[3653] = 12'h111;
rom[3654] = 12'h111;
rom[3655] = 12'h111;
rom[3656] = 12'h111;
rom[3657] = 12'h111;
rom[3658] = 12'h111;
rom[3659] = 12'h111;
rom[3660] = 12'h111;
rom[3661] = 12'h111;
rom[3662] = 12'h111;
rom[3663] = 12'h111;
rom[3664] = 12'h111;
rom[3665] = 12'h111;
rom[3666] = 12'h111;
rom[3667] = 12'h111;
rom[3668] = 12'h111;
rom[3669] = 12'h111;
rom[3670] = 12'h111;
rom[3671] = 12'h111;
rom[3672] = 12'h111;
rom[3673] = 12'h111;
rom[3674] = 12'h111;
rom[3675] = 12'h111;
rom[3676] = 12'h111;
rom[3677] = 12'h111;
rom[3678] = 12'h111;
rom[3679] = 12'h111;
rom[3680] = 12'h222;
rom[3681] = 12'h222;
rom[3682] = 12'h222;
rom[3683] = 12'h222;
rom[3684] = 12'h222;
rom[3685] = 12'h222;
rom[3686] = 12'h333;
rom[3687] = 12'h333;
rom[3688] = 12'h333;
rom[3689] = 12'h333;
rom[3690] = 12'h333;
rom[3691] = 12'h444;
rom[3692] = 12'h444;
rom[3693] = 12'h444;
rom[3694] = 12'h555;
rom[3695] = 12'h555;
rom[3696] = 12'h555;
rom[3697] = 12'h555;
rom[3698] = 12'h666;
rom[3699] = 12'h666;
rom[3700] = 12'h777;
rom[3701] = 12'h777;
rom[3702] = 12'h888;
rom[3703] = 12'h888;
rom[3704] = 12'h999;
rom[3705] = 12'h999;
rom[3706] = 12'h999;
rom[3707] = 12'h999;
rom[3708] = 12'haaa;
rom[3709] = 12'haaa;
rom[3710] = 12'haaa;
rom[3711] = 12'haaa;
rom[3712] = 12'haaa;
rom[3713] = 12'hbbb;
rom[3714] = 12'hbbb;
rom[3715] = 12'hbcb;
rom[3716] = 12'hccc;
rom[3717] = 12'hccc;
rom[3718] = 12'hcdc;
rom[3719] = 12'hcdc;
rom[3720] = 12'hddc;
rom[3721] = 12'hcdc;
rom[3722] = 12'hcdc;
rom[3723] = 12'hcdd;
rom[3724] = 12'hcdd;
rom[3725] = 12'hcdd;
rom[3726] = 12'hddd;
rom[3727] = 12'hddd;
rom[3728] = 12'hddd;
rom[3729] = 12'hddd;
rom[3730] = 12'hddd;
rom[3731] = 12'hddd;
rom[3732] = 12'hcdd;
rom[3733] = 12'hcdc;
rom[3734] = 12'hcdc;
rom[3735] = 12'hcdc;
rom[3736] = 12'hccc;
rom[3737] = 12'hccc;
rom[3738] = 12'hccc;
rom[3739] = 12'hbcc;
rom[3740] = 12'hbcb;
rom[3741] = 12'hbcb;
rom[3742] = 12'hbcb;
rom[3743] = 12'hbcc;
rom[3744] = 12'hbbc;
rom[3745] = 12'hbbb;
rom[3746] = 12'habb;
rom[3747] = 12'haaa;
rom[3748] = 12'haaa;
rom[3749] = 12'h99a;
rom[3750] = 12'h999;
rom[3751] = 12'h899;
rom[3752] = 12'h888;
rom[3753] = 12'h888;
rom[3754] = 12'h888;
rom[3755] = 12'h889;
rom[3756] = 12'h889;
rom[3757] = 12'h889;
rom[3758] = 12'h889;
rom[3759] = 12'h899;
rom[3760] = 12'h888;
rom[3761] = 12'h888;
rom[3762] = 12'h888;
rom[3763] = 12'h777;
rom[3764] = 12'h777;
rom[3765] = 12'h666;
rom[3766] = 12'h666;
rom[3767] = 12'h666;
rom[3768] = 12'h666;
rom[3769] = 12'h666;
rom[3770] = 12'h666;
rom[3771] = 12'h666;
rom[3772] = 12'h666;
rom[3773] = 12'h666;
rom[3774] = 12'h555;
rom[3775] = 12'h555;
rom[3776] = 12'h555;
rom[3777] = 12'h555;
rom[3778] = 12'h444;
rom[3779] = 12'h555;
rom[3780] = 12'h555;
rom[3781] = 12'h555;
rom[3782] = 12'h555;
rom[3783] = 12'h555;
rom[3784] = 12'h444;
rom[3785] = 12'h444;
rom[3786] = 12'h444;
rom[3787] = 12'h444;
rom[3788] = 12'h444;
rom[3789] = 12'h444;
rom[3790] = 12'h555;
rom[3791] = 12'h555;
rom[3792] = 12'h666;
rom[3793] = 12'h666;
rom[3794] = 12'h555;
rom[3795] = 12'h555;
rom[3796] = 12'h666;
rom[3797] = 12'h777;
rom[3798] = 12'h777;
rom[3799] = 12'h777;
rom[3800] = 12'h888;
rom[3801] = 12'h777;
rom[3802] = 12'h666;
rom[3803] = 12'h666;
rom[3804] = 12'h555;
rom[3805] = 12'h444;
rom[3806] = 12'h444;
rom[3807] = 12'h333;
rom[3808] = 12'h222;
rom[3809] = 12'h222;
rom[3810] = 12'h111;
rom[3811] = 12'h222;
rom[3812] = 12'h222;
rom[3813] = 12'h222;
rom[3814] = 12'h111;
rom[3815] = 12'h222;
rom[3816] = 12'h333;
rom[3817] = 12'h222;
rom[3818] = 12'h111;
rom[3819] = 12'h  0;
rom[3820] = 12'h  0;
rom[3821] = 12'h  0;
rom[3822] = 12'h  0;
rom[3823] = 12'h  0;
rom[3824] = 12'h  0;
rom[3825] = 12'h  0;
rom[3826] = 12'h  0;
rom[3827] = 12'h  0;
rom[3828] = 12'h  0;
rom[3829] = 12'h  0;
rom[3830] = 12'h  0;
rom[3831] = 12'h  0;
rom[3832] = 12'h  0;
rom[3833] = 12'h  0;
rom[3834] = 12'h  0;
rom[3835] = 12'h  0;
rom[3836] = 12'h  0;
rom[3837] = 12'h  0;
rom[3838] = 12'h  0;
rom[3839] = 12'h  0;
rom[3840] = 12'h  0;
rom[3841] = 12'h  0;
rom[3842] = 12'h  0;
rom[3843] = 12'h  0;
rom[3844] = 12'h  0;
rom[3845] = 12'h  0;
rom[3846] = 12'h111;
rom[3847] = 12'h111;
rom[3848] = 12'h111;
rom[3849] = 12'h111;
rom[3850] = 12'h111;
rom[3851] = 12'h111;
rom[3852] = 12'h111;
rom[3853] = 12'h111;
rom[3854] = 12'h111;
rom[3855] = 12'h111;
rom[3856] = 12'h222;
rom[3857] = 12'h333;
rom[3858] = 12'h333;
rom[3859] = 12'h222;
rom[3860] = 12'h222;
rom[3861] = 12'h222;
rom[3862] = 12'h222;
rom[3863] = 12'h222;
rom[3864] = 12'h111;
rom[3865] = 12'h111;
rom[3866] = 12'h  0;
rom[3867] = 12'h111;
rom[3868] = 12'h111;
rom[3869] = 12'h111;
rom[3870] = 12'h  0;
rom[3871] = 12'h  0;
rom[3872] = 12'h  0;
rom[3873] = 12'h  0;
rom[3874] = 12'h  0;
rom[3875] = 12'h  0;
rom[3876] = 12'h  0;
rom[3877] = 12'h  0;
rom[3878] = 12'h  0;
rom[3879] = 12'h  0;
rom[3880] = 12'h  0;
rom[3881] = 12'h  0;
rom[3882] = 12'h  0;
rom[3883] = 12'h  0;
rom[3884] = 12'h  0;
rom[3885] = 12'h  0;
rom[3886] = 12'h  0;
rom[3887] = 12'h  0;
rom[3888] = 12'h  0;
rom[3889] = 12'h  0;
rom[3890] = 12'h  0;
rom[3891] = 12'h  0;
rom[3892] = 12'h  0;
rom[3893] = 12'h  0;
rom[3894] = 12'h  0;
rom[3895] = 12'h  0;
rom[3896] = 12'h  0;
rom[3897] = 12'h  0;
rom[3898] = 12'h  0;
rom[3899] = 12'h  0;
rom[3900] = 12'h111;
rom[3901] = 12'h111;
rom[3902] = 12'h111;
rom[3903] = 12'h111;
rom[3904] = 12'h111;
rom[3905] = 12'h  0;
rom[3906] = 12'h  0;
rom[3907] = 12'h  0;
rom[3908] = 12'h  0;
rom[3909] = 12'h  0;
rom[3910] = 12'h  0;
rom[3911] = 12'h  0;
rom[3912] = 12'h  0;
rom[3913] = 12'h  0;
rom[3914] = 12'h  0;
rom[3915] = 12'h  0;
rom[3916] = 12'h  0;
rom[3917] = 12'h111;
rom[3918] = 12'h111;
rom[3919] = 12'h111;
rom[3920] = 12'h222;
rom[3921] = 12'h333;
rom[3922] = 12'h444;
rom[3923] = 12'h555;
rom[3924] = 12'h555;
rom[3925] = 12'h444;
rom[3926] = 12'h444;
rom[3927] = 12'h444;
rom[3928] = 12'h333;
rom[3929] = 12'h222;
rom[3930] = 12'h222;
rom[3931] = 12'h222;
rom[3932] = 12'h111;
rom[3933] = 12'h111;
rom[3934] = 12'h111;
rom[3935] = 12'h111;
rom[3936] = 12'h111;
rom[3937] = 12'h111;
rom[3938] = 12'h111;
rom[3939] = 12'h111;
rom[3940] = 12'h111;
rom[3941] = 12'h111;
rom[3942] = 12'h111;
rom[3943] = 12'h111;
rom[3944] = 12'h111;
rom[3945] = 12'h222;
rom[3946] = 12'h222;
rom[3947] = 12'h222;
rom[3948] = 12'h333;
rom[3949] = 12'h444;
rom[3950] = 12'h555;
rom[3951] = 12'h555;
rom[3952] = 12'h444;
rom[3953] = 12'h444;
rom[3954] = 12'h333;
rom[3955] = 12'h444;
rom[3956] = 12'h444;
rom[3957] = 12'h444;
rom[3958] = 12'h555;
rom[3959] = 12'h555;
rom[3960] = 12'h555;
rom[3961] = 12'h555;
rom[3962] = 12'h444;
rom[3963] = 12'h555;
rom[3964] = 12'h666;
rom[3965] = 12'h777;
rom[3966] = 12'h888;
rom[3967] = 12'h888;
rom[3968] = 12'h888;
rom[3969] = 12'h888;
rom[3970] = 12'h777;
rom[3971] = 12'h666;
rom[3972] = 12'h666;
rom[3973] = 12'h555;
rom[3974] = 12'h555;
rom[3975] = 12'h555;
rom[3976] = 12'h555;
rom[3977] = 12'h555;
rom[3978] = 12'h555;
rom[3979] = 12'h666;
rom[3980] = 12'h666;
rom[3981] = 12'h666;
rom[3982] = 12'h666;
rom[3983] = 12'h666;
rom[3984] = 12'h666;
rom[3985] = 12'h666;
rom[3986] = 12'h666;
rom[3987] = 12'h666;
rom[3988] = 12'h666;
rom[3989] = 12'h777;
rom[3990] = 12'h888;
rom[3991] = 12'h888;
rom[3992] = 12'h999;
rom[3993] = 12'h999;
rom[3994] = 12'h999;
rom[3995] = 12'h999;
rom[3996] = 12'h999;
rom[3997] = 12'h999;
rom[3998] = 12'h999;
rom[3999] = 12'h999;
rom[4000] = 12'h555;
rom[4001] = 12'h555;
rom[4002] = 12'h555;
rom[4003] = 12'h555;
rom[4004] = 12'h444;
rom[4005] = 12'h444;
rom[4006] = 12'h444;
rom[4007] = 12'h444;
rom[4008] = 12'h444;
rom[4009] = 12'h444;
rom[4010] = 12'h444;
rom[4011] = 12'h444;
rom[4012] = 12'h444;
rom[4013] = 12'h444;
rom[4014] = 12'h444;
rom[4015] = 12'h444;
rom[4016] = 12'h444;
rom[4017] = 12'h444;
rom[4018] = 12'h444;
rom[4019] = 12'h333;
rom[4020] = 12'h333;
rom[4021] = 12'h333;
rom[4022] = 12'h333;
rom[4023] = 12'h333;
rom[4024] = 12'h222;
rom[4025] = 12'h222;
rom[4026] = 12'h222;
rom[4027] = 12'h222;
rom[4028] = 12'h222;
rom[4029] = 12'h222;
rom[4030] = 12'h222;
rom[4031] = 12'h222;
rom[4032] = 12'h222;
rom[4033] = 12'h222;
rom[4034] = 12'h222;
rom[4035] = 12'h222;
rom[4036] = 12'h222;
rom[4037] = 12'h111;
rom[4038] = 12'h111;
rom[4039] = 12'h111;
rom[4040] = 12'h111;
rom[4041] = 12'h111;
rom[4042] = 12'h111;
rom[4043] = 12'h111;
rom[4044] = 12'h111;
rom[4045] = 12'h111;
rom[4046] = 12'h111;
rom[4047] = 12'h111;
rom[4048] = 12'h111;
rom[4049] = 12'h111;
rom[4050] = 12'h111;
rom[4051] = 12'h111;
rom[4052] = 12'h111;
rom[4053] = 12'h111;
rom[4054] = 12'h111;
rom[4055] = 12'h111;
rom[4056] = 12'h111;
rom[4057] = 12'h111;
rom[4058] = 12'h111;
rom[4059] = 12'h111;
rom[4060] = 12'h111;
rom[4061] = 12'h111;
rom[4062] = 12'h111;
rom[4063] = 12'h111;
rom[4064] = 12'h111;
rom[4065] = 12'h111;
rom[4066] = 12'h111;
rom[4067] = 12'h111;
rom[4068] = 12'h111;
rom[4069] = 12'h111;
rom[4070] = 12'h111;
rom[4071] = 12'h111;
rom[4072] = 12'h111;
rom[4073] = 12'h111;
rom[4074] = 12'h111;
rom[4075] = 12'h111;
rom[4076] = 12'h111;
rom[4077] = 12'h111;
rom[4078] = 12'h111;
rom[4079] = 12'h111;
rom[4080] = 12'h111;
rom[4081] = 12'h111;
rom[4082] = 12'h111;
rom[4083] = 12'h222;
rom[4084] = 12'h222;
rom[4085] = 12'h222;
rom[4086] = 12'h222;
rom[4087] = 12'h222;
rom[4088] = 12'h222;
rom[4089] = 12'h222;
rom[4090] = 12'h333;
rom[4091] = 12'h333;
rom[4092] = 12'h333;
rom[4093] = 12'h333;
rom[4094] = 12'h444;
rom[4095] = 12'h444;
rom[4096] = 12'h444;
rom[4097] = 12'h555;
rom[4098] = 12'h555;
rom[4099] = 12'h555;
rom[4100] = 12'h666;
rom[4101] = 12'h666;
rom[4102] = 12'h777;
rom[4103] = 12'h777;
rom[4104] = 12'h888;
rom[4105] = 12'h888;
rom[4106] = 12'h888;
rom[4107] = 12'h999;
rom[4108] = 12'h999;
rom[4109] = 12'haaa;
rom[4110] = 12'haaa;
rom[4111] = 12'hbbb;
rom[4112] = 12'hcbb;
rom[4113] = 12'hccc;
rom[4114] = 12'hdcc;
rom[4115] = 12'hddd;
rom[4116] = 12'hddd;
rom[4117] = 12'hddd;
rom[4118] = 12'hedd;
rom[4119] = 12'heed;
rom[4120] = 12'heed;
rom[4121] = 12'heed;
rom[4122] = 12'heed;
rom[4123] = 12'heed;
rom[4124] = 12'heed;
rom[4125] = 12'heed;
rom[4126] = 12'heee;
rom[4127] = 12'heee;
rom[4128] = 12'heee;
rom[4129] = 12'heed;
rom[4130] = 12'hded;
rom[4131] = 12'hddd;
rom[4132] = 12'hddd;
rom[4133] = 12'hddd;
rom[4134] = 12'hddc;
rom[4135] = 12'hcdc;
rom[4136] = 12'hccc;
rom[4137] = 12'hccc;
rom[4138] = 12'hccb;
rom[4139] = 12'hbcb;
rom[4140] = 12'hbbb;
rom[4141] = 12'hbbb;
rom[4142] = 12'hbcb;
rom[4143] = 12'hbcb;
rom[4144] = 12'hccc;
rom[4145] = 12'hbcc;
rom[4146] = 12'hbbb;
rom[4147] = 12'hbbb;
rom[4148] = 12'hbbb;
rom[4149] = 12'haab;
rom[4150] = 12'haaa;
rom[4151] = 12'h9aa;
rom[4152] = 12'h99a;
rom[4153] = 12'h999;
rom[4154] = 12'h999;
rom[4155] = 12'h899;
rom[4156] = 12'h899;
rom[4157] = 12'h888;
rom[4158] = 12'h888;
rom[4159] = 12'h888;
rom[4160] = 12'h999;
rom[4161] = 12'h998;
rom[4162] = 12'h888;
rom[4163] = 12'h888;
rom[4164] = 12'h888;
rom[4165] = 12'h888;
rom[4166] = 12'h777;
rom[4167] = 12'h777;
rom[4168] = 12'h777;
rom[4169] = 12'h666;
rom[4170] = 12'h666;
rom[4171] = 12'h666;
rom[4172] = 12'h776;
rom[4173] = 12'h777;
rom[4174] = 12'h666;
rom[4175] = 12'h666;
rom[4176] = 12'h555;
rom[4177] = 12'h555;
rom[4178] = 12'h444;
rom[4179] = 12'h444;
rom[4180] = 12'h555;
rom[4181] = 12'h555;
rom[4182] = 12'h555;
rom[4183] = 12'h444;
rom[4184] = 12'h555;
rom[4185] = 12'h555;
rom[4186] = 12'h555;
rom[4187] = 12'h444;
rom[4188] = 12'h444;
rom[4189] = 12'h444;
rom[4190] = 12'h555;
rom[4191] = 12'h555;
rom[4192] = 12'h666;
rom[4193] = 12'h666;
rom[4194] = 12'h666;
rom[4195] = 12'h555;
rom[4196] = 12'h666;
rom[4197] = 12'h777;
rom[4198] = 12'h777;
rom[4199] = 12'h888;
rom[4200] = 12'h888;
rom[4201] = 12'h777;
rom[4202] = 12'h777;
rom[4203] = 12'h666;
rom[4204] = 12'h444;
rom[4205] = 12'h444;
rom[4206] = 12'h444;
rom[4207] = 12'h333;
rom[4208] = 12'h222;
rom[4209] = 12'h222;
rom[4210] = 12'h222;
rom[4211] = 12'h222;
rom[4212] = 12'h222;
rom[4213] = 12'h222;
rom[4214] = 12'h222;
rom[4215] = 12'h222;
rom[4216] = 12'h222;
rom[4217] = 12'h222;
rom[4218] = 12'h  0;
rom[4219] = 12'h  0;
rom[4220] = 12'h  0;
rom[4221] = 12'h  0;
rom[4222] = 12'h  0;
rom[4223] = 12'h  0;
rom[4224] = 12'h  0;
rom[4225] = 12'h  0;
rom[4226] = 12'h  0;
rom[4227] = 12'h  0;
rom[4228] = 12'h  0;
rom[4229] = 12'h  0;
rom[4230] = 12'h  0;
rom[4231] = 12'h  0;
rom[4232] = 12'h  0;
rom[4233] = 12'h  0;
rom[4234] = 12'h  0;
rom[4235] = 12'h  0;
rom[4236] = 12'h  0;
rom[4237] = 12'h  0;
rom[4238] = 12'h  0;
rom[4239] = 12'h  0;
rom[4240] = 12'h  0;
rom[4241] = 12'h  0;
rom[4242] = 12'h  0;
rom[4243] = 12'h  0;
rom[4244] = 12'h  0;
rom[4245] = 12'h111;
rom[4246] = 12'h111;
rom[4247] = 12'h111;
rom[4248] = 12'h111;
rom[4249] = 12'h111;
rom[4250] = 12'h111;
rom[4251] = 12'h111;
rom[4252] = 12'h111;
rom[4253] = 12'h111;
rom[4254] = 12'h111;
rom[4255] = 12'h222;
rom[4256] = 12'h333;
rom[4257] = 12'h333;
rom[4258] = 12'h333;
rom[4259] = 12'h222;
rom[4260] = 12'h222;
rom[4261] = 12'h222;
rom[4262] = 12'h222;
rom[4263] = 12'h222;
rom[4264] = 12'h111;
rom[4265] = 12'h111;
rom[4266] = 12'h111;
rom[4267] = 12'h111;
rom[4268] = 12'h111;
rom[4269] = 12'h111;
rom[4270] = 12'h111;
rom[4271] = 12'h  0;
rom[4272] = 12'h  0;
rom[4273] = 12'h  0;
rom[4274] = 12'h  0;
rom[4275] = 12'h  0;
rom[4276] = 12'h  0;
rom[4277] = 12'h  0;
rom[4278] = 12'h  0;
rom[4279] = 12'h  0;
rom[4280] = 12'h  0;
rom[4281] = 12'h  0;
rom[4282] = 12'h  0;
rom[4283] = 12'h  0;
rom[4284] = 12'h  0;
rom[4285] = 12'h  0;
rom[4286] = 12'h  0;
rom[4287] = 12'h  0;
rom[4288] = 12'h  0;
rom[4289] = 12'h  0;
rom[4290] = 12'h  0;
rom[4291] = 12'h  0;
rom[4292] = 12'h  0;
rom[4293] = 12'h  0;
rom[4294] = 12'h  0;
rom[4295] = 12'h  0;
rom[4296] = 12'h  0;
rom[4297] = 12'h  0;
rom[4298] = 12'h  0;
rom[4299] = 12'h  0;
rom[4300] = 12'h111;
rom[4301] = 12'h111;
rom[4302] = 12'h111;
rom[4303] = 12'h111;
rom[4304] = 12'h  0;
rom[4305] = 12'h  0;
rom[4306] = 12'h  0;
rom[4307] = 12'h  0;
rom[4308] = 12'h  0;
rom[4309] = 12'h  0;
rom[4310] = 12'h  0;
rom[4311] = 12'h  0;
rom[4312] = 12'h  0;
rom[4313] = 12'h  0;
rom[4314] = 12'h  0;
rom[4315] = 12'h  0;
rom[4316] = 12'h  0;
rom[4317] = 12'h111;
rom[4318] = 12'h111;
rom[4319] = 12'h111;
rom[4320] = 12'h222;
rom[4321] = 12'h333;
rom[4322] = 12'h444;
rom[4323] = 12'h555;
rom[4324] = 12'h555;
rom[4325] = 12'h555;
rom[4326] = 12'h444;
rom[4327] = 12'h444;
rom[4328] = 12'h333;
rom[4329] = 12'h222;
rom[4330] = 12'h222;
rom[4331] = 12'h222;
rom[4332] = 12'h111;
rom[4333] = 12'h111;
rom[4334] = 12'h111;
rom[4335] = 12'h111;
rom[4336] = 12'h111;
rom[4337] = 12'h111;
rom[4338] = 12'h111;
rom[4339] = 12'h111;
rom[4340] = 12'h111;
rom[4341] = 12'h111;
rom[4342] = 12'h111;
rom[4343] = 12'h111;
rom[4344] = 12'h111;
rom[4345] = 12'h222;
rom[4346] = 12'h111;
rom[4347] = 12'h111;
rom[4348] = 12'h333;
rom[4349] = 12'h555;
rom[4350] = 12'h555;
rom[4351] = 12'h444;
rom[4352] = 12'h444;
rom[4353] = 12'h444;
rom[4354] = 12'h333;
rom[4355] = 12'h444;
rom[4356] = 12'h444;
rom[4357] = 12'h444;
rom[4358] = 12'h555;
rom[4359] = 12'h555;
rom[4360] = 12'h555;
rom[4361] = 12'h555;
rom[4362] = 12'h555;
rom[4363] = 12'h666;
rom[4364] = 12'h777;
rom[4365] = 12'h999;
rom[4366] = 12'h999;
rom[4367] = 12'h888;
rom[4368] = 12'h777;
rom[4369] = 12'h666;
rom[4370] = 12'h555;
rom[4371] = 12'h444;
rom[4372] = 12'h444;
rom[4373] = 12'h444;
rom[4374] = 12'h555;
rom[4375] = 12'h555;
rom[4376] = 12'h555;
rom[4377] = 12'h555;
rom[4378] = 12'h555;
rom[4379] = 12'h555;
rom[4380] = 12'h555;
rom[4381] = 12'h666;
rom[4382] = 12'h666;
rom[4383] = 12'h666;
rom[4384] = 12'h666;
rom[4385] = 12'h666;
rom[4386] = 12'h666;
rom[4387] = 12'h666;
rom[4388] = 12'h666;
rom[4389] = 12'h777;
rom[4390] = 12'h888;
rom[4391] = 12'h888;
rom[4392] = 12'h999;
rom[4393] = 12'h999;
rom[4394] = 12'h999;
rom[4395] = 12'h999;
rom[4396] = 12'h999;
rom[4397] = 12'h999;
rom[4398] = 12'h999;
rom[4399] = 12'h999;
rom[4400] = 12'h555;
rom[4401] = 12'h555;
rom[4402] = 12'h555;
rom[4403] = 12'h555;
rom[4404] = 12'h555;
rom[4405] = 12'h555;
rom[4406] = 12'h444;
rom[4407] = 12'h444;
rom[4408] = 12'h444;
rom[4409] = 12'h444;
rom[4410] = 12'h444;
rom[4411] = 12'h444;
rom[4412] = 12'h444;
rom[4413] = 12'h444;
rom[4414] = 12'h444;
rom[4415] = 12'h444;
rom[4416] = 12'h444;
rom[4417] = 12'h444;
rom[4418] = 12'h333;
rom[4419] = 12'h333;
rom[4420] = 12'h333;
rom[4421] = 12'h222;
rom[4422] = 12'h222;
rom[4423] = 12'h222;
rom[4424] = 12'h222;
rom[4425] = 12'h222;
rom[4426] = 12'h222;
rom[4427] = 12'h111;
rom[4428] = 12'h111;
rom[4429] = 12'h111;
rom[4430] = 12'h111;
rom[4431] = 12'h222;
rom[4432] = 12'h111;
rom[4433] = 12'h111;
rom[4434] = 12'h111;
rom[4435] = 12'h111;
rom[4436] = 12'h111;
rom[4437] = 12'h111;
rom[4438] = 12'h111;
rom[4439] = 12'h111;
rom[4440] = 12'h111;
rom[4441] = 12'h111;
rom[4442] = 12'h111;
rom[4443] = 12'h111;
rom[4444] = 12'h111;
rom[4445] = 12'h111;
rom[4446] = 12'h  0;
rom[4447] = 12'h  0;
rom[4448] = 12'h  0;
rom[4449] = 12'h  0;
rom[4450] = 12'h  0;
rom[4451] = 12'h  0;
rom[4452] = 12'h  0;
rom[4453] = 12'h  0;
rom[4454] = 12'h111;
rom[4455] = 12'h111;
rom[4456] = 12'h111;
rom[4457] = 12'h111;
rom[4458] = 12'h111;
rom[4459] = 12'h111;
rom[4460] = 12'h111;
rom[4461] = 12'h111;
rom[4462] = 12'h111;
rom[4463] = 12'h111;
rom[4464] = 12'h111;
rom[4465] = 12'h111;
rom[4466] = 12'h111;
rom[4467] = 12'h111;
rom[4468] = 12'h111;
rom[4469] = 12'h111;
rom[4470] = 12'h111;
rom[4471] = 12'h111;
rom[4472] = 12'h111;
rom[4473] = 12'h111;
rom[4474] = 12'h111;
rom[4475] = 12'h111;
rom[4476] = 12'h111;
rom[4477] = 12'h111;
rom[4478] = 12'h111;
rom[4479] = 12'h111;
rom[4480] = 12'h111;
rom[4481] = 12'h111;
rom[4482] = 12'h111;
rom[4483] = 12'h111;
rom[4484] = 12'h111;
rom[4485] = 12'h111;
rom[4486] = 12'h111;
rom[4487] = 12'h111;
rom[4488] = 12'h111;
rom[4489] = 12'h111;
rom[4490] = 12'h222;
rom[4491] = 12'h222;
rom[4492] = 12'h222;
rom[4493] = 12'h333;
rom[4494] = 12'h333;
rom[4495] = 12'h333;
rom[4496] = 12'h444;
rom[4497] = 12'h444;
rom[4498] = 12'h555;
rom[4499] = 12'h555;
rom[4500] = 12'h555;
rom[4501] = 12'h555;
rom[4502] = 12'h666;
rom[4503] = 12'h777;
rom[4504] = 12'h777;
rom[4505] = 12'h777;
rom[4506] = 12'h888;
rom[4507] = 12'h999;
rom[4508] = 12'h999;
rom[4509] = 12'haaa;
rom[4510] = 12'hbbb;
rom[4511] = 12'hccc;
rom[4512] = 12'hdcc;
rom[4513] = 12'hddc;
rom[4514] = 12'heed;
rom[4515] = 12'heed;
rom[4516] = 12'heed;
rom[4517] = 12'heed;
rom[4518] = 12'heed;
rom[4519] = 12'heed;
rom[4520] = 12'hfed;
rom[4521] = 12'hfed;
rom[4522] = 12'hfed;
rom[4523] = 12'hfed;
rom[4524] = 12'hfed;
rom[4525] = 12'hfed;
rom[4526] = 12'hfed;
rom[4527] = 12'heed;
rom[4528] = 12'hddc;
rom[4529] = 12'hddc;
rom[4530] = 12'hddc;
rom[4531] = 12'hcdc;
rom[4532] = 12'hccc;
rom[4533] = 12'hccc;
rom[4534] = 12'hccc;
rom[4535] = 12'hccc;
rom[4536] = 12'hccb;
rom[4537] = 12'hbbb;
rom[4538] = 12'hbbb;
rom[4539] = 12'hbba;
rom[4540] = 12'hbba;
rom[4541] = 12'hbba;
rom[4542] = 12'hbba;
rom[4543] = 12'hbba;
rom[4544] = 12'hbba;
rom[4545] = 12'hbbb;
rom[4546] = 12'hbbb;
rom[4547] = 12'hbbb;
rom[4548] = 12'hbbb;
rom[4549] = 12'hbbb;
rom[4550] = 12'hbbb;
rom[4551] = 12'hbbb;
rom[4552] = 12'hbbb;
rom[4553] = 12'habb;
rom[4554] = 12'haaa;
rom[4555] = 12'h9aa;
rom[4556] = 12'h999;
rom[4557] = 12'h999;
rom[4558] = 12'h888;
rom[4559] = 12'h888;
rom[4560] = 12'h888;
rom[4561] = 12'h888;
rom[4562] = 12'h999;
rom[4563] = 12'h999;
rom[4564] = 12'h999;
rom[4565] = 12'h999;
rom[4566] = 12'h999;
rom[4567] = 12'h898;
rom[4568] = 12'h777;
rom[4569] = 12'h777;
rom[4570] = 12'h666;
rom[4571] = 12'h666;
rom[4572] = 12'h776;
rom[4573] = 12'h777;
rom[4574] = 12'h777;
rom[4575] = 12'h777;
rom[4576] = 12'h666;
rom[4577] = 12'h555;
rom[4578] = 12'h555;
rom[4579] = 12'h444;
rom[4580] = 12'h444;
rom[4581] = 12'h444;
rom[4582] = 12'h444;
rom[4583] = 12'h444;
rom[4584] = 12'h555;
rom[4585] = 12'h555;
rom[4586] = 12'h555;
rom[4587] = 12'h555;
rom[4588] = 12'h555;
rom[4589] = 12'h444;
rom[4590] = 12'h444;
rom[4591] = 12'h555;
rom[4592] = 12'h555;
rom[4593] = 12'h666;
rom[4594] = 12'h666;
rom[4595] = 12'h666;
rom[4596] = 12'h666;
rom[4597] = 12'h777;
rom[4598] = 12'h888;
rom[4599] = 12'h888;
rom[4600] = 12'h777;
rom[4601] = 12'h777;
rom[4602] = 12'h777;
rom[4603] = 12'h666;
rom[4604] = 12'h444;
rom[4605] = 12'h555;
rom[4606] = 12'h444;
rom[4607] = 12'h333;
rom[4608] = 12'h222;
rom[4609] = 12'h222;
rom[4610] = 12'h222;
rom[4611] = 12'h222;
rom[4612] = 12'h222;
rom[4613] = 12'h222;
rom[4614] = 12'h222;
rom[4615] = 12'h333;
rom[4616] = 12'h222;
rom[4617] = 12'h111;
rom[4618] = 12'h  0;
rom[4619] = 12'h  0;
rom[4620] = 12'h  0;
rom[4621] = 12'h  0;
rom[4622] = 12'h  0;
rom[4623] = 12'h  0;
rom[4624] = 12'h  0;
rom[4625] = 12'h  0;
rom[4626] = 12'h  0;
rom[4627] = 12'h  0;
rom[4628] = 12'h  0;
rom[4629] = 12'h  0;
rom[4630] = 12'h  0;
rom[4631] = 12'h  0;
rom[4632] = 12'h  0;
rom[4633] = 12'h  0;
rom[4634] = 12'h  0;
rom[4635] = 12'h  0;
rom[4636] = 12'h  0;
rom[4637] = 12'h  0;
rom[4638] = 12'h  0;
rom[4639] = 12'h  0;
rom[4640] = 12'h  0;
rom[4641] = 12'h  0;
rom[4642] = 12'h  0;
rom[4643] = 12'h  0;
rom[4644] = 12'h  0;
rom[4645] = 12'h111;
rom[4646] = 12'h111;
rom[4647] = 12'h111;
rom[4648] = 12'h111;
rom[4649] = 12'h111;
rom[4650] = 12'h111;
rom[4651] = 12'h111;
rom[4652] = 12'h111;
rom[4653] = 12'h111;
rom[4654] = 12'h222;
rom[4655] = 12'h222;
rom[4656] = 12'h333;
rom[4657] = 12'h333;
rom[4658] = 12'h222;
rom[4659] = 12'h222;
rom[4660] = 12'h222;
rom[4661] = 12'h222;
rom[4662] = 12'h222;
rom[4663] = 12'h111;
rom[4664] = 12'h111;
rom[4665] = 12'h111;
rom[4666] = 12'h111;
rom[4667] = 12'h111;
rom[4668] = 12'h111;
rom[4669] = 12'h111;
rom[4670] = 12'h111;
rom[4671] = 12'h  0;
rom[4672] = 12'h  0;
rom[4673] = 12'h  0;
rom[4674] = 12'h  0;
rom[4675] = 12'h  0;
rom[4676] = 12'h  0;
rom[4677] = 12'h  0;
rom[4678] = 12'h  0;
rom[4679] = 12'h  0;
rom[4680] = 12'h  0;
rom[4681] = 12'h  0;
rom[4682] = 12'h  0;
rom[4683] = 12'h  0;
rom[4684] = 12'h  0;
rom[4685] = 12'h  0;
rom[4686] = 12'h  0;
rom[4687] = 12'h  0;
rom[4688] = 12'h  0;
rom[4689] = 12'h  0;
rom[4690] = 12'h  0;
rom[4691] = 12'h  0;
rom[4692] = 12'h  0;
rom[4693] = 12'h  0;
rom[4694] = 12'h  0;
rom[4695] = 12'h  0;
rom[4696] = 12'h  0;
rom[4697] = 12'h  0;
rom[4698] = 12'h  0;
rom[4699] = 12'h  0;
rom[4700] = 12'h111;
rom[4701] = 12'h111;
rom[4702] = 12'h111;
rom[4703] = 12'h111;
rom[4704] = 12'h  0;
rom[4705] = 12'h  0;
rom[4706] = 12'h  0;
rom[4707] = 12'h  0;
rom[4708] = 12'h  0;
rom[4709] = 12'h  0;
rom[4710] = 12'h  0;
rom[4711] = 12'h  0;
rom[4712] = 12'h  0;
rom[4713] = 12'h  0;
rom[4714] = 12'h  0;
rom[4715] = 12'h  0;
rom[4716] = 12'h  0;
rom[4717] = 12'h111;
rom[4718] = 12'h111;
rom[4719] = 12'h111;
rom[4720] = 12'h222;
rom[4721] = 12'h444;
rom[4722] = 12'h555;
rom[4723] = 12'h555;
rom[4724] = 12'h555;
rom[4725] = 12'h555;
rom[4726] = 12'h555;
rom[4727] = 12'h444;
rom[4728] = 12'h222;
rom[4729] = 12'h222;
rom[4730] = 12'h222;
rom[4731] = 12'h222;
rom[4732] = 12'h111;
rom[4733] = 12'h111;
rom[4734] = 12'h111;
rom[4735] = 12'h111;
rom[4736] = 12'h111;
rom[4737] = 12'h111;
rom[4738] = 12'h111;
rom[4739] = 12'h111;
rom[4740] = 12'h111;
rom[4741] = 12'h111;
rom[4742] = 12'h111;
rom[4743] = 12'h111;
rom[4744] = 12'h111;
rom[4745] = 12'h111;
rom[4746] = 12'h111;
rom[4747] = 12'h222;
rom[4748] = 12'h444;
rom[4749] = 12'h555;
rom[4750] = 12'h555;
rom[4751] = 12'h444;
rom[4752] = 12'h444;
rom[4753] = 12'h444;
rom[4754] = 12'h444;
rom[4755] = 12'h444;
rom[4756] = 12'h444;
rom[4757] = 12'h444;
rom[4758] = 12'h444;
rom[4759] = 12'h555;
rom[4760] = 12'h555;
rom[4761] = 12'h555;
rom[4762] = 12'h666;
rom[4763] = 12'h888;
rom[4764] = 12'h999;
rom[4765] = 12'h999;
rom[4766] = 12'h888;
rom[4767] = 12'h777;
rom[4768] = 12'h555;
rom[4769] = 12'h555;
rom[4770] = 12'h444;
rom[4771] = 12'h444;
rom[4772] = 12'h444;
rom[4773] = 12'h444;
rom[4774] = 12'h444;
rom[4775] = 12'h444;
rom[4776] = 12'h444;
rom[4777] = 12'h444;
rom[4778] = 12'h555;
rom[4779] = 12'h555;
rom[4780] = 12'h555;
rom[4781] = 12'h555;
rom[4782] = 12'h666;
rom[4783] = 12'h666;
rom[4784] = 12'h666;
rom[4785] = 12'h666;
rom[4786] = 12'h666;
rom[4787] = 12'h666;
rom[4788] = 12'h666;
rom[4789] = 12'h777;
rom[4790] = 12'h777;
rom[4791] = 12'h888;
rom[4792] = 12'h999;
rom[4793] = 12'h999;
rom[4794] = 12'h999;
rom[4795] = 12'h999;
rom[4796] = 12'h999;
rom[4797] = 12'h999;
rom[4798] = 12'h999;
rom[4799] = 12'h999;
rom[4800] = 12'h555;
rom[4801] = 12'h555;
rom[4802] = 12'h555;
rom[4803] = 12'h444;
rom[4804] = 12'h444;
rom[4805] = 12'h444;
rom[4806] = 12'h444;
rom[4807] = 12'h444;
rom[4808] = 12'h555;
rom[4809] = 12'h444;
rom[4810] = 12'h444;
rom[4811] = 12'h444;
rom[4812] = 12'h444;
rom[4813] = 12'h444;
rom[4814] = 12'h444;
rom[4815] = 12'h444;
rom[4816] = 12'h444;
rom[4817] = 12'h333;
rom[4818] = 12'h333;
rom[4819] = 12'h333;
rom[4820] = 12'h222;
rom[4821] = 12'h222;
rom[4822] = 12'h222;
rom[4823] = 12'h222;
rom[4824] = 12'h222;
rom[4825] = 12'h111;
rom[4826] = 12'h111;
rom[4827] = 12'h111;
rom[4828] = 12'h111;
rom[4829] = 12'h111;
rom[4830] = 12'h111;
rom[4831] = 12'h111;
rom[4832] = 12'h111;
rom[4833] = 12'h111;
rom[4834] = 12'h111;
rom[4835] = 12'h111;
rom[4836] = 12'h111;
rom[4837] = 12'h111;
rom[4838] = 12'h111;
rom[4839] = 12'h111;
rom[4840] = 12'h111;
rom[4841] = 12'h111;
rom[4842] = 12'h111;
rom[4843] = 12'h111;
rom[4844] = 12'h111;
rom[4845] = 12'h  0;
rom[4846] = 12'h  0;
rom[4847] = 12'h  0;
rom[4848] = 12'h  0;
rom[4849] = 12'h  0;
rom[4850] = 12'h  0;
rom[4851] = 12'h  0;
rom[4852] = 12'h  0;
rom[4853] = 12'h  0;
rom[4854] = 12'h  0;
rom[4855] = 12'h111;
rom[4856] = 12'h  0;
rom[4857] = 12'h  0;
rom[4858] = 12'h  0;
rom[4859] = 12'h111;
rom[4860] = 12'h111;
rom[4861] = 12'h111;
rom[4862] = 12'h111;
rom[4863] = 12'h111;
rom[4864] = 12'h111;
rom[4865] = 12'h111;
rom[4866] = 12'h111;
rom[4867] = 12'h111;
rom[4868] = 12'h111;
rom[4869] = 12'h111;
rom[4870] = 12'h111;
rom[4871] = 12'h111;
rom[4872] = 12'h111;
rom[4873] = 12'h111;
rom[4874] = 12'h111;
rom[4875] = 12'h111;
rom[4876] = 12'h111;
rom[4877] = 12'h111;
rom[4878] = 12'h111;
rom[4879] = 12'h111;
rom[4880] = 12'h111;
rom[4881] = 12'h111;
rom[4882] = 12'h111;
rom[4883] = 12'h111;
rom[4884] = 12'h111;
rom[4885] = 12'h111;
rom[4886] = 12'h111;
rom[4887] = 12'h111;
rom[4888] = 12'h111;
rom[4889] = 12'h111;
rom[4890] = 12'h111;
rom[4891] = 12'h111;
rom[4892] = 12'h222;
rom[4893] = 12'h222;
rom[4894] = 12'h222;
rom[4895] = 12'h333;
rom[4896] = 12'h333;
rom[4897] = 12'h444;
rom[4898] = 12'h444;
rom[4899] = 12'h444;
rom[4900] = 12'h555;
rom[4901] = 12'h555;
rom[4902] = 12'h666;
rom[4903] = 12'h777;
rom[4904] = 12'h888;
rom[4905] = 12'h999;
rom[4906] = 12'haaa;
rom[4907] = 12'haaa;
rom[4908] = 12'hbbb;
rom[4909] = 12'hbbb;
rom[4910] = 12'hccc;
rom[4911] = 12'hccc;
rom[4912] = 12'hdcc;
rom[4913] = 12'hedc;
rom[4914] = 12'hedc;
rom[4915] = 12'hedc;
rom[4916] = 12'hedc;
rom[4917] = 12'hedc;
rom[4918] = 12'hedc;
rom[4919] = 12'hedc;
rom[4920] = 12'hedc;
rom[4921] = 12'hedc;
rom[4922] = 12'hedc;
rom[4923] = 12'hedc;
rom[4924] = 12'hecb;
rom[4925] = 12'hdcb;
rom[4926] = 12'hdbb;
rom[4927] = 12'hcbb;
rom[4928] = 12'hbba;
rom[4929] = 12'hbba;
rom[4930] = 12'hbba;
rom[4931] = 12'hbba;
rom[4932] = 12'hbba;
rom[4933] = 12'hbba;
rom[4934] = 12'hbba;
rom[4935] = 12'hbba;
rom[4936] = 12'hbaa;
rom[4937] = 12'hbaa;
rom[4938] = 12'hbaa;
rom[4939] = 12'hbaa;
rom[4940] = 12'hbaa;
rom[4941] = 12'haaa;
rom[4942] = 12'haa9;
rom[4943] = 12'haa9;
rom[4944] = 12'haa9;
rom[4945] = 12'haa9;
rom[4946] = 12'haa9;
rom[4947] = 12'hbaa;
rom[4948] = 12'hbaa;
rom[4949] = 12'hbaa;
rom[4950] = 12'hbba;
rom[4951] = 12'hbba;
rom[4952] = 12'hbba;
rom[4953] = 12'hbba;
rom[4954] = 12'hbba;
rom[4955] = 12'hbaa;
rom[4956] = 12'haaa;
rom[4957] = 12'haaa;
rom[4958] = 12'haaa;
rom[4959] = 12'haaa;
rom[4960] = 12'h999;
rom[4961] = 12'h999;
rom[4962] = 12'h999;
rom[4963] = 12'h999;
rom[4964] = 12'h999;
rom[4965] = 12'h999;
rom[4966] = 12'h999;
rom[4967] = 12'h999;
rom[4968] = 12'h888;
rom[4969] = 12'h888;
rom[4970] = 12'h887;
rom[4971] = 12'h777;
rom[4972] = 12'h777;
rom[4973] = 12'h776;
rom[4974] = 12'h777;
rom[4975] = 12'h777;
rom[4976] = 12'h777;
rom[4977] = 12'h666;
rom[4978] = 12'h666;
rom[4979] = 12'h555;
rom[4980] = 12'h555;
rom[4981] = 12'h555;
rom[4982] = 12'h555;
rom[4983] = 12'h555;
rom[4984] = 12'h555;
rom[4985] = 12'h555;
rom[4986] = 12'h555;
rom[4987] = 12'h555;
rom[4988] = 12'h555;
rom[4989] = 12'h555;
rom[4990] = 12'h555;
rom[4991] = 12'h555;
rom[4992] = 12'h555;
rom[4993] = 12'h666;
rom[4994] = 12'h666;
rom[4995] = 12'h666;
rom[4996] = 12'h666;
rom[4997] = 12'h777;
rom[4998] = 12'h888;
rom[4999] = 12'h888;
rom[5000] = 12'h777;
rom[5001] = 12'h777;
rom[5002] = 12'h777;
rom[5003] = 12'h666;
rom[5004] = 12'h444;
rom[5005] = 12'h444;
rom[5006] = 12'h444;
rom[5007] = 12'h333;
rom[5008] = 12'h222;
rom[5009] = 12'h222;
rom[5010] = 12'h222;
rom[5011] = 12'h222;
rom[5012] = 12'h222;
rom[5013] = 12'h222;
rom[5014] = 12'h333;
rom[5015] = 12'h333;
rom[5016] = 12'h222;
rom[5017] = 12'h111;
rom[5018] = 12'h  0;
rom[5019] = 12'h  0;
rom[5020] = 12'h  0;
rom[5021] = 12'h  0;
rom[5022] = 12'h  0;
rom[5023] = 12'h  0;
rom[5024] = 12'h  0;
rom[5025] = 12'h  0;
rom[5026] = 12'h  0;
rom[5027] = 12'h  0;
rom[5028] = 12'h  0;
rom[5029] = 12'h  0;
rom[5030] = 12'h  0;
rom[5031] = 12'h  0;
rom[5032] = 12'h  0;
rom[5033] = 12'h  0;
rom[5034] = 12'h  0;
rom[5035] = 12'h  0;
rom[5036] = 12'h  0;
rom[5037] = 12'h  0;
rom[5038] = 12'h  0;
rom[5039] = 12'h  0;
rom[5040] = 12'h  0;
rom[5041] = 12'h  0;
rom[5042] = 12'h  0;
rom[5043] = 12'h  0;
rom[5044] = 12'h111;
rom[5045] = 12'h111;
rom[5046] = 12'h111;
rom[5047] = 12'h111;
rom[5048] = 12'h222;
rom[5049] = 12'h111;
rom[5050] = 12'h111;
rom[5051] = 12'h111;
rom[5052] = 12'h111;
rom[5053] = 12'h222;
rom[5054] = 12'h222;
rom[5055] = 12'h333;
rom[5056] = 12'h333;
rom[5057] = 12'h222;
rom[5058] = 12'h222;
rom[5059] = 12'h111;
rom[5060] = 12'h222;
rom[5061] = 12'h222;
rom[5062] = 12'h222;
rom[5063] = 12'h111;
rom[5064] = 12'h111;
rom[5065] = 12'h111;
rom[5066] = 12'h111;
rom[5067] = 12'h111;
rom[5068] = 12'h111;
rom[5069] = 12'h111;
rom[5070] = 12'h  0;
rom[5071] = 12'h  0;
rom[5072] = 12'h  0;
rom[5073] = 12'h  0;
rom[5074] = 12'h  0;
rom[5075] = 12'h  0;
rom[5076] = 12'h  0;
rom[5077] = 12'h  0;
rom[5078] = 12'h  0;
rom[5079] = 12'h  0;
rom[5080] = 12'h  0;
rom[5081] = 12'h  0;
rom[5082] = 12'h  0;
rom[5083] = 12'h  0;
rom[5084] = 12'h  0;
rom[5085] = 12'h  0;
rom[5086] = 12'h  0;
rom[5087] = 12'h  0;
rom[5088] = 12'h  0;
rom[5089] = 12'h  0;
rom[5090] = 12'h  0;
rom[5091] = 12'h  0;
rom[5092] = 12'h  0;
rom[5093] = 12'h  0;
rom[5094] = 12'h  0;
rom[5095] = 12'h  0;
rom[5096] = 12'h  0;
rom[5097] = 12'h  0;
rom[5098] = 12'h  0;
rom[5099] = 12'h  0;
rom[5100] = 12'h  0;
rom[5101] = 12'h111;
rom[5102] = 12'h111;
rom[5103] = 12'h  0;
rom[5104] = 12'h  0;
rom[5105] = 12'h  0;
rom[5106] = 12'h  0;
rom[5107] = 12'h  0;
rom[5108] = 12'h  0;
rom[5109] = 12'h  0;
rom[5110] = 12'h  0;
rom[5111] = 12'h  0;
rom[5112] = 12'h  0;
rom[5113] = 12'h  0;
rom[5114] = 12'h  0;
rom[5115] = 12'h  0;
rom[5116] = 12'h  0;
rom[5117] = 12'h  0;
rom[5118] = 12'h111;
rom[5119] = 12'h111;
rom[5120] = 12'h222;
rom[5121] = 12'h444;
rom[5122] = 12'h555;
rom[5123] = 12'h555;
rom[5124] = 12'h555;
rom[5125] = 12'h555;
rom[5126] = 12'h555;
rom[5127] = 12'h444;
rom[5128] = 12'h222;
rom[5129] = 12'h222;
rom[5130] = 12'h222;
rom[5131] = 12'h222;
rom[5132] = 12'h111;
rom[5133] = 12'h111;
rom[5134] = 12'h111;
rom[5135] = 12'h111;
rom[5136] = 12'h111;
rom[5137] = 12'h111;
rom[5138] = 12'h111;
rom[5139] = 12'h111;
rom[5140] = 12'h111;
rom[5141] = 12'h111;
rom[5142] = 12'h111;
rom[5143] = 12'h222;
rom[5144] = 12'h111;
rom[5145] = 12'h111;
rom[5146] = 12'h222;
rom[5147] = 12'h444;
rom[5148] = 12'h444;
rom[5149] = 12'h444;
rom[5150] = 12'h444;
rom[5151] = 12'h333;
rom[5152] = 12'h444;
rom[5153] = 12'h444;
rom[5154] = 12'h444;
rom[5155] = 12'h444;
rom[5156] = 12'h444;
rom[5157] = 12'h444;
rom[5158] = 12'h444;
rom[5159] = 12'h555;
rom[5160] = 12'h555;
rom[5161] = 12'h777;
rom[5162] = 12'h888;
rom[5163] = 12'h999;
rom[5164] = 12'h888;
rom[5165] = 12'h777;
rom[5166] = 12'h555;
rom[5167] = 12'h444;
rom[5168] = 12'h444;
rom[5169] = 12'h444;
rom[5170] = 12'h444;
rom[5171] = 12'h444;
rom[5172] = 12'h444;
rom[5173] = 12'h444;
rom[5174] = 12'h444;
rom[5175] = 12'h444;
rom[5176] = 12'h444;
rom[5177] = 12'h555;
rom[5178] = 12'h555;
rom[5179] = 12'h555;
rom[5180] = 12'h555;
rom[5181] = 12'h555;
rom[5182] = 12'h666;
rom[5183] = 12'h666;
rom[5184] = 12'h666;
rom[5185] = 12'h666;
rom[5186] = 12'h666;
rom[5187] = 12'h666;
rom[5188] = 12'h666;
rom[5189] = 12'h777;
rom[5190] = 12'h777;
rom[5191] = 12'h888;
rom[5192] = 12'h999;
rom[5193] = 12'h999;
rom[5194] = 12'h999;
rom[5195] = 12'h999;
rom[5196] = 12'h999;
rom[5197] = 12'h999;
rom[5198] = 12'h999;
rom[5199] = 12'h999;
rom[5200] = 12'h444;
rom[5201] = 12'h444;
rom[5202] = 12'h444;
rom[5203] = 12'h444;
rom[5204] = 12'h444;
rom[5205] = 12'h444;
rom[5206] = 12'h444;
rom[5207] = 12'h444;
rom[5208] = 12'h555;
rom[5209] = 12'h555;
rom[5210] = 12'h555;
rom[5211] = 12'h444;
rom[5212] = 12'h444;
rom[5213] = 12'h444;
rom[5214] = 12'h444;
rom[5215] = 12'h333;
rom[5216] = 12'h333;
rom[5217] = 12'h333;
rom[5218] = 12'h333;
rom[5219] = 12'h222;
rom[5220] = 12'h222;
rom[5221] = 12'h222;
rom[5222] = 12'h222;
rom[5223] = 12'h111;
rom[5224] = 12'h111;
rom[5225] = 12'h111;
rom[5226] = 12'h111;
rom[5227] = 12'h111;
rom[5228] = 12'h111;
rom[5229] = 12'h111;
rom[5230] = 12'h111;
rom[5231] = 12'h111;
rom[5232] = 12'h111;
rom[5233] = 12'h111;
rom[5234] = 12'h111;
rom[5235] = 12'h111;
rom[5236] = 12'h111;
rom[5237] = 12'h111;
rom[5238] = 12'h111;
rom[5239] = 12'h111;
rom[5240] = 12'h111;
rom[5241] = 12'h111;
rom[5242] = 12'h111;
rom[5243] = 12'h111;
rom[5244] = 12'h  0;
rom[5245] = 12'h  0;
rom[5246] = 12'h  0;
rom[5247] = 12'h  0;
rom[5248] = 12'h  0;
rom[5249] = 12'h  0;
rom[5250] = 12'h  0;
rom[5251] = 12'h  0;
rom[5252] = 12'h  0;
rom[5253] = 12'h  0;
rom[5254] = 12'h  0;
rom[5255] = 12'h  0;
rom[5256] = 12'h  0;
rom[5257] = 12'h  0;
rom[5258] = 12'h  0;
rom[5259] = 12'h  0;
rom[5260] = 12'h111;
rom[5261] = 12'h111;
rom[5262] = 12'h111;
rom[5263] = 12'h111;
rom[5264] = 12'h111;
rom[5265] = 12'h111;
rom[5266] = 12'h111;
rom[5267] = 12'h111;
rom[5268] = 12'h111;
rom[5269] = 12'h111;
rom[5270] = 12'h111;
rom[5271] = 12'h111;
rom[5272] = 12'h111;
rom[5273] = 12'h111;
rom[5274] = 12'h111;
rom[5275] = 12'h  0;
rom[5276] = 12'h  0;
rom[5277] = 12'h111;
rom[5278] = 12'h111;
rom[5279] = 12'h111;
rom[5280] = 12'h111;
rom[5281] = 12'h111;
rom[5282] = 12'h111;
rom[5283] = 12'h111;
rom[5284] = 12'h111;
rom[5285] = 12'h111;
rom[5286] = 12'h111;
rom[5287] = 12'h111;
rom[5288] = 12'h  0;
rom[5289] = 12'h111;
rom[5290] = 12'h111;
rom[5291] = 12'h111;
rom[5292] = 12'h222;
rom[5293] = 12'h222;
rom[5294] = 12'h222;
rom[5295] = 12'h333;
rom[5296] = 12'h444;
rom[5297] = 12'h444;
rom[5298] = 12'h555;
rom[5299] = 12'h555;
rom[5300] = 12'h666;
rom[5301] = 12'h666;
rom[5302] = 12'h777;
rom[5303] = 12'h888;
rom[5304] = 12'h999;
rom[5305] = 12'haaa;
rom[5306] = 12'haaa;
rom[5307] = 12'haaa;
rom[5308] = 12'haaa;
rom[5309] = 12'haaa;
rom[5310] = 12'haaa;
rom[5311] = 12'hbba;
rom[5312] = 12'hbba;
rom[5313] = 12'hcba;
rom[5314] = 12'hcba;
rom[5315] = 12'hcba;
rom[5316] = 12'hcba;
rom[5317] = 12'hcb9;
rom[5318] = 12'hcb9;
rom[5319] = 12'hcb9;
rom[5320] = 12'hcb9;
rom[5321] = 12'hcb9;
rom[5322] = 12'hcb9;
rom[5323] = 12'hca9;
rom[5324] = 12'hba8;
rom[5325] = 12'hb98;
rom[5326] = 12'ha87;
rom[5327] = 12'ha87;
rom[5328] = 12'ha98;
rom[5329] = 12'h998;
rom[5330] = 12'h998;
rom[5331] = 12'h998;
rom[5332] = 12'h998;
rom[5333] = 12'h998;
rom[5334] = 12'ha98;
rom[5335] = 12'ha98;
rom[5336] = 12'h998;
rom[5337] = 12'ha98;
rom[5338] = 12'ha98;
rom[5339] = 12'ha98;
rom[5340] = 12'ha99;
rom[5341] = 12'ha99;
rom[5342] = 12'ha99;
rom[5343] = 12'ha99;
rom[5344] = 12'ha99;
rom[5345] = 12'haa9;
rom[5346] = 12'hba9;
rom[5347] = 12'hba9;
rom[5348] = 12'hba9;
rom[5349] = 12'haa9;
rom[5350] = 12'hba9;
rom[5351] = 12'hba9;
rom[5352] = 12'hbaa;
rom[5353] = 12'hbaa;
rom[5354] = 12'hbaa;
rom[5355] = 12'hbba;
rom[5356] = 12'hbba;
rom[5357] = 12'hbba;
rom[5358] = 12'hbba;
rom[5359] = 12'hbba;
rom[5360] = 12'haaa;
rom[5361] = 12'haaa;
rom[5362] = 12'haaa;
rom[5363] = 12'haaa;
rom[5364] = 12'haaa;
rom[5365] = 12'haaa;
rom[5366] = 12'haa9;
rom[5367] = 12'h9a9;
rom[5368] = 12'h999;
rom[5369] = 12'h999;
rom[5370] = 12'h999;
rom[5371] = 12'h888;
rom[5372] = 12'h787;
rom[5373] = 12'h777;
rom[5374] = 12'h776;
rom[5375] = 12'h777;
rom[5376] = 12'h777;
rom[5377] = 12'h777;
rom[5378] = 12'h777;
rom[5379] = 12'h666;
rom[5380] = 12'h666;
rom[5381] = 12'h555;
rom[5382] = 12'h555;
rom[5383] = 12'h555;
rom[5384] = 12'h555;
rom[5385] = 12'h555;
rom[5386] = 12'h555;
rom[5387] = 12'h555;
rom[5388] = 12'h555;
rom[5389] = 12'h555;
rom[5390] = 12'h555;
rom[5391] = 12'h555;
rom[5392] = 12'h555;
rom[5393] = 12'h555;
rom[5394] = 12'h666;
rom[5395] = 12'h666;
rom[5396] = 12'h666;
rom[5397] = 12'h777;
rom[5398] = 12'h888;
rom[5399] = 12'h777;
rom[5400] = 12'h777;
rom[5401] = 12'h777;
rom[5402] = 12'h777;
rom[5403] = 12'h666;
rom[5404] = 12'h555;
rom[5405] = 12'h444;
rom[5406] = 12'h444;
rom[5407] = 12'h333;
rom[5408] = 12'h333;
rom[5409] = 12'h333;
rom[5410] = 12'h222;
rom[5411] = 12'h222;
rom[5412] = 12'h222;
rom[5413] = 12'h222;
rom[5414] = 12'h333;
rom[5415] = 12'h333;
rom[5416] = 12'h222;
rom[5417] = 12'h  0;
rom[5418] = 12'h  0;
rom[5419] = 12'h  0;
rom[5420] = 12'h  0;
rom[5421] = 12'h  0;
rom[5422] = 12'h  0;
rom[5423] = 12'h  0;
rom[5424] = 12'h  0;
rom[5425] = 12'h  0;
rom[5426] = 12'h  0;
rom[5427] = 12'h  0;
rom[5428] = 12'h  0;
rom[5429] = 12'h  0;
rom[5430] = 12'h  0;
rom[5431] = 12'h  0;
rom[5432] = 12'h  0;
rom[5433] = 12'h  0;
rom[5434] = 12'h  0;
rom[5435] = 12'h  0;
rom[5436] = 12'h  0;
rom[5437] = 12'h  0;
rom[5438] = 12'h  0;
rom[5439] = 12'h  0;
rom[5440] = 12'h  0;
rom[5441] = 12'h  0;
rom[5442] = 12'h111;
rom[5443] = 12'h111;
rom[5444] = 12'h111;
rom[5445] = 12'h111;
rom[5446] = 12'h111;
rom[5447] = 12'h111;
rom[5448] = 12'h222;
rom[5449] = 12'h111;
rom[5450] = 12'h111;
rom[5451] = 12'h111;
rom[5452] = 12'h111;
rom[5453] = 12'h222;
rom[5454] = 12'h333;
rom[5455] = 12'h333;
rom[5456] = 12'h222;
rom[5457] = 12'h222;
rom[5458] = 12'h111;
rom[5459] = 12'h111;
rom[5460] = 12'h222;
rom[5461] = 12'h222;
rom[5462] = 12'h222;
rom[5463] = 12'h111;
rom[5464] = 12'h111;
rom[5465] = 12'h111;
rom[5466] = 12'h111;
rom[5467] = 12'h111;
rom[5468] = 12'h111;
rom[5469] = 12'h111;
rom[5470] = 12'h  0;
rom[5471] = 12'h  0;
rom[5472] = 12'h  0;
rom[5473] = 12'h  0;
rom[5474] = 12'h  0;
rom[5475] = 12'h  0;
rom[5476] = 12'h  0;
rom[5477] = 12'h  0;
rom[5478] = 12'h  0;
rom[5479] = 12'h  0;
rom[5480] = 12'h  0;
rom[5481] = 12'h  0;
rom[5482] = 12'h  0;
rom[5483] = 12'h  0;
rom[5484] = 12'h  0;
rom[5485] = 12'h  0;
rom[5486] = 12'h  0;
rom[5487] = 12'h  0;
rom[5488] = 12'h  0;
rom[5489] = 12'h  0;
rom[5490] = 12'h  0;
rom[5491] = 12'h  0;
rom[5492] = 12'h  0;
rom[5493] = 12'h  0;
rom[5494] = 12'h  0;
rom[5495] = 12'h  0;
rom[5496] = 12'h  0;
rom[5497] = 12'h  0;
rom[5498] = 12'h  0;
rom[5499] = 12'h  0;
rom[5500] = 12'h  0;
rom[5501] = 12'h111;
rom[5502] = 12'h111;
rom[5503] = 12'h  0;
rom[5504] = 12'h  0;
rom[5505] = 12'h  0;
rom[5506] = 12'h  0;
rom[5507] = 12'h  0;
rom[5508] = 12'h  0;
rom[5509] = 12'h  0;
rom[5510] = 12'h  0;
rom[5511] = 12'h  0;
rom[5512] = 12'h  0;
rom[5513] = 12'h  0;
rom[5514] = 12'h  0;
rom[5515] = 12'h  0;
rom[5516] = 12'h  0;
rom[5517] = 12'h  0;
rom[5518] = 12'h111;
rom[5519] = 12'h222;
rom[5520] = 12'h333;
rom[5521] = 12'h444;
rom[5522] = 12'h555;
rom[5523] = 12'h555;
rom[5524] = 12'h555;
rom[5525] = 12'h555;
rom[5526] = 12'h444;
rom[5527] = 12'h333;
rom[5528] = 12'h222;
rom[5529] = 12'h222;
rom[5530] = 12'h222;
rom[5531] = 12'h222;
rom[5532] = 12'h111;
rom[5533] = 12'h111;
rom[5534] = 12'h111;
rom[5535] = 12'h111;
rom[5536] = 12'h111;
rom[5537] = 12'h111;
rom[5538] = 12'h111;
rom[5539] = 12'h111;
rom[5540] = 12'h111;
rom[5541] = 12'h111;
rom[5542] = 12'h111;
rom[5543] = 12'h111;
rom[5544] = 12'h111;
rom[5545] = 12'h111;
rom[5546] = 12'h333;
rom[5547] = 12'h444;
rom[5548] = 12'h555;
rom[5549] = 12'h333;
rom[5550] = 12'h333;
rom[5551] = 12'h333;
rom[5552] = 12'h444;
rom[5553] = 12'h444;
rom[5554] = 12'h444;
rom[5555] = 12'h444;
rom[5556] = 12'h444;
rom[5557] = 12'h444;
rom[5558] = 12'h555;
rom[5559] = 12'h555;
rom[5560] = 12'h666;
rom[5561] = 12'h777;
rom[5562] = 12'h888;
rom[5563] = 12'h888;
rom[5564] = 12'h666;
rom[5565] = 12'h444;
rom[5566] = 12'h444;
rom[5567] = 12'h444;
rom[5568] = 12'h444;
rom[5569] = 12'h444;
rom[5570] = 12'h444;
rom[5571] = 12'h444;
rom[5572] = 12'h444;
rom[5573] = 12'h444;
rom[5574] = 12'h444;
rom[5575] = 12'h444;
rom[5576] = 12'h555;
rom[5577] = 12'h555;
rom[5578] = 12'h666;
rom[5579] = 12'h666;
rom[5580] = 12'h666;
rom[5581] = 12'h555;
rom[5582] = 12'h555;
rom[5583] = 12'h666;
rom[5584] = 12'h666;
rom[5585] = 12'h666;
rom[5586] = 12'h666;
rom[5587] = 12'h666;
rom[5588] = 12'h666;
rom[5589] = 12'h777;
rom[5590] = 12'h777;
rom[5591] = 12'h777;
rom[5592] = 12'h999;
rom[5593] = 12'h999;
rom[5594] = 12'h999;
rom[5595] = 12'haaa;
rom[5596] = 12'h999;
rom[5597] = 12'h999;
rom[5598] = 12'h999;
rom[5599] = 12'h999;
rom[5600] = 12'h444;
rom[5601] = 12'h444;
rom[5602] = 12'h444;
rom[5603] = 12'h444;
rom[5604] = 12'h444;
rom[5605] = 12'h555;
rom[5606] = 12'h555;
rom[5607] = 12'h555;
rom[5608] = 12'h555;
rom[5609] = 12'h555;
rom[5610] = 12'h555;
rom[5611] = 12'h444;
rom[5612] = 12'h444;
rom[5613] = 12'h444;
rom[5614] = 12'h333;
rom[5615] = 12'h333;
rom[5616] = 12'h222;
rom[5617] = 12'h222;
rom[5618] = 12'h222;
rom[5619] = 12'h222;
rom[5620] = 12'h222;
rom[5621] = 12'h111;
rom[5622] = 12'h111;
rom[5623] = 12'h111;
rom[5624] = 12'h111;
rom[5625] = 12'h111;
rom[5626] = 12'h111;
rom[5627] = 12'h111;
rom[5628] = 12'h111;
rom[5629] = 12'h111;
rom[5630] = 12'h111;
rom[5631] = 12'h111;
rom[5632] = 12'h111;
rom[5633] = 12'h111;
rom[5634] = 12'h111;
rom[5635] = 12'h111;
rom[5636] = 12'h111;
rom[5637] = 12'h111;
rom[5638] = 12'h111;
rom[5639] = 12'h111;
rom[5640] = 12'h  0;
rom[5641] = 12'h  0;
rom[5642] = 12'h  0;
rom[5643] = 12'h  0;
rom[5644] = 12'h  0;
rom[5645] = 12'h  0;
rom[5646] = 12'h  0;
rom[5647] = 12'h  0;
rom[5648] = 12'h  0;
rom[5649] = 12'h  0;
rom[5650] = 12'h  0;
rom[5651] = 12'h  0;
rom[5652] = 12'h  0;
rom[5653] = 12'h  0;
rom[5654] = 12'h  0;
rom[5655] = 12'h  0;
rom[5656] = 12'h  0;
rom[5657] = 12'h  0;
rom[5658] = 12'h  0;
rom[5659] = 12'h  0;
rom[5660] = 12'h  0;
rom[5661] = 12'h111;
rom[5662] = 12'h111;
rom[5663] = 12'h111;
rom[5664] = 12'h111;
rom[5665] = 12'h111;
rom[5666] = 12'h111;
rom[5667] = 12'h111;
rom[5668] = 12'h111;
rom[5669] = 12'h111;
rom[5670] = 12'h111;
rom[5671] = 12'h111;
rom[5672] = 12'h111;
rom[5673] = 12'h111;
rom[5674] = 12'h  0;
rom[5675] = 12'h  0;
rom[5676] = 12'h  0;
rom[5677] = 12'h  0;
rom[5678] = 12'h111;
rom[5679] = 12'h111;
rom[5680] = 12'h111;
rom[5681] = 12'h111;
rom[5682] = 12'h111;
rom[5683] = 12'h111;
rom[5684] = 12'h111;
rom[5685] = 12'h111;
rom[5686] = 12'h111;
rom[5687] = 12'h111;
rom[5688] = 12'h111;
rom[5689] = 12'h111;
rom[5690] = 12'h111;
rom[5691] = 12'h222;
rom[5692] = 12'h222;
rom[5693] = 12'h333;
rom[5694] = 12'h333;
rom[5695] = 12'h333;
rom[5696] = 12'h444;
rom[5697] = 12'h444;
rom[5698] = 12'h555;
rom[5699] = 12'h666;
rom[5700] = 12'h666;
rom[5701] = 12'h777;
rom[5702] = 12'h888;
rom[5703] = 12'h888;
rom[5704] = 12'h888;
rom[5705] = 12'h888;
rom[5706] = 12'h888;
rom[5707] = 12'h888;
rom[5708] = 12'h888;
rom[5709] = 12'h888;
rom[5710] = 12'h888;
rom[5711] = 12'h988;
rom[5712] = 12'h998;
rom[5713] = 12'ha97;
rom[5714] = 12'ha97;
rom[5715] = 12'ha97;
rom[5716] = 12'ha97;
rom[5717] = 12'ha97;
rom[5718] = 12'ha97;
rom[5719] = 12'ha97;
rom[5720] = 12'ha97;
rom[5721] = 12'ha97;
rom[5722] = 12'ha97;
rom[5723] = 12'ha87;
rom[5724] = 12'ha86;
rom[5725] = 12'h976;
rom[5726] = 12'h965;
rom[5727] = 12'h865;
rom[5728] = 12'h866;
rom[5729] = 12'h766;
rom[5730] = 12'h766;
rom[5731] = 12'h765;
rom[5732] = 12'h765;
rom[5733] = 12'h765;
rom[5734] = 12'h765;
rom[5735] = 12'h765;
rom[5736] = 12'h765;
rom[5737] = 12'h765;
rom[5738] = 12'h766;
rom[5739] = 12'h876;
rom[5740] = 12'h876;
rom[5741] = 12'h876;
rom[5742] = 12'h877;
rom[5743] = 12'h987;
rom[5744] = 12'h987;
rom[5745] = 12'h988;
rom[5746] = 12'ha88;
rom[5747] = 12'ha98;
rom[5748] = 12'ha98;
rom[5749] = 12'ha98;
rom[5750] = 12'ha98;
rom[5751] = 12'ha98;
rom[5752] = 12'ha99;
rom[5753] = 12'ha99;
rom[5754] = 12'haa9;
rom[5755] = 12'hba9;
rom[5756] = 12'hba9;
rom[5757] = 12'hba9;
rom[5758] = 12'hba9;
rom[5759] = 12'hbaa;
rom[5760] = 12'hbbb;
rom[5761] = 12'hbbb;
rom[5762] = 12'hbbb;
rom[5763] = 12'hbbb;
rom[5764] = 12'hbbb;
rom[5765] = 12'hbba;
rom[5766] = 12'haaa;
rom[5767] = 12'haaa;
rom[5768] = 12'haaa;
rom[5769] = 12'haaa;
rom[5770] = 12'haaa;
rom[5771] = 12'haaa;
rom[5772] = 12'h999;
rom[5773] = 12'h888;
rom[5774] = 12'h887;
rom[5775] = 12'h777;
rom[5776] = 12'h777;
rom[5777] = 12'h777;
rom[5778] = 12'h777;
rom[5779] = 12'h777;
rom[5780] = 12'h777;
rom[5781] = 12'h666;
rom[5782] = 12'h666;
rom[5783] = 12'h555;
rom[5784] = 12'h555;
rom[5785] = 12'h555;
rom[5786] = 12'h555;
rom[5787] = 12'h555;
rom[5788] = 12'h555;
rom[5789] = 12'h555;
rom[5790] = 12'h555;
rom[5791] = 12'h555;
rom[5792] = 12'h444;
rom[5793] = 12'h555;
rom[5794] = 12'h666;
rom[5795] = 12'h666;
rom[5796] = 12'h777;
rom[5797] = 12'h777;
rom[5798] = 12'h888;
rom[5799] = 12'h888;
rom[5800] = 12'h777;
rom[5801] = 12'h777;
rom[5802] = 12'h777;
rom[5803] = 12'h777;
rom[5804] = 12'h555;
rom[5805] = 12'h444;
rom[5806] = 12'h444;
rom[5807] = 12'h333;
rom[5808] = 12'h333;
rom[5809] = 12'h333;
rom[5810] = 12'h333;
rom[5811] = 12'h222;
rom[5812] = 12'h222;
rom[5813] = 12'h333;
rom[5814] = 12'h333;
rom[5815] = 12'h222;
rom[5816] = 12'h111;
rom[5817] = 12'h  0;
rom[5818] = 12'h  0;
rom[5819] = 12'h  0;
rom[5820] = 12'h  0;
rom[5821] = 12'h  0;
rom[5822] = 12'h  0;
rom[5823] = 12'h  0;
rom[5824] = 12'h  0;
rom[5825] = 12'h  0;
rom[5826] = 12'h  0;
rom[5827] = 12'h  0;
rom[5828] = 12'h  0;
rom[5829] = 12'h  0;
rom[5830] = 12'h  0;
rom[5831] = 12'h  0;
rom[5832] = 12'h  0;
rom[5833] = 12'h  0;
rom[5834] = 12'h  0;
rom[5835] = 12'h  0;
rom[5836] = 12'h  0;
rom[5837] = 12'h  0;
rom[5838] = 12'h  0;
rom[5839] = 12'h  0;
rom[5840] = 12'h  0;
rom[5841] = 12'h111;
rom[5842] = 12'h111;
rom[5843] = 12'h111;
rom[5844] = 12'h111;
rom[5845] = 12'h222;
rom[5846] = 12'h222;
rom[5847] = 12'h222;
rom[5848] = 12'h111;
rom[5849] = 12'h111;
rom[5850] = 12'h111;
rom[5851] = 12'h111;
rom[5852] = 12'h222;
rom[5853] = 12'h333;
rom[5854] = 12'h333;
rom[5855] = 12'h333;
rom[5856] = 12'h222;
rom[5857] = 12'h222;
rom[5858] = 12'h111;
rom[5859] = 12'h111;
rom[5860] = 12'h222;
rom[5861] = 12'h222;
rom[5862] = 12'h222;
rom[5863] = 12'h111;
rom[5864] = 12'h111;
rom[5865] = 12'h111;
rom[5866] = 12'h111;
rom[5867] = 12'h111;
rom[5868] = 12'h111;
rom[5869] = 12'h111;
rom[5870] = 12'h  0;
rom[5871] = 12'h  0;
rom[5872] = 12'h  0;
rom[5873] = 12'h  0;
rom[5874] = 12'h  0;
rom[5875] = 12'h  0;
rom[5876] = 12'h  0;
rom[5877] = 12'h  0;
rom[5878] = 12'h  0;
rom[5879] = 12'h  0;
rom[5880] = 12'h  0;
rom[5881] = 12'h  0;
rom[5882] = 12'h  0;
rom[5883] = 12'h  0;
rom[5884] = 12'h  0;
rom[5885] = 12'h  0;
rom[5886] = 12'h  0;
rom[5887] = 12'h  0;
rom[5888] = 12'h  0;
rom[5889] = 12'h  0;
rom[5890] = 12'h  0;
rom[5891] = 12'h  0;
rom[5892] = 12'h  0;
rom[5893] = 12'h  0;
rom[5894] = 12'h  0;
rom[5895] = 12'h  0;
rom[5896] = 12'h  0;
rom[5897] = 12'h  0;
rom[5898] = 12'h  0;
rom[5899] = 12'h  0;
rom[5900] = 12'h  0;
rom[5901] = 12'h111;
rom[5902] = 12'h111;
rom[5903] = 12'h  0;
rom[5904] = 12'h  0;
rom[5905] = 12'h  0;
rom[5906] = 12'h  0;
rom[5907] = 12'h  0;
rom[5908] = 12'h  0;
rom[5909] = 12'h  0;
rom[5910] = 12'h  0;
rom[5911] = 12'h  0;
rom[5912] = 12'h  0;
rom[5913] = 12'h  0;
rom[5914] = 12'h  0;
rom[5915] = 12'h  0;
rom[5916] = 12'h  0;
rom[5917] = 12'h  0;
rom[5918] = 12'h111;
rom[5919] = 12'h222;
rom[5920] = 12'h333;
rom[5921] = 12'h444;
rom[5922] = 12'h555;
rom[5923] = 12'h555;
rom[5924] = 12'h555;
rom[5925] = 12'h555;
rom[5926] = 12'h444;
rom[5927] = 12'h333;
rom[5928] = 12'h222;
rom[5929] = 12'h333;
rom[5930] = 12'h222;
rom[5931] = 12'h222;
rom[5932] = 12'h111;
rom[5933] = 12'h111;
rom[5934] = 12'h111;
rom[5935] = 12'h111;
rom[5936] = 12'h111;
rom[5937] = 12'h111;
rom[5938] = 12'h111;
rom[5939] = 12'h111;
rom[5940] = 12'h111;
rom[5941] = 12'h222;
rom[5942] = 12'h111;
rom[5943] = 12'h111;
rom[5944] = 12'h222;
rom[5945] = 12'h222;
rom[5946] = 12'h333;
rom[5947] = 12'h444;
rom[5948] = 12'h444;
rom[5949] = 12'h333;
rom[5950] = 12'h333;
rom[5951] = 12'h333;
rom[5952] = 12'h444;
rom[5953] = 12'h333;
rom[5954] = 12'h444;
rom[5955] = 12'h444;
rom[5956] = 12'h555;
rom[5957] = 12'h555;
rom[5958] = 12'h666;
rom[5959] = 12'h666;
rom[5960] = 12'h777;
rom[5961] = 12'h777;
rom[5962] = 12'h777;
rom[5963] = 12'h666;
rom[5964] = 12'h444;
rom[5965] = 12'h333;
rom[5966] = 12'h333;
rom[5967] = 12'h444;
rom[5968] = 12'h444;
rom[5969] = 12'h444;
rom[5970] = 12'h444;
rom[5971] = 12'h444;
rom[5972] = 12'h444;
rom[5973] = 12'h444;
rom[5974] = 12'h444;
rom[5975] = 12'h444;
rom[5976] = 12'h555;
rom[5977] = 12'h555;
rom[5978] = 12'h555;
rom[5979] = 12'h555;
rom[5980] = 12'h555;
rom[5981] = 12'h555;
rom[5982] = 12'h555;
rom[5983] = 12'h555;
rom[5984] = 12'h666;
rom[5985] = 12'h666;
rom[5986] = 12'h666;
rom[5987] = 12'h666;
rom[5988] = 12'h666;
rom[5989] = 12'h777;
rom[5990] = 12'h777;
rom[5991] = 12'h777;
rom[5992] = 12'h888;
rom[5993] = 12'h999;
rom[5994] = 12'h999;
rom[5995] = 12'haaa;
rom[5996] = 12'haaa;
rom[5997] = 12'h999;
rom[5998] = 12'h999;
rom[5999] = 12'h999;
rom[6000] = 12'h444;
rom[6001] = 12'h444;
rom[6002] = 12'h555;
rom[6003] = 12'h555;
rom[6004] = 12'h555;
rom[6005] = 12'h666;
rom[6006] = 12'h666;
rom[6007] = 12'h666;
rom[6008] = 12'h555;
rom[6009] = 12'h555;
rom[6010] = 12'h444;
rom[6011] = 12'h444;
rom[6012] = 12'h444;
rom[6013] = 12'h333;
rom[6014] = 12'h333;
rom[6015] = 12'h222;
rom[6016] = 12'h222;
rom[6017] = 12'h222;
rom[6018] = 12'h222;
rom[6019] = 12'h222;
rom[6020] = 12'h222;
rom[6021] = 12'h111;
rom[6022] = 12'h111;
rom[6023] = 12'h111;
rom[6024] = 12'h111;
rom[6025] = 12'h111;
rom[6026] = 12'h111;
rom[6027] = 12'h111;
rom[6028] = 12'h111;
rom[6029] = 12'h111;
rom[6030] = 12'h111;
rom[6031] = 12'h111;
rom[6032] = 12'h111;
rom[6033] = 12'h111;
rom[6034] = 12'h111;
rom[6035] = 12'h111;
rom[6036] = 12'h111;
rom[6037] = 12'h111;
rom[6038] = 12'h111;
rom[6039] = 12'h111;
rom[6040] = 12'h  0;
rom[6041] = 12'h  0;
rom[6042] = 12'h  0;
rom[6043] = 12'h  0;
rom[6044] = 12'h  0;
rom[6045] = 12'h  0;
rom[6046] = 12'h  0;
rom[6047] = 12'h  0;
rom[6048] = 12'h  0;
rom[6049] = 12'h  0;
rom[6050] = 12'h  0;
rom[6051] = 12'h  0;
rom[6052] = 12'h  0;
rom[6053] = 12'h  0;
rom[6054] = 12'h  0;
rom[6055] = 12'h  0;
rom[6056] = 12'h  0;
rom[6057] = 12'h  0;
rom[6058] = 12'h  0;
rom[6059] = 12'h  0;
rom[6060] = 12'h  0;
rom[6061] = 12'h  0;
rom[6062] = 12'h111;
rom[6063] = 12'h111;
rom[6064] = 12'h111;
rom[6065] = 12'h111;
rom[6066] = 12'h111;
rom[6067] = 12'h111;
rom[6068] = 12'h111;
rom[6069] = 12'h111;
rom[6070] = 12'h111;
rom[6071] = 12'h111;
rom[6072] = 12'h111;
rom[6073] = 12'h111;
rom[6074] = 12'h  0;
rom[6075] = 12'h  0;
rom[6076] = 12'h  0;
rom[6077] = 12'h  0;
rom[6078] = 12'h  0;
rom[6079] = 12'h111;
rom[6080] = 12'h  0;
rom[6081] = 12'h  0;
rom[6082] = 12'h  0;
rom[6083] = 12'h  0;
rom[6084] = 12'h  0;
rom[6085] = 12'h111;
rom[6086] = 12'h111;
rom[6087] = 12'h111;
rom[6088] = 12'h111;
rom[6089] = 12'h222;
rom[6090] = 12'h222;
rom[6091] = 12'h222;
rom[6092] = 12'h333;
rom[6093] = 12'h333;
rom[6094] = 12'h333;
rom[6095] = 12'h333;
rom[6096] = 12'h444;
rom[6097] = 12'h444;
rom[6098] = 12'h555;
rom[6099] = 12'h555;
rom[6100] = 12'h666;
rom[6101] = 12'h777;
rom[6102] = 12'h777;
rom[6103] = 12'h777;
rom[6104] = 12'h666;
rom[6105] = 12'h666;
rom[6106] = 12'h666;
rom[6107] = 12'h666;
rom[6108] = 12'h666;
rom[6109] = 12'h766;
rom[6110] = 12'h777;
rom[6111] = 12'h877;
rom[6112] = 12'h876;
rom[6113] = 12'h876;
rom[6114] = 12'h875;
rom[6115] = 12'h875;
rom[6116] = 12'h986;
rom[6117] = 12'h986;
rom[6118] = 12'ha86;
rom[6119] = 12'ha86;
rom[6120] = 12'ha85;
rom[6121] = 12'ha86;
rom[6122] = 12'ha86;
rom[6123] = 12'ha86;
rom[6124] = 12'ha75;
rom[6125] = 12'h975;
rom[6126] = 12'h965;
rom[6127] = 12'h864;
rom[6128] = 12'h754;
rom[6129] = 12'h654;
rom[6130] = 12'h653;
rom[6131] = 12'h643;
rom[6132] = 12'h643;
rom[6133] = 12'h543;
rom[6134] = 12'h543;
rom[6135] = 12'h542;
rom[6136] = 12'h643;
rom[6137] = 12'h643;
rom[6138] = 12'h643;
rom[6139] = 12'h643;
rom[6140] = 12'h643;
rom[6141] = 12'h654;
rom[6142] = 12'h754;
rom[6143] = 12'h754;
rom[6144] = 12'h765;
rom[6145] = 12'h865;
rom[6146] = 12'h865;
rom[6147] = 12'h976;
rom[6148] = 12'h976;
rom[6149] = 12'h976;
rom[6150] = 12'h987;
rom[6151] = 12'ha87;
rom[6152] = 12'ha87;
rom[6153] = 12'ha87;
rom[6154] = 12'ha87;
rom[6155] = 12'ha98;
rom[6156] = 12'ha98;
rom[6157] = 12'hb98;
rom[6158] = 12'hba9;
rom[6159] = 12'hba9;
rom[6160] = 12'haa9;
rom[6161] = 12'haa9;
rom[6162] = 12'haaa;
rom[6163] = 12'haaa;
rom[6164] = 12'hbba;
rom[6165] = 12'hbba;
rom[6166] = 12'hbba;
rom[6167] = 12'hbba;
rom[6168] = 12'hbbb;
rom[6169] = 12'hbbb;
rom[6170] = 12'hbbb;
rom[6171] = 12'hbbb;
rom[6172] = 12'hbbb;
rom[6173] = 12'haaa;
rom[6174] = 12'h999;
rom[6175] = 12'h999;
rom[6176] = 12'h888;
rom[6177] = 12'h778;
rom[6178] = 12'h777;
rom[6179] = 12'h777;
rom[6180] = 12'h777;
rom[6181] = 12'h777;
rom[6182] = 12'h666;
rom[6183] = 12'h666;
rom[6184] = 12'h555;
rom[6185] = 12'h555;
rom[6186] = 12'h555;
rom[6187] = 12'h555;
rom[6188] = 12'h555;
rom[6189] = 12'h555;
rom[6190] = 12'h555;
rom[6191] = 12'h555;
rom[6192] = 12'h444;
rom[6193] = 12'h555;
rom[6194] = 12'h666;
rom[6195] = 12'h666;
rom[6196] = 12'h666;
rom[6197] = 12'h888;
rom[6198] = 12'h888;
rom[6199] = 12'h888;
rom[6200] = 12'h888;
rom[6201] = 12'h777;
rom[6202] = 12'h888;
rom[6203] = 12'h777;
rom[6204] = 12'h555;
rom[6205] = 12'h444;
rom[6206] = 12'h444;
rom[6207] = 12'h444;
rom[6208] = 12'h333;
rom[6209] = 12'h333;
rom[6210] = 12'h333;
rom[6211] = 12'h222;
rom[6212] = 12'h222;
rom[6213] = 12'h333;
rom[6214] = 12'h333;
rom[6215] = 12'h222;
rom[6216] = 12'h111;
rom[6217] = 12'h  0;
rom[6218] = 12'h  0;
rom[6219] = 12'h  0;
rom[6220] = 12'h  0;
rom[6221] = 12'h  0;
rom[6222] = 12'h  0;
rom[6223] = 12'h  0;
rom[6224] = 12'h  0;
rom[6225] = 12'h  0;
rom[6226] = 12'h  0;
rom[6227] = 12'h  0;
rom[6228] = 12'h  0;
rom[6229] = 12'h  0;
rom[6230] = 12'h  0;
rom[6231] = 12'h  0;
rom[6232] = 12'h  0;
rom[6233] = 12'h  0;
rom[6234] = 12'h  0;
rom[6235] = 12'h  0;
rom[6236] = 12'h  0;
rom[6237] = 12'h  0;
rom[6238] = 12'h  0;
rom[6239] = 12'h  0;
rom[6240] = 12'h111;
rom[6241] = 12'h111;
rom[6242] = 12'h111;
rom[6243] = 12'h222;
rom[6244] = 12'h222;
rom[6245] = 12'h222;
rom[6246] = 12'h222;
rom[6247] = 12'h222;
rom[6248] = 12'h111;
rom[6249] = 12'h111;
rom[6250] = 12'h111;
rom[6251] = 12'h222;
rom[6252] = 12'h222;
rom[6253] = 12'h333;
rom[6254] = 12'h333;
rom[6255] = 12'h333;
rom[6256] = 12'h222;
rom[6257] = 12'h222;
rom[6258] = 12'h111;
rom[6259] = 12'h222;
rom[6260] = 12'h222;
rom[6261] = 12'h222;
rom[6262] = 12'h222;
rom[6263] = 12'h222;
rom[6264] = 12'h111;
rom[6265] = 12'h222;
rom[6266] = 12'h111;
rom[6267] = 12'h111;
rom[6268] = 12'h  0;
rom[6269] = 12'h  0;
rom[6270] = 12'h  0;
rom[6271] = 12'h  0;
rom[6272] = 12'h  0;
rom[6273] = 12'h  0;
rom[6274] = 12'h  0;
rom[6275] = 12'h  0;
rom[6276] = 12'h  0;
rom[6277] = 12'h  0;
rom[6278] = 12'h  0;
rom[6279] = 12'h  0;
rom[6280] = 12'h  0;
rom[6281] = 12'h  0;
rom[6282] = 12'h  0;
rom[6283] = 12'h  0;
rom[6284] = 12'h  0;
rom[6285] = 12'h  0;
rom[6286] = 12'h  0;
rom[6287] = 12'h  0;
rom[6288] = 12'h  0;
rom[6289] = 12'h  0;
rom[6290] = 12'h  0;
rom[6291] = 12'h  0;
rom[6292] = 12'h  0;
rom[6293] = 12'h  0;
rom[6294] = 12'h  0;
rom[6295] = 12'h  0;
rom[6296] = 12'h  0;
rom[6297] = 12'h  0;
rom[6298] = 12'h  0;
rom[6299] = 12'h  0;
rom[6300] = 12'h  0;
rom[6301] = 12'h111;
rom[6302] = 12'h111;
rom[6303] = 12'h  0;
rom[6304] = 12'h  0;
rom[6305] = 12'h  0;
rom[6306] = 12'h  0;
rom[6307] = 12'h  0;
rom[6308] = 12'h  0;
rom[6309] = 12'h  0;
rom[6310] = 12'h  0;
rom[6311] = 12'h  0;
rom[6312] = 12'h  0;
rom[6313] = 12'h  0;
rom[6314] = 12'h  0;
rom[6315] = 12'h  0;
rom[6316] = 12'h  0;
rom[6317] = 12'h  0;
rom[6318] = 12'h111;
rom[6319] = 12'h222;
rom[6320] = 12'h333;
rom[6321] = 12'h444;
rom[6322] = 12'h555;
rom[6323] = 12'h666;
rom[6324] = 12'h666;
rom[6325] = 12'h555;
rom[6326] = 12'h444;
rom[6327] = 12'h333;
rom[6328] = 12'h222;
rom[6329] = 12'h333;
rom[6330] = 12'h222;
rom[6331] = 12'h111;
rom[6332] = 12'h111;
rom[6333] = 12'h111;
rom[6334] = 12'h222;
rom[6335] = 12'h111;
rom[6336] = 12'h111;
rom[6337] = 12'h111;
rom[6338] = 12'h111;
rom[6339] = 12'h111;
rom[6340] = 12'h222;
rom[6341] = 12'h222;
rom[6342] = 12'h111;
rom[6343] = 12'h111;
rom[6344] = 12'h222;
rom[6345] = 12'h333;
rom[6346] = 12'h333;
rom[6347] = 12'h333;
rom[6348] = 12'h333;
rom[6349] = 12'h333;
rom[6350] = 12'h333;
rom[6351] = 12'h333;
rom[6352] = 12'h444;
rom[6353] = 12'h444;
rom[6354] = 12'h444;
rom[6355] = 12'h444;
rom[6356] = 12'h555;
rom[6357] = 12'h666;
rom[6358] = 12'h666;
rom[6359] = 12'h777;
rom[6360] = 12'h666;
rom[6361] = 12'h666;
rom[6362] = 12'h555;
rom[6363] = 12'h444;
rom[6364] = 12'h444;
rom[6365] = 12'h333;
rom[6366] = 12'h444;
rom[6367] = 12'h444;
rom[6368] = 12'h444;
rom[6369] = 12'h444;
rom[6370] = 12'h333;
rom[6371] = 12'h444;
rom[6372] = 12'h444;
rom[6373] = 12'h555;
rom[6374] = 12'h555;
rom[6375] = 12'h555;
rom[6376] = 12'h444;
rom[6377] = 12'h555;
rom[6378] = 12'h555;
rom[6379] = 12'h555;
rom[6380] = 12'h444;
rom[6381] = 12'h444;
rom[6382] = 12'h555;
rom[6383] = 12'h555;
rom[6384] = 12'h666;
rom[6385] = 12'h666;
rom[6386] = 12'h666;
rom[6387] = 12'h777;
rom[6388] = 12'h777;
rom[6389] = 12'h777;
rom[6390] = 12'h777;
rom[6391] = 12'h777;
rom[6392] = 12'h888;
rom[6393] = 12'h999;
rom[6394] = 12'h999;
rom[6395] = 12'haaa;
rom[6396] = 12'haaa;
rom[6397] = 12'h999;
rom[6398] = 12'h999;
rom[6399] = 12'h999;
rom[6400] = 12'h666;
rom[6401] = 12'h666;
rom[6402] = 12'h666;
rom[6403] = 12'h666;
rom[6404] = 12'h666;
rom[6405] = 12'h666;
rom[6406] = 12'h555;
rom[6407] = 12'h555;
rom[6408] = 12'h444;
rom[6409] = 12'h444;
rom[6410] = 12'h333;
rom[6411] = 12'h333;
rom[6412] = 12'h333;
rom[6413] = 12'h333;
rom[6414] = 12'h222;
rom[6415] = 12'h222;
rom[6416] = 12'h222;
rom[6417] = 12'h222;
rom[6418] = 12'h222;
rom[6419] = 12'h222;
rom[6420] = 12'h111;
rom[6421] = 12'h111;
rom[6422] = 12'h111;
rom[6423] = 12'h111;
rom[6424] = 12'h111;
rom[6425] = 12'h111;
rom[6426] = 12'h111;
rom[6427] = 12'h  0;
rom[6428] = 12'h  0;
rom[6429] = 12'h111;
rom[6430] = 12'h111;
rom[6431] = 12'h111;
rom[6432] = 12'h111;
rom[6433] = 12'h111;
rom[6434] = 12'h111;
rom[6435] = 12'h111;
rom[6436] = 12'h111;
rom[6437] = 12'h111;
rom[6438] = 12'h111;
rom[6439] = 12'h111;
rom[6440] = 12'h  0;
rom[6441] = 12'h  0;
rom[6442] = 12'h  0;
rom[6443] = 12'h  0;
rom[6444] = 12'h  0;
rom[6445] = 12'h  0;
rom[6446] = 12'h  0;
rom[6447] = 12'h  0;
rom[6448] = 12'h  0;
rom[6449] = 12'h  0;
rom[6450] = 12'h  0;
rom[6451] = 12'h  0;
rom[6452] = 12'h  0;
rom[6453] = 12'h  0;
rom[6454] = 12'h  0;
rom[6455] = 12'h  0;
rom[6456] = 12'h  0;
rom[6457] = 12'h  0;
rom[6458] = 12'h  0;
rom[6459] = 12'h  0;
rom[6460] = 12'h  0;
rom[6461] = 12'h  0;
rom[6462] = 12'h111;
rom[6463] = 12'h111;
rom[6464] = 12'h111;
rom[6465] = 12'h111;
rom[6466] = 12'h111;
rom[6467] = 12'h111;
rom[6468] = 12'h111;
rom[6469] = 12'h111;
rom[6470] = 12'h111;
rom[6471] = 12'h111;
rom[6472] = 12'h  0;
rom[6473] = 12'h  0;
rom[6474] = 12'h  0;
rom[6475] = 12'h  0;
rom[6476] = 12'h  0;
rom[6477] = 12'h111;
rom[6478] = 12'h111;
rom[6479] = 12'h111;
rom[6480] = 12'h111;
rom[6481] = 12'h  0;
rom[6482] = 12'h  0;
rom[6483] = 12'h  0;
rom[6484] = 12'h  0;
rom[6485] = 12'h111;
rom[6486] = 12'h111;
rom[6487] = 12'h111;
rom[6488] = 12'h222;
rom[6489] = 12'h111;
rom[6490] = 12'h111;
rom[6491] = 12'h111;
rom[6492] = 12'h111;
rom[6493] = 12'h222;
rom[6494] = 12'h333;
rom[6495] = 12'h333;
rom[6496] = 12'h333;
rom[6497] = 12'h444;
rom[6498] = 12'h555;
rom[6499] = 12'h666;
rom[6500] = 12'h666;
rom[6501] = 12'h565;
rom[6502] = 12'h555;
rom[6503] = 12'h444;
rom[6504] = 12'h444;
rom[6505] = 12'h444;
rom[6506] = 12'h555;
rom[6507] = 12'h666;
rom[6508] = 12'h666;
rom[6509] = 12'h666;
rom[6510] = 12'h766;
rom[6511] = 12'h877;
rom[6512] = 12'h876;
rom[6513] = 12'h865;
rom[6514] = 12'h864;
rom[6515] = 12'h864;
rom[6516] = 12'h975;
rom[6517] = 12'h975;
rom[6518] = 12'ha85;
rom[6519] = 12'ha85;
rom[6520] = 12'hb85;
rom[6521] = 12'hb95;
rom[6522] = 12'hb85;
rom[6523] = 12'hb85;
rom[6524] = 12'ha75;
rom[6525] = 12'ha74;
rom[6526] = 12'h964;
rom[6527] = 12'h853;
rom[6528] = 12'h753;
rom[6529] = 12'h643;
rom[6530] = 12'h642;
rom[6531] = 12'h531;
rom[6532] = 12'h521;
rom[6533] = 12'h521;
rom[6534] = 12'h521;
rom[6535] = 12'h521;
rom[6536] = 12'h521;
rom[6537] = 12'h521;
rom[6538] = 12'h521;
rom[6539] = 12'h531;
rom[6540] = 12'h531;
rom[6541] = 12'h631;
rom[6542] = 12'h632;
rom[6543] = 12'h631;
rom[6544] = 12'h642;
rom[6545] = 12'h742;
rom[6546] = 12'h742;
rom[6547] = 12'h742;
rom[6548] = 12'h743;
rom[6549] = 12'h853;
rom[6550] = 12'h854;
rom[6551] = 12'h854;
rom[6552] = 12'h864;
rom[6553] = 12'h864;
rom[6554] = 12'h864;
rom[6555] = 12'h864;
rom[6556] = 12'h865;
rom[6557] = 12'h975;
rom[6558] = 12'h976;
rom[6559] = 12'h976;
rom[6560] = 12'h986;
rom[6561] = 12'h987;
rom[6562] = 12'h987;
rom[6563] = 12'ha98;
rom[6564] = 12'ha98;
rom[6565] = 12'ha99;
rom[6566] = 12'haa9;
rom[6567] = 12'haa9;
rom[6568] = 12'hbaa;
rom[6569] = 12'haaa;
rom[6570] = 12'haaa;
rom[6571] = 12'haaa;
rom[6572] = 12'hbbb;
rom[6573] = 12'hbbb;
rom[6574] = 12'hbbb;
rom[6575] = 12'habb;
rom[6576] = 12'haaa;
rom[6577] = 12'h99a;
rom[6578] = 12'h999;
rom[6579] = 12'h899;
rom[6580] = 12'h899;
rom[6581] = 12'h888;
rom[6582] = 12'h778;
rom[6583] = 12'h777;
rom[6584] = 12'h666;
rom[6585] = 12'h666;
rom[6586] = 12'h655;
rom[6587] = 12'h655;
rom[6588] = 12'h555;
rom[6589] = 12'h555;
rom[6590] = 12'h555;
rom[6591] = 12'h555;
rom[6592] = 12'h555;
rom[6593] = 12'h555;
rom[6594] = 12'h555;
rom[6595] = 12'h666;
rom[6596] = 12'h666;
rom[6597] = 12'h777;
rom[6598] = 12'h888;
rom[6599] = 12'h999;
rom[6600] = 12'h888;
rom[6601] = 12'h888;
rom[6602] = 12'h888;
rom[6603] = 12'h777;
rom[6604] = 12'h666;
rom[6605] = 12'h444;
rom[6606] = 12'h444;
rom[6607] = 12'h444;
rom[6608] = 12'h444;
rom[6609] = 12'h222;
rom[6610] = 12'h222;
rom[6611] = 12'h333;
rom[6612] = 12'h333;
rom[6613] = 12'h333;
rom[6614] = 12'h222;
rom[6615] = 12'h222;
rom[6616] = 12'h111;
rom[6617] = 12'h  0;
rom[6618] = 12'h  0;
rom[6619] = 12'h  0;
rom[6620] = 12'h  0;
rom[6621] = 12'h  0;
rom[6622] = 12'h  0;
rom[6623] = 12'h  0;
rom[6624] = 12'h  0;
rom[6625] = 12'h  0;
rom[6626] = 12'h  0;
rom[6627] = 12'h  0;
rom[6628] = 12'h  0;
rom[6629] = 12'h  0;
rom[6630] = 12'h  0;
rom[6631] = 12'h  0;
rom[6632] = 12'h  0;
rom[6633] = 12'h  0;
rom[6634] = 12'h  0;
rom[6635] = 12'h  0;
rom[6636] = 12'h  0;
rom[6637] = 12'h  0;
rom[6638] = 12'h  0;
rom[6639] = 12'h  0;
rom[6640] = 12'h111;
rom[6641] = 12'h111;
rom[6642] = 12'h111;
rom[6643] = 12'h222;
rom[6644] = 12'h222;
rom[6645] = 12'h222;
rom[6646] = 12'h222;
rom[6647] = 12'h111;
rom[6648] = 12'h111;
rom[6649] = 12'h111;
rom[6650] = 12'h222;
rom[6651] = 12'h333;
rom[6652] = 12'h333;
rom[6653] = 12'h333;
rom[6654] = 12'h222;
rom[6655] = 12'h222;
rom[6656] = 12'h222;
rom[6657] = 12'h222;
rom[6658] = 12'h111;
rom[6659] = 12'h111;
rom[6660] = 12'h222;
rom[6661] = 12'h222;
rom[6662] = 12'h222;
rom[6663] = 12'h222;
rom[6664] = 12'h111;
rom[6665] = 12'h111;
rom[6666] = 12'h111;
rom[6667] = 12'h111;
rom[6668] = 12'h111;
rom[6669] = 12'h  0;
rom[6670] = 12'h  0;
rom[6671] = 12'h  0;
rom[6672] = 12'h  0;
rom[6673] = 12'h  0;
rom[6674] = 12'h  0;
rom[6675] = 12'h  0;
rom[6676] = 12'h  0;
rom[6677] = 12'h  0;
rom[6678] = 12'h  0;
rom[6679] = 12'h  0;
rom[6680] = 12'h  0;
rom[6681] = 12'h  0;
rom[6682] = 12'h  0;
rom[6683] = 12'h  0;
rom[6684] = 12'h  0;
rom[6685] = 12'h  0;
rom[6686] = 12'h  0;
rom[6687] = 12'h  0;
rom[6688] = 12'h  0;
rom[6689] = 12'h  0;
rom[6690] = 12'h  0;
rom[6691] = 12'h  0;
rom[6692] = 12'h  0;
rom[6693] = 12'h  0;
rom[6694] = 12'h  0;
rom[6695] = 12'h  0;
rom[6696] = 12'h  0;
rom[6697] = 12'h  0;
rom[6698] = 12'h  0;
rom[6699] = 12'h  0;
rom[6700] = 12'h111;
rom[6701] = 12'h111;
rom[6702] = 12'h111;
rom[6703] = 12'h  0;
rom[6704] = 12'h  0;
rom[6705] = 12'h  0;
rom[6706] = 12'h  0;
rom[6707] = 12'h  0;
rom[6708] = 12'h  0;
rom[6709] = 12'h  0;
rom[6710] = 12'h  0;
rom[6711] = 12'h  0;
rom[6712] = 12'h  0;
rom[6713] = 12'h  0;
rom[6714] = 12'h  0;
rom[6715] = 12'h  0;
rom[6716] = 12'h  0;
rom[6717] = 12'h111;
rom[6718] = 12'h111;
rom[6719] = 12'h222;
rom[6720] = 12'h444;
rom[6721] = 12'h555;
rom[6722] = 12'h666;
rom[6723] = 12'h666;
rom[6724] = 12'h555;
rom[6725] = 12'h555;
rom[6726] = 12'h444;
rom[6727] = 12'h333;
rom[6728] = 12'h333;
rom[6729] = 12'h333;
rom[6730] = 12'h222;
rom[6731] = 12'h222;
rom[6732] = 12'h222;
rom[6733] = 12'h111;
rom[6734] = 12'h111;
rom[6735] = 12'h111;
rom[6736] = 12'h111;
rom[6737] = 12'h111;
rom[6738] = 12'h111;
rom[6739] = 12'h111;
rom[6740] = 12'h111;
rom[6741] = 12'h111;
rom[6742] = 12'h111;
rom[6743] = 12'h111;
rom[6744] = 12'h333;
rom[6745] = 12'h333;
rom[6746] = 12'h333;
rom[6747] = 12'h222;
rom[6748] = 12'h222;
rom[6749] = 12'h333;
rom[6750] = 12'h333;
rom[6751] = 12'h333;
rom[6752] = 12'h444;
rom[6753] = 12'h444;
rom[6754] = 12'h444;
rom[6755] = 12'h555;
rom[6756] = 12'h555;
rom[6757] = 12'h666;
rom[6758] = 12'h666;
rom[6759] = 12'h666;
rom[6760] = 12'h555;
rom[6761] = 12'h555;
rom[6762] = 12'h444;
rom[6763] = 12'h444;
rom[6764] = 12'h444;
rom[6765] = 12'h444;
rom[6766] = 12'h444;
rom[6767] = 12'h444;
rom[6768] = 12'h444;
rom[6769] = 12'h444;
rom[6770] = 12'h444;
rom[6771] = 12'h555;
rom[6772] = 12'h555;
rom[6773] = 12'h555;
rom[6774] = 12'h555;
rom[6775] = 12'h555;
rom[6776] = 12'h444;
rom[6777] = 12'h444;
rom[6778] = 12'h444;
rom[6779] = 12'h444;
rom[6780] = 12'h444;
rom[6781] = 12'h444;
rom[6782] = 12'h555;
rom[6783] = 12'h555;
rom[6784] = 12'h555;
rom[6785] = 12'h555;
rom[6786] = 12'h666;
rom[6787] = 12'h666;
rom[6788] = 12'h777;
rom[6789] = 12'h777;
rom[6790] = 12'h777;
rom[6791] = 12'h777;
rom[6792] = 12'h888;
rom[6793] = 12'h999;
rom[6794] = 12'h999;
rom[6795] = 12'haaa;
rom[6796] = 12'haaa;
rom[6797] = 12'h999;
rom[6798] = 12'h999;
rom[6799] = 12'h999;
rom[6800] = 12'h666;
rom[6801] = 12'h666;
rom[6802] = 12'h666;
rom[6803] = 12'h666;
rom[6804] = 12'h555;
rom[6805] = 12'h555;
rom[6806] = 12'h555;
rom[6807] = 12'h444;
rom[6808] = 12'h444;
rom[6809] = 12'h333;
rom[6810] = 12'h333;
rom[6811] = 12'h333;
rom[6812] = 12'h222;
rom[6813] = 12'h222;
rom[6814] = 12'h222;
rom[6815] = 12'h222;
rom[6816] = 12'h222;
rom[6817] = 12'h222;
rom[6818] = 12'h222;
rom[6819] = 12'h111;
rom[6820] = 12'h111;
rom[6821] = 12'h111;
rom[6822] = 12'h111;
rom[6823] = 12'h111;
rom[6824] = 12'h111;
rom[6825] = 12'h111;
rom[6826] = 12'h111;
rom[6827] = 12'h  0;
rom[6828] = 12'h  0;
rom[6829] = 12'h111;
rom[6830] = 12'h111;
rom[6831] = 12'h111;
rom[6832] = 12'h111;
rom[6833] = 12'h111;
rom[6834] = 12'h111;
rom[6835] = 12'h111;
rom[6836] = 12'h111;
rom[6837] = 12'h111;
rom[6838] = 12'h111;
rom[6839] = 12'h111;
rom[6840] = 12'h  0;
rom[6841] = 12'h  0;
rom[6842] = 12'h  0;
rom[6843] = 12'h  0;
rom[6844] = 12'h  0;
rom[6845] = 12'h  0;
rom[6846] = 12'h  0;
rom[6847] = 12'h  0;
rom[6848] = 12'h  0;
rom[6849] = 12'h  0;
rom[6850] = 12'h  0;
rom[6851] = 12'h  0;
rom[6852] = 12'h  0;
rom[6853] = 12'h  0;
rom[6854] = 12'h  0;
rom[6855] = 12'h  0;
rom[6856] = 12'h  0;
rom[6857] = 12'h  0;
rom[6858] = 12'h  0;
rom[6859] = 12'h  0;
rom[6860] = 12'h111;
rom[6861] = 12'h111;
rom[6862] = 12'h111;
rom[6863] = 12'h111;
rom[6864] = 12'h111;
rom[6865] = 12'h111;
rom[6866] = 12'h111;
rom[6867] = 12'h111;
rom[6868] = 12'h111;
rom[6869] = 12'h111;
rom[6870] = 12'h111;
rom[6871] = 12'h111;
rom[6872] = 12'h  0;
rom[6873] = 12'h  0;
rom[6874] = 12'h  0;
rom[6875] = 12'h  0;
rom[6876] = 12'h111;
rom[6877] = 12'h111;
rom[6878] = 12'h111;
rom[6879] = 12'h111;
rom[6880] = 12'h111;
rom[6881] = 12'h111;
rom[6882] = 12'h  0;
rom[6883] = 12'h  0;
rom[6884] = 12'h  0;
rom[6885] = 12'h111;
rom[6886] = 12'h111;
rom[6887] = 12'h111;
rom[6888] = 12'h111;
rom[6889] = 12'h111;
rom[6890] = 12'h111;
rom[6891] = 12'h111;
rom[6892] = 12'h111;
rom[6893] = 12'h222;
rom[6894] = 12'h333;
rom[6895] = 12'h333;
rom[6896] = 12'h444;
rom[6897] = 12'h444;
rom[6898] = 12'h444;
rom[6899] = 12'h444;
rom[6900] = 12'h444;
rom[6901] = 12'h444;
rom[6902] = 12'h344;
rom[6903] = 12'h343;
rom[6904] = 12'h444;
rom[6905] = 12'h444;
rom[6906] = 12'h555;
rom[6907] = 12'h666;
rom[6908] = 12'h656;
rom[6909] = 12'h655;
rom[6910] = 12'h655;
rom[6911] = 12'h765;
rom[6912] = 12'h754;
rom[6913] = 12'h754;
rom[6914] = 12'h753;
rom[6915] = 12'h753;
rom[6916] = 12'h863;
rom[6917] = 12'h974;
rom[6918] = 12'ha74;
rom[6919] = 12'ha74;
rom[6920] = 12'hb84;
rom[6921] = 12'hb84;
rom[6922] = 12'hb84;
rom[6923] = 12'hb74;
rom[6924] = 12'ha73;
rom[6925] = 12'h963;
rom[6926] = 12'h952;
rom[6927] = 12'h842;
rom[6928] = 12'h742;
rom[6929] = 12'h631;
rom[6930] = 12'h531;
rom[6931] = 12'h520;
rom[6932] = 12'h520;
rom[6933] = 12'h520;
rom[6934] = 12'h520;
rom[6935] = 12'h520;
rom[6936] = 12'h521;
rom[6937] = 12'h520;
rom[6938] = 12'h621;
rom[6939] = 12'h620;
rom[6940] = 12'h621;
rom[6941] = 12'h621;
rom[6942] = 12'h631;
rom[6943] = 12'h631;
rom[6944] = 12'h631;
rom[6945] = 12'h631;
rom[6946] = 12'h631;
rom[6947] = 12'h631;
rom[6948] = 12'h631;
rom[6949] = 12'h731;
rom[6950] = 12'h731;
rom[6951] = 12'h731;
rom[6952] = 12'h742;
rom[6953] = 12'h642;
rom[6954] = 12'h642;
rom[6955] = 12'h642;
rom[6956] = 12'h642;
rom[6957] = 12'h642;
rom[6958] = 12'h743;
rom[6959] = 12'h753;
rom[6960] = 12'h764;
rom[6961] = 12'h865;
rom[6962] = 12'h875;
rom[6963] = 12'h876;
rom[6964] = 12'h986;
rom[6965] = 12'h987;
rom[6966] = 12'h987;
rom[6967] = 12'h988;
rom[6968] = 12'h998;
rom[6969] = 12'h999;
rom[6970] = 12'h999;
rom[6971] = 12'h999;
rom[6972] = 12'h999;
rom[6973] = 12'ha9a;
rom[6974] = 12'haaa;
rom[6975] = 12'haab;
rom[6976] = 12'hbbb;
rom[6977] = 12'habb;
rom[6978] = 12'haab;
rom[6979] = 12'haaa;
rom[6980] = 12'h9aa;
rom[6981] = 12'h99a;
rom[6982] = 12'h999;
rom[6983] = 12'h999;
rom[6984] = 12'h888;
rom[6985] = 12'h777;
rom[6986] = 12'h766;
rom[6987] = 12'h666;
rom[6988] = 12'h666;
rom[6989] = 12'h666;
rom[6990] = 12'h655;
rom[6991] = 12'h655;
rom[6992] = 12'h666;
rom[6993] = 12'h555;
rom[6994] = 12'h555;
rom[6995] = 12'h555;
rom[6996] = 12'h666;
rom[6997] = 12'h777;
rom[6998] = 12'h888;
rom[6999] = 12'h999;
rom[7000] = 12'h888;
rom[7001] = 12'h888;
rom[7002] = 12'h888;
rom[7003] = 12'h777;
rom[7004] = 12'h666;
rom[7005] = 12'h555;
rom[7006] = 12'h444;
rom[7007] = 12'h444;
rom[7008] = 12'h444;
rom[7009] = 12'h333;
rom[7010] = 12'h333;
rom[7011] = 12'h444;
rom[7012] = 12'h333;
rom[7013] = 12'h333;
rom[7014] = 12'h222;
rom[7015] = 12'h222;
rom[7016] = 12'h111;
rom[7017] = 12'h111;
rom[7018] = 12'h  0;
rom[7019] = 12'h  0;
rom[7020] = 12'h  0;
rom[7021] = 12'h  0;
rom[7022] = 12'h  0;
rom[7023] = 12'h  0;
rom[7024] = 12'h  0;
rom[7025] = 12'h  0;
rom[7026] = 12'h  0;
rom[7027] = 12'h  0;
rom[7028] = 12'h  0;
rom[7029] = 12'h  0;
rom[7030] = 12'h  0;
rom[7031] = 12'h  0;
rom[7032] = 12'h  0;
rom[7033] = 12'h  0;
rom[7034] = 12'h  0;
rom[7035] = 12'h  0;
rom[7036] = 12'h  0;
rom[7037] = 12'h  0;
rom[7038] = 12'h111;
rom[7039] = 12'h111;
rom[7040] = 12'h111;
rom[7041] = 12'h111;
rom[7042] = 12'h222;
rom[7043] = 12'h222;
rom[7044] = 12'h222;
rom[7045] = 12'h222;
rom[7046] = 12'h111;
rom[7047] = 12'h111;
rom[7048] = 12'h111;
rom[7049] = 12'h222;
rom[7050] = 12'h222;
rom[7051] = 12'h333;
rom[7052] = 12'h333;
rom[7053] = 12'h333;
rom[7054] = 12'h222;
rom[7055] = 12'h222;
rom[7056] = 12'h222;
rom[7057] = 12'h222;
rom[7058] = 12'h222;
rom[7059] = 12'h222;
rom[7060] = 12'h222;
rom[7061] = 12'h222;
rom[7062] = 12'h222;
rom[7063] = 12'h222;
rom[7064] = 12'h111;
rom[7065] = 12'h111;
rom[7066] = 12'h111;
rom[7067] = 12'h111;
rom[7068] = 12'h  0;
rom[7069] = 12'h  0;
rom[7070] = 12'h  0;
rom[7071] = 12'h  0;
rom[7072] = 12'h  0;
rom[7073] = 12'h  0;
rom[7074] = 12'h  0;
rom[7075] = 12'h  0;
rom[7076] = 12'h  0;
rom[7077] = 12'h  0;
rom[7078] = 12'h  0;
rom[7079] = 12'h  0;
rom[7080] = 12'h  0;
rom[7081] = 12'h  0;
rom[7082] = 12'h  0;
rom[7083] = 12'h  0;
rom[7084] = 12'h  0;
rom[7085] = 12'h  0;
rom[7086] = 12'h  0;
rom[7087] = 12'h  0;
rom[7088] = 12'h  0;
rom[7089] = 12'h  0;
rom[7090] = 12'h  0;
rom[7091] = 12'h  0;
rom[7092] = 12'h  0;
rom[7093] = 12'h  0;
rom[7094] = 12'h  0;
rom[7095] = 12'h  0;
rom[7096] = 12'h  0;
rom[7097] = 12'h  0;
rom[7098] = 12'h  0;
rom[7099] = 12'h  0;
rom[7100] = 12'h111;
rom[7101] = 12'h111;
rom[7102] = 12'h  0;
rom[7103] = 12'h  0;
rom[7104] = 12'h  0;
rom[7105] = 12'h  0;
rom[7106] = 12'h  0;
rom[7107] = 12'h  0;
rom[7108] = 12'h  0;
rom[7109] = 12'h  0;
rom[7110] = 12'h  0;
rom[7111] = 12'h  0;
rom[7112] = 12'h  0;
rom[7113] = 12'h  0;
rom[7114] = 12'h  0;
rom[7115] = 12'h  0;
rom[7116] = 12'h  0;
rom[7117] = 12'h111;
rom[7118] = 12'h111;
rom[7119] = 12'h222;
rom[7120] = 12'h444;
rom[7121] = 12'h555;
rom[7122] = 12'h666;
rom[7123] = 12'h666;
rom[7124] = 12'h666;
rom[7125] = 12'h444;
rom[7126] = 12'h333;
rom[7127] = 12'h333;
rom[7128] = 12'h333;
rom[7129] = 12'h333;
rom[7130] = 12'h222;
rom[7131] = 12'h222;
rom[7132] = 12'h111;
rom[7133] = 12'h111;
rom[7134] = 12'h111;
rom[7135] = 12'h111;
rom[7136] = 12'h111;
rom[7137] = 12'h111;
rom[7138] = 12'h111;
rom[7139] = 12'h111;
rom[7140] = 12'h111;
rom[7141] = 12'h111;
rom[7142] = 12'h222;
rom[7143] = 12'h222;
rom[7144] = 12'h333;
rom[7145] = 12'h222;
rom[7146] = 12'h222;
rom[7147] = 12'h222;
rom[7148] = 12'h222;
rom[7149] = 12'h222;
rom[7150] = 12'h333;
rom[7151] = 12'h444;
rom[7152] = 12'h444;
rom[7153] = 12'h444;
rom[7154] = 12'h444;
rom[7155] = 12'h555;
rom[7156] = 12'h555;
rom[7157] = 12'h666;
rom[7158] = 12'h666;
rom[7159] = 12'h666;
rom[7160] = 12'h555;
rom[7161] = 12'h555;
rom[7162] = 12'h444;
rom[7163] = 12'h444;
rom[7164] = 12'h444;
rom[7165] = 12'h444;
rom[7166] = 12'h444;
rom[7167] = 12'h444;
rom[7168] = 12'h444;
rom[7169] = 12'h555;
rom[7170] = 12'h555;
rom[7171] = 12'h555;
rom[7172] = 12'h555;
rom[7173] = 12'h444;
rom[7174] = 12'h444;
rom[7175] = 12'h444;
rom[7176] = 12'h444;
rom[7177] = 12'h444;
rom[7178] = 12'h444;
rom[7179] = 12'h444;
rom[7180] = 12'h444;
rom[7181] = 12'h444;
rom[7182] = 12'h444;
rom[7183] = 12'h555;
rom[7184] = 12'h555;
rom[7185] = 12'h666;
rom[7186] = 12'h666;
rom[7187] = 12'h666;
rom[7188] = 12'h777;
rom[7189] = 12'h777;
rom[7190] = 12'h777;
rom[7191] = 12'h777;
rom[7192] = 12'h888;
rom[7193] = 12'h999;
rom[7194] = 12'h999;
rom[7195] = 12'haaa;
rom[7196] = 12'haaa;
rom[7197] = 12'h999;
rom[7198] = 12'h999;
rom[7199] = 12'h999;
rom[7200] = 12'h666;
rom[7201] = 12'h666;
rom[7202] = 12'h666;
rom[7203] = 12'h555;
rom[7204] = 12'h555;
rom[7205] = 12'h444;
rom[7206] = 12'h444;
rom[7207] = 12'h333;
rom[7208] = 12'h333;
rom[7209] = 12'h333;
rom[7210] = 12'h222;
rom[7211] = 12'h222;
rom[7212] = 12'h222;
rom[7213] = 12'h222;
rom[7214] = 12'h222;
rom[7215] = 12'h111;
rom[7216] = 12'h222;
rom[7217] = 12'h111;
rom[7218] = 12'h111;
rom[7219] = 12'h111;
rom[7220] = 12'h111;
rom[7221] = 12'h111;
rom[7222] = 12'h111;
rom[7223] = 12'h111;
rom[7224] = 12'h111;
rom[7225] = 12'h111;
rom[7226] = 12'h111;
rom[7227] = 12'h  0;
rom[7228] = 12'h  0;
rom[7229] = 12'h  0;
rom[7230] = 12'h111;
rom[7231] = 12'h111;
rom[7232] = 12'h111;
rom[7233] = 12'h111;
rom[7234] = 12'h111;
rom[7235] = 12'h111;
rom[7236] = 12'h111;
rom[7237] = 12'h111;
rom[7238] = 12'h111;
rom[7239] = 12'h111;
rom[7240] = 12'h111;
rom[7241] = 12'h  0;
rom[7242] = 12'h  0;
rom[7243] = 12'h  0;
rom[7244] = 12'h  0;
rom[7245] = 12'h  0;
rom[7246] = 12'h  0;
rom[7247] = 12'h  0;
rom[7248] = 12'h  0;
rom[7249] = 12'h  0;
rom[7250] = 12'h  0;
rom[7251] = 12'h  0;
rom[7252] = 12'h  0;
rom[7253] = 12'h  0;
rom[7254] = 12'h  0;
rom[7255] = 12'h111;
rom[7256] = 12'h  0;
rom[7257] = 12'h  0;
rom[7258] = 12'h  0;
rom[7259] = 12'h111;
rom[7260] = 12'h111;
rom[7261] = 12'h111;
rom[7262] = 12'h111;
rom[7263] = 12'h111;
rom[7264] = 12'h111;
rom[7265] = 12'h111;
rom[7266] = 12'h111;
rom[7267] = 12'h111;
rom[7268] = 12'h111;
rom[7269] = 12'h111;
rom[7270] = 12'h111;
rom[7271] = 12'h111;
rom[7272] = 12'h  0;
rom[7273] = 12'h  0;
rom[7274] = 12'h111;
rom[7275] = 12'h111;
rom[7276] = 12'h111;
rom[7277] = 12'h111;
rom[7278] = 12'h111;
rom[7279] = 12'h111;
rom[7280] = 12'h111;
rom[7281] = 12'h111;
rom[7282] = 12'h111;
rom[7283] = 12'h111;
rom[7284] = 12'h111;
rom[7285] = 12'h111;
rom[7286] = 12'h111;
rom[7287] = 12'h111;
rom[7288] = 12'h  0;
rom[7289] = 12'h  0;
rom[7290] = 12'h111;
rom[7291] = 12'h111;
rom[7292] = 12'h222;
rom[7293] = 12'h222;
rom[7294] = 12'h333;
rom[7295] = 12'h444;
rom[7296] = 12'h444;
rom[7297] = 12'h444;
rom[7298] = 12'h333;
rom[7299] = 12'h333;
rom[7300] = 12'h233;
rom[7301] = 12'h233;
rom[7302] = 12'h333;
rom[7303] = 12'h333;
rom[7304] = 12'h444;
rom[7305] = 12'h444;
rom[7306] = 12'h555;
rom[7307] = 12'h655;
rom[7308] = 12'h655;
rom[7309] = 12'h544;
rom[7310] = 12'h544;
rom[7311] = 12'h544;
rom[7312] = 12'h643;
rom[7313] = 12'h643;
rom[7314] = 12'h642;
rom[7315] = 12'h642;
rom[7316] = 12'h853;
rom[7317] = 12'h963;
rom[7318] = 12'ha74;
rom[7319] = 12'ha74;
rom[7320] = 12'hb74;
rom[7321] = 12'hb84;
rom[7322] = 12'hb84;
rom[7323] = 12'ha73;
rom[7324] = 12'h963;
rom[7325] = 12'h952;
rom[7326] = 12'h841;
rom[7327] = 12'h731;
rom[7328] = 12'h631;
rom[7329] = 12'h521;
rom[7330] = 12'h520;
rom[7331] = 12'h510;
rom[7332] = 12'h510;
rom[7333] = 12'h510;
rom[7334] = 12'h520;
rom[7335] = 12'h520;
rom[7336] = 12'h520;
rom[7337] = 12'h520;
rom[7338] = 12'h520;
rom[7339] = 12'h520;
rom[7340] = 12'h520;
rom[7341] = 12'h620;
rom[7342] = 12'h620;
rom[7343] = 12'h620;
rom[7344] = 12'h621;
rom[7345] = 12'h620;
rom[7346] = 12'h620;
rom[7347] = 12'h620;
rom[7348] = 12'h620;
rom[7349] = 12'h620;
rom[7350] = 12'h621;
rom[7351] = 12'h621;
rom[7352] = 12'h521;
rom[7353] = 12'h521;
rom[7354] = 12'h520;
rom[7355] = 12'h521;
rom[7356] = 12'h521;
rom[7357] = 12'h521;
rom[7358] = 12'h521;
rom[7359] = 12'h521;
rom[7360] = 12'h531;
rom[7361] = 12'h532;
rom[7362] = 12'h543;
rom[7363] = 12'h643;
rom[7364] = 12'h754;
rom[7365] = 12'h765;
rom[7366] = 12'h866;
rom[7367] = 12'h876;
rom[7368] = 12'h877;
rom[7369] = 12'h988;
rom[7370] = 12'h988;
rom[7371] = 12'h999;
rom[7372] = 12'h988;
rom[7373] = 12'h988;
rom[7374] = 12'h999;
rom[7375] = 12'ha9a;
rom[7376] = 12'haaa;
rom[7377] = 12'haab;
rom[7378] = 12'haab;
rom[7379] = 12'haaa;
rom[7380] = 12'haaa;
rom[7381] = 12'haaa;
rom[7382] = 12'haaa;
rom[7383] = 12'haaa;
rom[7384] = 12'h999;
rom[7385] = 12'h888;
rom[7386] = 12'h877;
rom[7387] = 12'h777;
rom[7388] = 12'h777;
rom[7389] = 12'h766;
rom[7390] = 12'h666;
rom[7391] = 12'h666;
rom[7392] = 12'h666;
rom[7393] = 12'h666;
rom[7394] = 12'h555;
rom[7395] = 12'h555;
rom[7396] = 12'h666;
rom[7397] = 12'h777;
rom[7398] = 12'h888;
rom[7399] = 12'h999;
rom[7400] = 12'h999;
rom[7401] = 12'h888;
rom[7402] = 12'h888;
rom[7403] = 12'h888;
rom[7404] = 12'h777;
rom[7405] = 12'h555;
rom[7406] = 12'h444;
rom[7407] = 12'h444;
rom[7408] = 12'h444;
rom[7409] = 12'h333;
rom[7410] = 12'h333;
rom[7411] = 12'h444;
rom[7412] = 12'h333;
rom[7413] = 12'h333;
rom[7414] = 12'h222;
rom[7415] = 12'h222;
rom[7416] = 12'h111;
rom[7417] = 12'h111;
rom[7418] = 12'h111;
rom[7419] = 12'h  0;
rom[7420] = 12'h  0;
rom[7421] = 12'h  0;
rom[7422] = 12'h  0;
rom[7423] = 12'h  0;
rom[7424] = 12'h  0;
rom[7425] = 12'h  0;
rom[7426] = 12'h  0;
rom[7427] = 12'h  0;
rom[7428] = 12'h  0;
rom[7429] = 12'h  0;
rom[7430] = 12'h  0;
rom[7431] = 12'h  0;
rom[7432] = 12'h  0;
rom[7433] = 12'h  0;
rom[7434] = 12'h  0;
rom[7435] = 12'h  0;
rom[7436] = 12'h  0;
rom[7437] = 12'h111;
rom[7438] = 12'h111;
rom[7439] = 12'h111;
rom[7440] = 12'h222;
rom[7441] = 12'h222;
rom[7442] = 12'h222;
rom[7443] = 12'h222;
rom[7444] = 12'h222;
rom[7445] = 12'h222;
rom[7446] = 12'h222;
rom[7447] = 12'h111;
rom[7448] = 12'h222;
rom[7449] = 12'h222;
rom[7450] = 12'h333;
rom[7451] = 12'h333;
rom[7452] = 12'h333;
rom[7453] = 12'h333;
rom[7454] = 12'h222;
rom[7455] = 12'h222;
rom[7456] = 12'h222;
rom[7457] = 12'h222;
rom[7458] = 12'h222;
rom[7459] = 12'h222;
rom[7460] = 12'h222;
rom[7461] = 12'h222;
rom[7462] = 12'h222;
rom[7463] = 12'h222;
rom[7464] = 12'h111;
rom[7465] = 12'h111;
rom[7466] = 12'h111;
rom[7467] = 12'h111;
rom[7468] = 12'h  0;
rom[7469] = 12'h  0;
rom[7470] = 12'h  0;
rom[7471] = 12'h  0;
rom[7472] = 12'h  0;
rom[7473] = 12'h  0;
rom[7474] = 12'h  0;
rom[7475] = 12'h  0;
rom[7476] = 12'h  0;
rom[7477] = 12'h  0;
rom[7478] = 12'h  0;
rom[7479] = 12'h  0;
rom[7480] = 12'h  0;
rom[7481] = 12'h  0;
rom[7482] = 12'h  0;
rom[7483] = 12'h  0;
rom[7484] = 12'h  0;
rom[7485] = 12'h  0;
rom[7486] = 12'h  0;
rom[7487] = 12'h  0;
rom[7488] = 12'h  0;
rom[7489] = 12'h  0;
rom[7490] = 12'h  0;
rom[7491] = 12'h  0;
rom[7492] = 12'h  0;
rom[7493] = 12'h  0;
rom[7494] = 12'h  0;
rom[7495] = 12'h  0;
rom[7496] = 12'h  0;
rom[7497] = 12'h  0;
rom[7498] = 12'h  0;
rom[7499] = 12'h  0;
rom[7500] = 12'h111;
rom[7501] = 12'h111;
rom[7502] = 12'h  0;
rom[7503] = 12'h  0;
rom[7504] = 12'h  0;
rom[7505] = 12'h  0;
rom[7506] = 12'h  0;
rom[7507] = 12'h  0;
rom[7508] = 12'h  0;
rom[7509] = 12'h  0;
rom[7510] = 12'h  0;
rom[7511] = 12'h  0;
rom[7512] = 12'h  0;
rom[7513] = 12'h  0;
rom[7514] = 12'h  0;
rom[7515] = 12'h  0;
rom[7516] = 12'h  0;
rom[7517] = 12'h111;
rom[7518] = 12'h222;
rom[7519] = 12'h222;
rom[7520] = 12'h555;
rom[7521] = 12'h555;
rom[7522] = 12'h666;
rom[7523] = 12'h777;
rom[7524] = 12'h666;
rom[7525] = 12'h444;
rom[7526] = 12'h333;
rom[7527] = 12'h333;
rom[7528] = 12'h333;
rom[7529] = 12'h333;
rom[7530] = 12'h222;
rom[7531] = 12'h222;
rom[7532] = 12'h111;
rom[7533] = 12'h111;
rom[7534] = 12'h111;
rom[7535] = 12'h111;
rom[7536] = 12'h111;
rom[7537] = 12'h111;
rom[7538] = 12'h111;
rom[7539] = 12'h111;
rom[7540] = 12'h  0;
rom[7541] = 12'h111;
rom[7542] = 12'h222;
rom[7543] = 12'h333;
rom[7544] = 12'h333;
rom[7545] = 12'h222;
rom[7546] = 12'h111;
rom[7547] = 12'h222;
rom[7548] = 12'h222;
rom[7549] = 12'h222;
rom[7550] = 12'h333;
rom[7551] = 12'h444;
rom[7552] = 12'h444;
rom[7553] = 12'h444;
rom[7554] = 12'h555;
rom[7555] = 12'h555;
rom[7556] = 12'h555;
rom[7557] = 12'h555;
rom[7558] = 12'h555;
rom[7559] = 12'h555;
rom[7560] = 12'h555;
rom[7561] = 12'h555;
rom[7562] = 12'h444;
rom[7563] = 12'h444;
rom[7564] = 12'h444;
rom[7565] = 12'h444;
rom[7566] = 12'h444;
rom[7567] = 12'h444;
rom[7568] = 12'h555;
rom[7569] = 12'h555;
rom[7570] = 12'h555;
rom[7571] = 12'h555;
rom[7572] = 12'h444;
rom[7573] = 12'h444;
rom[7574] = 12'h333;
rom[7575] = 12'h444;
rom[7576] = 12'h444;
rom[7577] = 12'h444;
rom[7578] = 12'h444;
rom[7579] = 12'h444;
rom[7580] = 12'h444;
rom[7581] = 12'h444;
rom[7582] = 12'h444;
rom[7583] = 12'h555;
rom[7584] = 12'h555;
rom[7585] = 12'h666;
rom[7586] = 12'h666;
rom[7587] = 12'h777;
rom[7588] = 12'h777;
rom[7589] = 12'h777;
rom[7590] = 12'h777;
rom[7591] = 12'h777;
rom[7592] = 12'h888;
rom[7593] = 12'h888;
rom[7594] = 12'h999;
rom[7595] = 12'haaa;
rom[7596] = 12'haaa;
rom[7597] = 12'h999;
rom[7598] = 12'h999;
rom[7599] = 12'h999;
rom[7600] = 12'h555;
rom[7601] = 12'h555;
rom[7602] = 12'h444;
rom[7603] = 12'h444;
rom[7604] = 12'h444;
rom[7605] = 12'h333;
rom[7606] = 12'h333;
rom[7607] = 12'h333;
rom[7608] = 12'h222;
rom[7609] = 12'h222;
rom[7610] = 12'h222;
rom[7611] = 12'h222;
rom[7612] = 12'h222;
rom[7613] = 12'h222;
rom[7614] = 12'h111;
rom[7615] = 12'h111;
rom[7616] = 12'h111;
rom[7617] = 12'h111;
rom[7618] = 12'h111;
rom[7619] = 12'h111;
rom[7620] = 12'h111;
rom[7621] = 12'h111;
rom[7622] = 12'h111;
rom[7623] = 12'h111;
rom[7624] = 12'h111;
rom[7625] = 12'h111;
rom[7626] = 12'h111;
rom[7627] = 12'h  0;
rom[7628] = 12'h  0;
rom[7629] = 12'h  0;
rom[7630] = 12'h  0;
rom[7631] = 12'h  0;
rom[7632] = 12'h111;
rom[7633] = 12'h111;
rom[7634] = 12'h111;
rom[7635] = 12'h111;
rom[7636] = 12'h111;
rom[7637] = 12'h111;
rom[7638] = 12'h111;
rom[7639] = 12'h111;
rom[7640] = 12'h111;
rom[7641] = 12'h111;
rom[7642] = 12'h111;
rom[7643] = 12'h  0;
rom[7644] = 12'h  0;
rom[7645] = 12'h  0;
rom[7646] = 12'h  0;
rom[7647] = 12'h  0;
rom[7648] = 12'h  0;
rom[7649] = 12'h  0;
rom[7650] = 12'h  0;
rom[7651] = 12'h  0;
rom[7652] = 12'h  0;
rom[7653] = 12'h  0;
rom[7654] = 12'h  0;
rom[7655] = 12'h111;
rom[7656] = 12'h  0;
rom[7657] = 12'h  0;
rom[7658] = 12'h111;
rom[7659] = 12'h111;
rom[7660] = 12'h111;
rom[7661] = 12'h111;
rom[7662] = 12'h111;
rom[7663] = 12'h111;
rom[7664] = 12'h111;
rom[7665] = 12'h111;
rom[7666] = 12'h111;
rom[7667] = 12'h111;
rom[7668] = 12'h111;
rom[7669] = 12'h111;
rom[7670] = 12'h111;
rom[7671] = 12'h111;
rom[7672] = 12'h111;
rom[7673] = 12'h111;
rom[7674] = 12'h111;
rom[7675] = 12'h111;
rom[7676] = 12'h111;
rom[7677] = 12'h111;
rom[7678] = 12'h111;
rom[7679] = 12'h111;
rom[7680] = 12'h111;
rom[7681] = 12'h111;
rom[7682] = 12'h111;
rom[7683] = 12'h111;
rom[7684] = 12'h111;
rom[7685] = 12'h111;
rom[7686] = 12'h  0;
rom[7687] = 12'h  0;
rom[7688] = 12'h  0;
rom[7689] = 12'h111;
rom[7690] = 12'h111;
rom[7691] = 12'h222;
rom[7692] = 12'h222;
rom[7693] = 12'h333;
rom[7694] = 12'h333;
rom[7695] = 12'h333;
rom[7696] = 12'h333;
rom[7697] = 12'h222;
rom[7698] = 12'h222;
rom[7699] = 12'h222;
rom[7700] = 12'h222;
rom[7701] = 12'h222;
rom[7702] = 12'h333;
rom[7703] = 12'h333;
rom[7704] = 12'h444;
rom[7705] = 12'h444;
rom[7706] = 12'h544;
rom[7707] = 12'h545;
rom[7708] = 12'h544;
rom[7709] = 12'h444;
rom[7710] = 12'h433;
rom[7711] = 12'h533;
rom[7712] = 12'h533;
rom[7713] = 12'h532;
rom[7714] = 12'h532;
rom[7715] = 12'h642;
rom[7716] = 12'h752;
rom[7717] = 12'h963;
rom[7718] = 12'ha74;
rom[7719] = 12'hb74;
rom[7720] = 12'hb74;
rom[7721] = 12'hb84;
rom[7722] = 12'hb74;
rom[7723] = 12'ha63;
rom[7724] = 12'h952;
rom[7725] = 12'h841;
rom[7726] = 12'h731;
rom[7727] = 12'h630;
rom[7728] = 12'h520;
rom[7729] = 12'h510;
rom[7730] = 12'h510;
rom[7731] = 12'h510;
rom[7732] = 12'h510;
rom[7733] = 12'h510;
rom[7734] = 12'h510;
rom[7735] = 12'h510;
rom[7736] = 12'h510;
rom[7737] = 12'h510;
rom[7738] = 12'h510;
rom[7739] = 12'h510;
rom[7740] = 12'h610;
rom[7741] = 12'h610;
rom[7742] = 12'h610;
rom[7743] = 12'h610;
rom[7744] = 12'h620;
rom[7745] = 12'h620;
rom[7746] = 12'h620;
rom[7747] = 12'h620;
rom[7748] = 12'h620;
rom[7749] = 12'h620;
rom[7750] = 12'h621;
rom[7751] = 12'h621;
rom[7752] = 12'h621;
rom[7753] = 12'h521;
rom[7754] = 12'h521;
rom[7755] = 12'h521;
rom[7756] = 12'h521;
rom[7757] = 12'h521;
rom[7758] = 12'h521;
rom[7759] = 12'h521;
rom[7760] = 12'h410;
rom[7761] = 12'h420;
rom[7762] = 12'h421;
rom[7763] = 12'h421;
rom[7764] = 12'h532;
rom[7765] = 12'h532;
rom[7766] = 12'h643;
rom[7767] = 12'h644;
rom[7768] = 12'h765;
rom[7769] = 12'h876;
rom[7770] = 12'h988;
rom[7771] = 12'h988;
rom[7772] = 12'h988;
rom[7773] = 12'h988;
rom[7774] = 12'h988;
rom[7775] = 12'h988;
rom[7776] = 12'h999;
rom[7777] = 12'h999;
rom[7778] = 12'h999;
rom[7779] = 12'h9aa;
rom[7780] = 12'h999;
rom[7781] = 12'h999;
rom[7782] = 12'haaa;
rom[7783] = 12'haaa;
rom[7784] = 12'h999;
rom[7785] = 12'h999;
rom[7786] = 12'h999;
rom[7787] = 12'h888;
rom[7788] = 12'h888;
rom[7789] = 12'h777;
rom[7790] = 12'h777;
rom[7791] = 12'h777;
rom[7792] = 12'h777;
rom[7793] = 12'h666;
rom[7794] = 12'h666;
rom[7795] = 12'h666;
rom[7796] = 12'h666;
rom[7797] = 12'h777;
rom[7798] = 12'h888;
rom[7799] = 12'h999;
rom[7800] = 12'h999;
rom[7801] = 12'h888;
rom[7802] = 12'h888;
rom[7803] = 12'h888;
rom[7804] = 12'h777;
rom[7805] = 12'h555;
rom[7806] = 12'h444;
rom[7807] = 12'h444;
rom[7808] = 12'h444;
rom[7809] = 12'h333;
rom[7810] = 12'h333;
rom[7811] = 12'h444;
rom[7812] = 12'h333;
rom[7813] = 12'h222;
rom[7814] = 12'h222;
rom[7815] = 12'h222;
rom[7816] = 12'h111;
rom[7817] = 12'h111;
rom[7818] = 12'h111;
rom[7819] = 12'h111;
rom[7820] = 12'h  0;
rom[7821] = 12'h  0;
rom[7822] = 12'h  0;
rom[7823] = 12'h  0;
rom[7824] = 12'h  0;
rom[7825] = 12'h  0;
rom[7826] = 12'h  0;
rom[7827] = 12'h  0;
rom[7828] = 12'h  0;
rom[7829] = 12'h  0;
rom[7830] = 12'h  0;
rom[7831] = 12'h  0;
rom[7832] = 12'h  0;
rom[7833] = 12'h  0;
rom[7834] = 12'h  0;
rom[7835] = 12'h111;
rom[7836] = 12'h111;
rom[7837] = 12'h111;
rom[7838] = 12'h111;
rom[7839] = 12'h222;
rom[7840] = 12'h222;
rom[7841] = 12'h222;
rom[7842] = 12'h222;
rom[7843] = 12'h222;
rom[7844] = 12'h222;
rom[7845] = 12'h222;
rom[7846] = 12'h222;
rom[7847] = 12'h222;
rom[7848] = 12'h222;
rom[7849] = 12'h333;
rom[7850] = 12'h333;
rom[7851] = 12'h333;
rom[7852] = 12'h333;
rom[7853] = 12'h333;
rom[7854] = 12'h222;
rom[7855] = 12'h222;
rom[7856] = 12'h222;
rom[7857] = 12'h222;
rom[7858] = 12'h222;
rom[7859] = 12'h222;
rom[7860] = 12'h222;
rom[7861] = 12'h222;
rom[7862] = 12'h222;
rom[7863] = 12'h222;
rom[7864] = 12'h111;
rom[7865] = 12'h111;
rom[7866] = 12'h111;
rom[7867] = 12'h111;
rom[7868] = 12'h  0;
rom[7869] = 12'h  0;
rom[7870] = 12'h  0;
rom[7871] = 12'h  0;
rom[7872] = 12'h  0;
rom[7873] = 12'h  0;
rom[7874] = 12'h  0;
rom[7875] = 12'h  0;
rom[7876] = 12'h  0;
rom[7877] = 12'h  0;
rom[7878] = 12'h  0;
rom[7879] = 12'h  0;
rom[7880] = 12'h  0;
rom[7881] = 12'h  0;
rom[7882] = 12'h  0;
rom[7883] = 12'h  0;
rom[7884] = 12'h  0;
rom[7885] = 12'h  0;
rom[7886] = 12'h  0;
rom[7887] = 12'h  0;
rom[7888] = 12'h  0;
rom[7889] = 12'h  0;
rom[7890] = 12'h  0;
rom[7891] = 12'h  0;
rom[7892] = 12'h  0;
rom[7893] = 12'h  0;
rom[7894] = 12'h  0;
rom[7895] = 12'h  0;
rom[7896] = 12'h  0;
rom[7897] = 12'h  0;
rom[7898] = 12'h  0;
rom[7899] = 12'h  0;
rom[7900] = 12'h111;
rom[7901] = 12'h111;
rom[7902] = 12'h  0;
rom[7903] = 12'h  0;
rom[7904] = 12'h  0;
rom[7905] = 12'h  0;
rom[7906] = 12'h  0;
rom[7907] = 12'h  0;
rom[7908] = 12'h  0;
rom[7909] = 12'h  0;
rom[7910] = 12'h  0;
rom[7911] = 12'h  0;
rom[7912] = 12'h  0;
rom[7913] = 12'h  0;
rom[7914] = 12'h  0;
rom[7915] = 12'h  0;
rom[7916] = 12'h  0;
rom[7917] = 12'h111;
rom[7918] = 12'h222;
rom[7919] = 12'h333;
rom[7920] = 12'h555;
rom[7921] = 12'h555;
rom[7922] = 12'h666;
rom[7923] = 12'h777;
rom[7924] = 12'h666;
rom[7925] = 12'h444;
rom[7926] = 12'h333;
rom[7927] = 12'h444;
rom[7928] = 12'h333;
rom[7929] = 12'h333;
rom[7930] = 12'h222;
rom[7931] = 12'h222;
rom[7932] = 12'h111;
rom[7933] = 12'h111;
rom[7934] = 12'h111;
rom[7935] = 12'h111;
rom[7936] = 12'h111;
rom[7937] = 12'h111;
rom[7938] = 12'h111;
rom[7939] = 12'h111;
rom[7940] = 12'h111;
rom[7941] = 12'h111;
rom[7942] = 12'h222;
rom[7943] = 12'h222;
rom[7944] = 12'h222;
rom[7945] = 12'h111;
rom[7946] = 12'h111;
rom[7947] = 12'h222;
rom[7948] = 12'h222;
rom[7949] = 12'h222;
rom[7950] = 12'h333;
rom[7951] = 12'h444;
rom[7952] = 12'h444;
rom[7953] = 12'h444;
rom[7954] = 12'h555;
rom[7955] = 12'h555;
rom[7956] = 12'h555;
rom[7957] = 12'h555;
rom[7958] = 12'h555;
rom[7959] = 12'h555;
rom[7960] = 12'h555;
rom[7961] = 12'h444;
rom[7962] = 12'h444;
rom[7963] = 12'h444;
rom[7964] = 12'h444;
rom[7965] = 12'h444;
rom[7966] = 12'h555;
rom[7967] = 12'h555;
rom[7968] = 12'h444;
rom[7969] = 12'h555;
rom[7970] = 12'h444;
rom[7971] = 12'h444;
rom[7972] = 12'h444;
rom[7973] = 12'h333;
rom[7974] = 12'h444;
rom[7975] = 12'h444;
rom[7976] = 12'h444;
rom[7977] = 12'h444;
rom[7978] = 12'h444;
rom[7979] = 12'h444;
rom[7980] = 12'h444;
rom[7981] = 12'h444;
rom[7982] = 12'h555;
rom[7983] = 12'h555;
rom[7984] = 12'h555;
rom[7985] = 12'h666;
rom[7986] = 12'h666;
rom[7987] = 12'h777;
rom[7988] = 12'h777;
rom[7989] = 12'h777;
rom[7990] = 12'h777;
rom[7991] = 12'h777;
rom[7992] = 12'h888;
rom[7993] = 12'h888;
rom[7994] = 12'h999;
rom[7995] = 12'h999;
rom[7996] = 12'haaa;
rom[7997] = 12'h999;
rom[7998] = 12'h999;
rom[7999] = 12'h999;
rom[8000] = 12'h444;
rom[8001] = 12'h444;
rom[8002] = 12'h333;
rom[8003] = 12'h333;
rom[8004] = 12'h333;
rom[8005] = 12'h333;
rom[8006] = 12'h333;
rom[8007] = 12'h222;
rom[8008] = 12'h222;
rom[8009] = 12'h222;
rom[8010] = 12'h222;
rom[8011] = 12'h222;
rom[8012] = 12'h222;
rom[8013] = 12'h222;
rom[8014] = 12'h111;
rom[8015] = 12'h111;
rom[8016] = 12'h111;
rom[8017] = 12'h111;
rom[8018] = 12'h111;
rom[8019] = 12'h111;
rom[8020] = 12'h111;
rom[8021] = 12'h111;
rom[8022] = 12'h111;
rom[8023] = 12'h111;
rom[8024] = 12'h111;
rom[8025] = 12'h111;
rom[8026] = 12'h111;
rom[8027] = 12'h  0;
rom[8028] = 12'h  0;
rom[8029] = 12'h  0;
rom[8030] = 12'h  0;
rom[8031] = 12'h  0;
rom[8032] = 12'h111;
rom[8033] = 12'h111;
rom[8034] = 12'h111;
rom[8035] = 12'h111;
rom[8036] = 12'h111;
rom[8037] = 12'h111;
rom[8038] = 12'h111;
rom[8039] = 12'h111;
rom[8040] = 12'h111;
rom[8041] = 12'h111;
rom[8042] = 12'h111;
rom[8043] = 12'h111;
rom[8044] = 12'h  0;
rom[8045] = 12'h  0;
rom[8046] = 12'h  0;
rom[8047] = 12'h  0;
rom[8048] = 12'h  0;
rom[8049] = 12'h  0;
rom[8050] = 12'h  0;
rom[8051] = 12'h111;
rom[8052] = 12'h111;
rom[8053] = 12'h111;
rom[8054] = 12'h111;
rom[8055] = 12'h111;
rom[8056] = 12'h111;
rom[8057] = 12'h111;
rom[8058] = 12'h111;
rom[8059] = 12'h111;
rom[8060] = 12'h111;
rom[8061] = 12'h111;
rom[8062] = 12'h111;
rom[8063] = 12'h111;
rom[8064] = 12'h111;
rom[8065] = 12'h111;
rom[8066] = 12'h111;
rom[8067] = 12'h111;
rom[8068] = 12'h111;
rom[8069] = 12'h111;
rom[8070] = 12'h111;
rom[8071] = 12'h111;
rom[8072] = 12'h111;
rom[8073] = 12'h111;
rom[8074] = 12'h111;
rom[8075] = 12'h111;
rom[8076] = 12'h111;
rom[8077] = 12'h111;
rom[8078] = 12'h111;
rom[8079] = 12'h111;
rom[8080] = 12'h111;
rom[8081] = 12'h111;
rom[8082] = 12'h111;
rom[8083] = 12'h111;
rom[8084] = 12'h111;
rom[8085] = 12'h111;
rom[8086] = 12'h111;
rom[8087] = 12'h111;
rom[8088] = 12'h111;
rom[8089] = 12'h111;
rom[8090] = 12'h222;
rom[8091] = 12'h222;
rom[8092] = 12'h333;
rom[8093] = 12'h333;
rom[8094] = 12'h222;
rom[8095] = 12'h222;
rom[8096] = 12'h111;
rom[8097] = 12'h111;
rom[8098] = 12'h111;
rom[8099] = 12'h122;
rom[8100] = 12'h222;
rom[8101] = 12'h233;
rom[8102] = 12'h333;
rom[8103] = 12'h333;
rom[8104] = 12'h444;
rom[8105] = 12'h444;
rom[8106] = 12'h444;
rom[8107] = 12'h444;
rom[8108] = 12'h433;
rom[8109] = 12'h433;
rom[8110] = 12'h433;
rom[8111] = 12'h433;
rom[8112] = 12'h422;
rom[8113] = 12'h421;
rom[8114] = 12'h521;
rom[8115] = 12'h531;
rom[8116] = 12'h641;
rom[8117] = 12'h852;
rom[8118] = 12'h963;
rom[8119] = 12'ha63;
rom[8120] = 12'hb74;
rom[8121] = 12'hc74;
rom[8122] = 12'hb74;
rom[8123] = 12'ha63;
rom[8124] = 12'h942;
rom[8125] = 12'h831;
rom[8126] = 12'h730;
rom[8127] = 12'h620;
rom[8128] = 12'h510;
rom[8129] = 12'h510;
rom[8130] = 12'h510;
rom[8131] = 12'h510;
rom[8132] = 12'h510;
rom[8133] = 12'h510;
rom[8134] = 12'h510;
rom[8135] = 12'h510;
rom[8136] = 12'h510;
rom[8137] = 12'h510;
rom[8138] = 12'h510;
rom[8139] = 12'h510;
rom[8140] = 12'h610;
rom[8141] = 12'h610;
rom[8142] = 12'h610;
rom[8143] = 12'h610;
rom[8144] = 12'h610;
rom[8145] = 12'h510;
rom[8146] = 12'h510;
rom[8147] = 12'h510;
rom[8148] = 12'h510;
rom[8149] = 12'h520;
rom[8150] = 12'h520;
rom[8151] = 12'h520;
rom[8152] = 12'h520;
rom[8153] = 12'h520;
rom[8154] = 12'h520;
rom[8155] = 12'h520;
rom[8156] = 12'h520;
rom[8157] = 12'h520;
rom[8158] = 12'h520;
rom[8159] = 12'h520;
rom[8160] = 12'h521;
rom[8161] = 12'h421;
rom[8162] = 12'h421;
rom[8163] = 12'h420;
rom[8164] = 12'h410;
rom[8165] = 12'h411;
rom[8166] = 12'h421;
rom[8167] = 12'h421;
rom[8168] = 12'h533;
rom[8169] = 12'h644;
rom[8170] = 12'h755;
rom[8171] = 12'h866;
rom[8172] = 12'h877;
rom[8173] = 12'h977;
rom[8174] = 12'h978;
rom[8175] = 12'h988;
rom[8176] = 12'h988;
rom[8177] = 12'h998;
rom[8178] = 12'h999;
rom[8179] = 12'h9a9;
rom[8180] = 12'haaa;
rom[8181] = 12'haaa;
rom[8182] = 12'haaa;
rom[8183] = 12'h999;
rom[8184] = 12'h999;
rom[8185] = 12'haaa;
rom[8186] = 12'haaa;
rom[8187] = 12'h999;
rom[8188] = 12'h989;
rom[8189] = 12'h888;
rom[8190] = 12'h888;
rom[8191] = 12'h888;
rom[8192] = 12'h777;
rom[8193] = 12'h777;
rom[8194] = 12'h666;
rom[8195] = 12'h777;
rom[8196] = 12'h777;
rom[8197] = 12'h777;
rom[8198] = 12'h888;
rom[8199] = 12'h888;
rom[8200] = 12'h999;
rom[8201] = 12'h888;
rom[8202] = 12'h888;
rom[8203] = 12'h888;
rom[8204] = 12'h777;
rom[8205] = 12'h666;
rom[8206] = 12'h555;
rom[8207] = 12'h444;
rom[8208] = 12'h444;
rom[8209] = 12'h333;
rom[8210] = 12'h444;
rom[8211] = 12'h444;
rom[8212] = 12'h333;
rom[8213] = 12'h222;
rom[8214] = 12'h222;
rom[8215] = 12'h222;
rom[8216] = 12'h111;
rom[8217] = 12'h111;
rom[8218] = 12'h111;
rom[8219] = 12'h111;
rom[8220] = 12'h111;
rom[8221] = 12'h  0;
rom[8222] = 12'h  0;
rom[8223] = 12'h111;
rom[8224] = 12'h  0;
rom[8225] = 12'h  0;
rom[8226] = 12'h  0;
rom[8227] = 12'h  0;
rom[8228] = 12'h  0;
rom[8229] = 12'h  0;
rom[8230] = 12'h  0;
rom[8231] = 12'h  0;
rom[8232] = 12'h  0;
rom[8233] = 12'h  0;
rom[8234] = 12'h111;
rom[8235] = 12'h111;
rom[8236] = 12'h111;
rom[8237] = 12'h222;
rom[8238] = 12'h222;
rom[8239] = 12'h222;
rom[8240] = 12'h222;
rom[8241] = 12'h222;
rom[8242] = 12'h222;
rom[8243] = 12'h222;
rom[8244] = 12'h222;
rom[8245] = 12'h222;
rom[8246] = 12'h222;
rom[8247] = 12'h222;
rom[8248] = 12'h333;
rom[8249] = 12'h333;
rom[8250] = 12'h333;
rom[8251] = 12'h333;
rom[8252] = 12'h333;
rom[8253] = 12'h222;
rom[8254] = 12'h222;
rom[8255] = 12'h222;
rom[8256] = 12'h222;
rom[8257] = 12'h222;
rom[8258] = 12'h222;
rom[8259] = 12'h222;
rom[8260] = 12'h222;
rom[8261] = 12'h222;
rom[8262] = 12'h222;
rom[8263] = 12'h222;
rom[8264] = 12'h222;
rom[8265] = 12'h111;
rom[8266] = 12'h111;
rom[8267] = 12'h111;
rom[8268] = 12'h  0;
rom[8269] = 12'h  0;
rom[8270] = 12'h  0;
rom[8271] = 12'h  0;
rom[8272] = 12'h  0;
rom[8273] = 12'h  0;
rom[8274] = 12'h  0;
rom[8275] = 12'h  0;
rom[8276] = 12'h  0;
rom[8277] = 12'h  0;
rom[8278] = 12'h  0;
rom[8279] = 12'h  0;
rom[8280] = 12'h  0;
rom[8281] = 12'h  0;
rom[8282] = 12'h  0;
rom[8283] = 12'h  0;
rom[8284] = 12'h  0;
rom[8285] = 12'h  0;
rom[8286] = 12'h  0;
rom[8287] = 12'h  0;
rom[8288] = 12'h  0;
rom[8289] = 12'h  0;
rom[8290] = 12'h  0;
rom[8291] = 12'h  0;
rom[8292] = 12'h  0;
rom[8293] = 12'h  0;
rom[8294] = 12'h  0;
rom[8295] = 12'h  0;
rom[8296] = 12'h  0;
rom[8297] = 12'h  0;
rom[8298] = 12'h  0;
rom[8299] = 12'h  0;
rom[8300] = 12'h111;
rom[8301] = 12'h111;
rom[8302] = 12'h  0;
rom[8303] = 12'h  0;
rom[8304] = 12'h  0;
rom[8305] = 12'h  0;
rom[8306] = 12'h  0;
rom[8307] = 12'h  0;
rom[8308] = 12'h  0;
rom[8309] = 12'h  0;
rom[8310] = 12'h  0;
rom[8311] = 12'h  0;
rom[8312] = 12'h  0;
rom[8313] = 12'h  0;
rom[8314] = 12'h  0;
rom[8315] = 12'h  0;
rom[8316] = 12'h111;
rom[8317] = 12'h111;
rom[8318] = 12'h222;
rom[8319] = 12'h333;
rom[8320] = 12'h555;
rom[8321] = 12'h666;
rom[8322] = 12'h666;
rom[8323] = 12'h777;
rom[8324] = 12'h555;
rom[8325] = 12'h444;
rom[8326] = 12'h333;
rom[8327] = 12'h444;
rom[8328] = 12'h444;
rom[8329] = 12'h333;
rom[8330] = 12'h222;
rom[8331] = 12'h111;
rom[8332] = 12'h111;
rom[8333] = 12'h111;
rom[8334] = 12'h111;
rom[8335] = 12'h  0;
rom[8336] = 12'h111;
rom[8337] = 12'h111;
rom[8338] = 12'h  0;
rom[8339] = 12'h111;
rom[8340] = 12'h111;
rom[8341] = 12'h222;
rom[8342] = 12'h222;
rom[8343] = 12'h222;
rom[8344] = 12'h111;
rom[8345] = 12'h111;
rom[8346] = 12'h222;
rom[8347] = 12'h222;
rom[8348] = 12'h222;
rom[8349] = 12'h333;
rom[8350] = 12'h333;
rom[8351] = 12'h333;
rom[8352] = 12'h444;
rom[8353] = 12'h444;
rom[8354] = 12'h555;
rom[8355] = 12'h555;
rom[8356] = 12'h555;
rom[8357] = 12'h555;
rom[8358] = 12'h555;
rom[8359] = 12'h555;
rom[8360] = 12'h555;
rom[8361] = 12'h444;
rom[8362] = 12'h444;
rom[8363] = 12'h444;
rom[8364] = 12'h444;
rom[8365] = 12'h555;
rom[8366] = 12'h555;
rom[8367] = 12'h555;
rom[8368] = 12'h444;
rom[8369] = 12'h444;
rom[8370] = 12'h333;
rom[8371] = 12'h333;
rom[8372] = 12'h333;
rom[8373] = 12'h444;
rom[8374] = 12'h444;
rom[8375] = 12'h444;
rom[8376] = 12'h444;
rom[8377] = 12'h444;
rom[8378] = 12'h444;
rom[8379] = 12'h444;
rom[8380] = 12'h444;
rom[8381] = 12'h555;
rom[8382] = 12'h555;
rom[8383] = 12'h555;
rom[8384] = 12'h666;
rom[8385] = 12'h666;
rom[8386] = 12'h777;
rom[8387] = 12'h777;
rom[8388] = 12'h777;
rom[8389] = 12'h777;
rom[8390] = 12'h777;
rom[8391] = 12'h777;
rom[8392] = 12'h888;
rom[8393] = 12'h888;
rom[8394] = 12'h999;
rom[8395] = 12'h999;
rom[8396] = 12'haaa;
rom[8397] = 12'haaa;
rom[8398] = 12'h999;
rom[8399] = 12'h999;
rom[8400] = 12'h444;
rom[8401] = 12'h444;
rom[8402] = 12'h333;
rom[8403] = 12'h333;
rom[8404] = 12'h333;
rom[8405] = 12'h333;
rom[8406] = 12'h222;
rom[8407] = 12'h222;
rom[8408] = 12'h222;
rom[8409] = 12'h222;
rom[8410] = 12'h222;
rom[8411] = 12'h222;
rom[8412] = 12'h222;
rom[8413] = 12'h222;
rom[8414] = 12'h222;
rom[8415] = 12'h222;
rom[8416] = 12'h111;
rom[8417] = 12'h111;
rom[8418] = 12'h111;
rom[8419] = 12'h111;
rom[8420] = 12'h111;
rom[8421] = 12'h111;
rom[8422] = 12'h111;
rom[8423] = 12'h111;
rom[8424] = 12'h111;
rom[8425] = 12'h111;
rom[8426] = 12'h111;
rom[8427] = 12'h111;
rom[8428] = 12'h  0;
rom[8429] = 12'h  0;
rom[8430] = 12'h  0;
rom[8431] = 12'h  0;
rom[8432] = 12'h111;
rom[8433] = 12'h111;
rom[8434] = 12'h111;
rom[8435] = 12'h111;
rom[8436] = 12'h111;
rom[8437] = 12'h111;
rom[8438] = 12'h111;
rom[8439] = 12'h111;
rom[8440] = 12'h111;
rom[8441] = 12'h111;
rom[8442] = 12'h111;
rom[8443] = 12'h111;
rom[8444] = 12'h111;
rom[8445] = 12'h111;
rom[8446] = 12'h  0;
rom[8447] = 12'h  0;
rom[8448] = 12'h  0;
rom[8449] = 12'h111;
rom[8450] = 12'h111;
rom[8451] = 12'h111;
rom[8452] = 12'h111;
rom[8453] = 12'h111;
rom[8454] = 12'h111;
rom[8455] = 12'h111;
rom[8456] = 12'h111;
rom[8457] = 12'h111;
rom[8458] = 12'h111;
rom[8459] = 12'h111;
rom[8460] = 12'h111;
rom[8461] = 12'h111;
rom[8462] = 12'h111;
rom[8463] = 12'h111;
rom[8464] = 12'h111;
rom[8465] = 12'h111;
rom[8466] = 12'h111;
rom[8467] = 12'h111;
rom[8468] = 12'h111;
rom[8469] = 12'h111;
rom[8470] = 12'h111;
rom[8471] = 12'h111;
rom[8472] = 12'h111;
rom[8473] = 12'h111;
rom[8474] = 12'h111;
rom[8475] = 12'h111;
rom[8476] = 12'h111;
rom[8477] = 12'h111;
rom[8478] = 12'h111;
rom[8479] = 12'h111;
rom[8480] = 12'h111;
rom[8481] = 12'h111;
rom[8482] = 12'h111;
rom[8483] = 12'h111;
rom[8484] = 12'h111;
rom[8485] = 12'h111;
rom[8486] = 12'h111;
rom[8487] = 12'h111;
rom[8488] = 12'h222;
rom[8489] = 12'h222;
rom[8490] = 12'h222;
rom[8491] = 12'h333;
rom[8492] = 12'h222;
rom[8493] = 12'h222;
rom[8494] = 12'h222;
rom[8495] = 12'h111;
rom[8496] = 12'h111;
rom[8497] = 12'h111;
rom[8498] = 12'h111;
rom[8499] = 12'h222;
rom[8500] = 12'h222;
rom[8501] = 12'h233;
rom[8502] = 12'h333;
rom[8503] = 12'h333;
rom[8504] = 12'h444;
rom[8505] = 12'h444;
rom[8506] = 12'h433;
rom[8507] = 12'h333;
rom[8508] = 12'h333;
rom[8509] = 12'h433;
rom[8510] = 12'h433;
rom[8511] = 12'h433;
rom[8512] = 12'h421;
rom[8513] = 12'h421;
rom[8514] = 12'h421;
rom[8515] = 12'h520;
rom[8516] = 12'h631;
rom[8517] = 12'h741;
rom[8518] = 12'h852;
rom[8519] = 12'h952;
rom[8520] = 12'hb73;
rom[8521] = 12'hb74;
rom[8522] = 12'hb73;
rom[8523] = 12'ha52;
rom[8524] = 12'h841;
rom[8525] = 12'h730;
rom[8526] = 12'h620;
rom[8527] = 12'h610;
rom[8528] = 12'h510;
rom[8529] = 12'h510;
rom[8530] = 12'h510;
rom[8531] = 12'h510;
rom[8532] = 12'h510;
rom[8533] = 12'h510;
rom[8534] = 12'h500;
rom[8535] = 12'h500;
rom[8536] = 12'h500;
rom[8537] = 12'h500;
rom[8538] = 12'h500;
rom[8539] = 12'h500;
rom[8540] = 12'h610;
rom[8541] = 12'h610;
rom[8542] = 12'h610;
rom[8543] = 12'h610;
rom[8544] = 12'h610;
rom[8545] = 12'h510;
rom[8546] = 12'h510;
rom[8547] = 12'h510;
rom[8548] = 12'h510;
rom[8549] = 12'h510;
rom[8550] = 12'h510;
rom[8551] = 12'h510;
rom[8552] = 12'h510;
rom[8553] = 12'h510;
rom[8554] = 12'h410;
rom[8555] = 12'h410;
rom[8556] = 12'h410;
rom[8557] = 12'h410;
rom[8558] = 12'h410;
rom[8559] = 12'h410;
rom[8560] = 12'h420;
rom[8561] = 12'h420;
rom[8562] = 12'h410;
rom[8563] = 12'h410;
rom[8564] = 12'h410;
rom[8565] = 12'h410;
rom[8566] = 12'h410;
rom[8567] = 12'h411;
rom[8568] = 12'h421;
rom[8569] = 12'h421;
rom[8570] = 12'h422;
rom[8571] = 12'h533;
rom[8572] = 12'h754;
rom[8573] = 12'h866;
rom[8574] = 12'h977;
rom[8575] = 12'h987;
rom[8576] = 12'h988;
rom[8577] = 12'h998;
rom[8578] = 12'h998;
rom[8579] = 12'h9a9;
rom[8580] = 12'haa9;
rom[8581] = 12'haaa;
rom[8582] = 12'haaa;
rom[8583] = 12'h9a9;
rom[8584] = 12'h999;
rom[8585] = 12'haaa;
rom[8586] = 12'haaa;
rom[8587] = 12'h99a;
rom[8588] = 12'h999;
rom[8589] = 12'h888;
rom[8590] = 12'h878;
rom[8591] = 12'h878;
rom[8592] = 12'h777;
rom[8593] = 12'h777;
rom[8594] = 12'h777;
rom[8595] = 12'h777;
rom[8596] = 12'h777;
rom[8597] = 12'h777;
rom[8598] = 12'h888;
rom[8599] = 12'h888;
rom[8600] = 12'h999;
rom[8601] = 12'h888;
rom[8602] = 12'h888;
rom[8603] = 12'h888;
rom[8604] = 12'h888;
rom[8605] = 12'h666;
rom[8606] = 12'h555;
rom[8607] = 12'h555;
rom[8608] = 12'h444;
rom[8609] = 12'h444;
rom[8610] = 12'h444;
rom[8611] = 12'h444;
rom[8612] = 12'h333;
rom[8613] = 12'h333;
rom[8614] = 12'h333;
rom[8615] = 12'h222;
rom[8616] = 12'h222;
rom[8617] = 12'h111;
rom[8618] = 12'h111;
rom[8619] = 12'h111;
rom[8620] = 12'h111;
rom[8621] = 12'h  0;
rom[8622] = 12'h  0;
rom[8623] = 12'h111;
rom[8624] = 12'h111;
rom[8625] = 12'h  0;
rom[8626] = 12'h  0;
rom[8627] = 12'h  0;
rom[8628] = 12'h  0;
rom[8629] = 12'h  0;
rom[8630] = 12'h  0;
rom[8631] = 12'h  0;
rom[8632] = 12'h111;
rom[8633] = 12'h111;
rom[8634] = 12'h111;
rom[8635] = 12'h111;
rom[8636] = 12'h222;
rom[8637] = 12'h222;
rom[8638] = 12'h222;
rom[8639] = 12'h222;
rom[8640] = 12'h222;
rom[8641] = 12'h222;
rom[8642] = 12'h222;
rom[8643] = 12'h222;
rom[8644] = 12'h222;
rom[8645] = 12'h222;
rom[8646] = 12'h222;
rom[8647] = 12'h333;
rom[8648] = 12'h333;
rom[8649] = 12'h333;
rom[8650] = 12'h333;
rom[8651] = 12'h333;
rom[8652] = 12'h333;
rom[8653] = 12'h222;
rom[8654] = 12'h222;
rom[8655] = 12'h333;
rom[8656] = 12'h333;
rom[8657] = 12'h333;
rom[8658] = 12'h222;
rom[8659] = 12'h222;
rom[8660] = 12'h222;
rom[8661] = 12'h222;
rom[8662] = 12'h222;
rom[8663] = 12'h111;
rom[8664] = 12'h222;
rom[8665] = 12'h222;
rom[8666] = 12'h111;
rom[8667] = 12'h111;
rom[8668] = 12'h  0;
rom[8669] = 12'h  0;
rom[8670] = 12'h  0;
rom[8671] = 12'h  0;
rom[8672] = 12'h  0;
rom[8673] = 12'h  0;
rom[8674] = 12'h  0;
rom[8675] = 12'h  0;
rom[8676] = 12'h  0;
rom[8677] = 12'h  0;
rom[8678] = 12'h  0;
rom[8679] = 12'h  0;
rom[8680] = 12'h  0;
rom[8681] = 12'h  0;
rom[8682] = 12'h  0;
rom[8683] = 12'h  0;
rom[8684] = 12'h  0;
rom[8685] = 12'h  0;
rom[8686] = 12'h  0;
rom[8687] = 12'h  0;
rom[8688] = 12'h  0;
rom[8689] = 12'h  0;
rom[8690] = 12'h  0;
rom[8691] = 12'h  0;
rom[8692] = 12'h  0;
rom[8693] = 12'h  0;
rom[8694] = 12'h  0;
rom[8695] = 12'h  0;
rom[8696] = 12'h  0;
rom[8697] = 12'h  0;
rom[8698] = 12'h  0;
rom[8699] = 12'h  0;
rom[8700] = 12'h111;
rom[8701] = 12'h111;
rom[8702] = 12'h  0;
rom[8703] = 12'h  0;
rom[8704] = 12'h  0;
rom[8705] = 12'h  0;
rom[8706] = 12'h  0;
rom[8707] = 12'h  0;
rom[8708] = 12'h  0;
rom[8709] = 12'h  0;
rom[8710] = 12'h  0;
rom[8711] = 12'h  0;
rom[8712] = 12'h  0;
rom[8713] = 12'h  0;
rom[8714] = 12'h  0;
rom[8715] = 12'h111;
rom[8716] = 12'h111;
rom[8717] = 12'h111;
rom[8718] = 12'h333;
rom[8719] = 12'h444;
rom[8720] = 12'h555;
rom[8721] = 12'h666;
rom[8722] = 12'h777;
rom[8723] = 12'h666;
rom[8724] = 12'h555;
rom[8725] = 12'h444;
rom[8726] = 12'h444;
rom[8727] = 12'h444;
rom[8728] = 12'h444;
rom[8729] = 12'h333;
rom[8730] = 12'h222;
rom[8731] = 12'h111;
rom[8732] = 12'h111;
rom[8733] = 12'h111;
rom[8734] = 12'h111;
rom[8735] = 12'h  0;
rom[8736] = 12'h111;
rom[8737] = 12'h111;
rom[8738] = 12'h111;
rom[8739] = 12'h111;
rom[8740] = 12'h222;
rom[8741] = 12'h222;
rom[8742] = 12'h222;
rom[8743] = 12'h111;
rom[8744] = 12'h111;
rom[8745] = 12'h222;
rom[8746] = 12'h222;
rom[8747] = 12'h222;
rom[8748] = 12'h222;
rom[8749] = 12'h333;
rom[8750] = 12'h333;
rom[8751] = 12'h333;
rom[8752] = 12'h444;
rom[8753] = 12'h444;
rom[8754] = 12'h555;
rom[8755] = 12'h555;
rom[8756] = 12'h555;
rom[8757] = 12'h666;
rom[8758] = 12'h666;
rom[8759] = 12'h555;
rom[8760] = 12'h555;
rom[8761] = 12'h444;
rom[8762] = 12'h444;
rom[8763] = 12'h444;
rom[8764] = 12'h555;
rom[8765] = 12'h555;
rom[8766] = 12'h555;
rom[8767] = 12'h555;
rom[8768] = 12'h444;
rom[8769] = 12'h444;
rom[8770] = 12'h333;
rom[8771] = 12'h333;
rom[8772] = 12'h333;
rom[8773] = 12'h444;
rom[8774] = 12'h444;
rom[8775] = 12'h444;
rom[8776] = 12'h444;
rom[8777] = 12'h444;
rom[8778] = 12'h444;
rom[8779] = 12'h444;
rom[8780] = 12'h444;
rom[8781] = 12'h555;
rom[8782] = 12'h555;
rom[8783] = 12'h666;
rom[8784] = 12'h777;
rom[8785] = 12'h777;
rom[8786] = 12'h777;
rom[8787] = 12'h777;
rom[8788] = 12'h777;
rom[8789] = 12'h777;
rom[8790] = 12'h777;
rom[8791] = 12'h777;
rom[8792] = 12'h888;
rom[8793] = 12'h888;
rom[8794] = 12'h999;
rom[8795] = 12'h999;
rom[8796] = 12'haaa;
rom[8797] = 12'haaa;
rom[8798] = 12'haaa;
rom[8799] = 12'h999;
rom[8800] = 12'h444;
rom[8801] = 12'h444;
rom[8802] = 12'h333;
rom[8803] = 12'h333;
rom[8804] = 12'h333;
rom[8805] = 12'h222;
rom[8806] = 12'h222;
rom[8807] = 12'h222;
rom[8808] = 12'h222;
rom[8809] = 12'h222;
rom[8810] = 12'h111;
rom[8811] = 12'h111;
rom[8812] = 12'h222;
rom[8813] = 12'h222;
rom[8814] = 12'h222;
rom[8815] = 12'h222;
rom[8816] = 12'h111;
rom[8817] = 12'h111;
rom[8818] = 12'h111;
rom[8819] = 12'h111;
rom[8820] = 12'h111;
rom[8821] = 12'h111;
rom[8822] = 12'h111;
rom[8823] = 12'h111;
rom[8824] = 12'h111;
rom[8825] = 12'h111;
rom[8826] = 12'h111;
rom[8827] = 12'h111;
rom[8828] = 12'h111;
rom[8829] = 12'h111;
rom[8830] = 12'h111;
rom[8831] = 12'h111;
rom[8832] = 12'h111;
rom[8833] = 12'h111;
rom[8834] = 12'h111;
rom[8835] = 12'h111;
rom[8836] = 12'h111;
rom[8837] = 12'h111;
rom[8838] = 12'h111;
rom[8839] = 12'h111;
rom[8840] = 12'h111;
rom[8841] = 12'h111;
rom[8842] = 12'h111;
rom[8843] = 12'h111;
rom[8844] = 12'h111;
rom[8845] = 12'h111;
rom[8846] = 12'h111;
rom[8847] = 12'h111;
rom[8848] = 12'h111;
rom[8849] = 12'h111;
rom[8850] = 12'h111;
rom[8851] = 12'h111;
rom[8852] = 12'h111;
rom[8853] = 12'h111;
rom[8854] = 12'h111;
rom[8855] = 12'h111;
rom[8856] = 12'h111;
rom[8857] = 12'h111;
rom[8858] = 12'h111;
rom[8859] = 12'h222;
rom[8860] = 12'h222;
rom[8861] = 12'h222;
rom[8862] = 12'h222;
rom[8863] = 12'h222;
rom[8864] = 12'h111;
rom[8865] = 12'h111;
rom[8866] = 12'h222;
rom[8867] = 12'h222;
rom[8868] = 12'h222;
rom[8869] = 12'h222;
rom[8870] = 12'h111;
rom[8871] = 12'h111;
rom[8872] = 12'h111;
rom[8873] = 12'h111;
rom[8874] = 12'h111;
rom[8875] = 12'h111;
rom[8876] = 12'h111;
rom[8877] = 12'h111;
rom[8878] = 12'h111;
rom[8879] = 12'h111;
rom[8880] = 12'h111;
rom[8881] = 12'h111;
rom[8882] = 12'h111;
rom[8883] = 12'h111;
rom[8884] = 12'h111;
rom[8885] = 12'h111;
rom[8886] = 12'h111;
rom[8887] = 12'h222;
rom[8888] = 12'h222;
rom[8889] = 12'h222;
rom[8890] = 12'h222;
rom[8891] = 12'h222;
rom[8892] = 12'h222;
rom[8893] = 12'h111;
rom[8894] = 12'h111;
rom[8895] = 12'h111;
rom[8896] = 12'h111;
rom[8897] = 12'h111;
rom[8898] = 12'h111;
rom[8899] = 12'h222;
rom[8900] = 12'h222;
rom[8901] = 12'h233;
rom[8902] = 12'h333;
rom[8903] = 12'h333;
rom[8904] = 12'h333;
rom[8905] = 12'h333;
rom[8906] = 12'h333;
rom[8907] = 12'h322;
rom[8908] = 12'h322;
rom[8909] = 12'h322;
rom[8910] = 12'h322;
rom[8911] = 12'h322;
rom[8912] = 12'h311;
rom[8913] = 12'h310;
rom[8914] = 12'h410;
rom[8915] = 12'h410;
rom[8916] = 12'h520;
rom[8917] = 12'h731;
rom[8918] = 12'h841;
rom[8919] = 12'h952;
rom[8920] = 12'hb63;
rom[8921] = 12'hb63;
rom[8922] = 12'hb63;
rom[8923] = 12'ha52;
rom[8924] = 12'h831;
rom[8925] = 12'h720;
rom[8926] = 12'h620;
rom[8927] = 12'h610;
rom[8928] = 12'h500;
rom[8929] = 12'h500;
rom[8930] = 12'h500;
rom[8931] = 12'h500;
rom[8932] = 12'h500;
rom[8933] = 12'h500;
rom[8934] = 12'h500;
rom[8935] = 12'h500;
rom[8936] = 12'h500;
rom[8937] = 12'h500;
rom[8938] = 12'h500;
rom[8939] = 12'h500;
rom[8940] = 12'h500;
rom[8941] = 12'h610;
rom[8942] = 12'h610;
rom[8943] = 12'h610;
rom[8944] = 12'h610;
rom[8945] = 12'h610;
rom[8946] = 12'h510;
rom[8947] = 12'h510;
rom[8948] = 12'h510;
rom[8949] = 12'h510;
rom[8950] = 12'h510;
rom[8951] = 12'h410;
rom[8952] = 12'h410;
rom[8953] = 12'h410;
rom[8954] = 12'h410;
rom[8955] = 12'h410;
rom[8956] = 12'h410;
rom[8957] = 12'h410;
rom[8958] = 12'h410;
rom[8959] = 12'h410;
rom[8960] = 12'h410;
rom[8961] = 12'h410;
rom[8962] = 12'h410;
rom[8963] = 12'h410;
rom[8964] = 12'h410;
rom[8965] = 12'h410;
rom[8966] = 12'h410;
rom[8967] = 12'h411;
rom[8968] = 12'h410;
rom[8969] = 12'h410;
rom[8970] = 12'h410;
rom[8971] = 12'h421;
rom[8972] = 12'h532;
rom[8973] = 12'h644;
rom[8974] = 12'h855;
rom[8975] = 12'h866;
rom[8976] = 12'h876;
rom[8977] = 12'h776;
rom[8978] = 12'h887;
rom[8979] = 12'h998;
rom[8980] = 12'h998;
rom[8981] = 12'ha99;
rom[8982] = 12'haa9;
rom[8983] = 12'haaa;
rom[8984] = 12'haaa;
rom[8985] = 12'haaa;
rom[8986] = 12'h999;
rom[8987] = 12'h999;
rom[8988] = 12'h999;
rom[8989] = 12'h889;
rom[8990] = 12'h888;
rom[8991] = 12'h888;
rom[8992] = 12'h777;
rom[8993] = 12'h777;
rom[8994] = 12'h777;
rom[8995] = 12'h777;
rom[8996] = 12'h777;
rom[8997] = 12'h777;
rom[8998] = 12'h888;
rom[8999] = 12'h888;
rom[9000] = 12'h999;
rom[9001] = 12'h888;
rom[9002] = 12'h888;
rom[9003] = 12'h999;
rom[9004] = 12'h888;
rom[9005] = 12'h777;
rom[9006] = 12'h666;
rom[9007] = 12'h555;
rom[9008] = 12'h555;
rom[9009] = 12'h444;
rom[9010] = 12'h444;
rom[9011] = 12'h444;
rom[9012] = 12'h333;
rom[9013] = 12'h333;
rom[9014] = 12'h333;
rom[9015] = 12'h333;
rom[9016] = 12'h222;
rom[9017] = 12'h111;
rom[9018] = 12'h111;
rom[9019] = 12'h111;
rom[9020] = 12'h111;
rom[9021] = 12'h111;
rom[9022] = 12'h111;
rom[9023] = 12'h111;
rom[9024] = 12'h111;
rom[9025] = 12'h111;
rom[9026] = 12'h111;
rom[9027] = 12'h  0;
rom[9028] = 12'h  0;
rom[9029] = 12'h  0;
rom[9030] = 12'h111;
rom[9031] = 12'h111;
rom[9032] = 12'h111;
rom[9033] = 12'h111;
rom[9034] = 12'h111;
rom[9035] = 12'h111;
rom[9036] = 12'h222;
rom[9037] = 12'h222;
rom[9038] = 12'h222;
rom[9039] = 12'h222;
rom[9040] = 12'h333;
rom[9041] = 12'h333;
rom[9042] = 12'h222;
rom[9043] = 12'h222;
rom[9044] = 12'h222;
rom[9045] = 12'h222;
rom[9046] = 12'h333;
rom[9047] = 12'h333;
rom[9048] = 12'h333;
rom[9049] = 12'h333;
rom[9050] = 12'h333;
rom[9051] = 12'h333;
rom[9052] = 12'h333;
rom[9053] = 12'h333;
rom[9054] = 12'h333;
rom[9055] = 12'h333;
rom[9056] = 12'h333;
rom[9057] = 12'h333;
rom[9058] = 12'h222;
rom[9059] = 12'h222;
rom[9060] = 12'h222;
rom[9061] = 12'h222;
rom[9062] = 12'h222;
rom[9063] = 12'h222;
rom[9064] = 12'h222;
rom[9065] = 12'h111;
rom[9066] = 12'h111;
rom[9067] = 12'h111;
rom[9068] = 12'h  0;
rom[9069] = 12'h  0;
rom[9070] = 12'h  0;
rom[9071] = 12'h  0;
rom[9072] = 12'h  0;
rom[9073] = 12'h  0;
rom[9074] = 12'h  0;
rom[9075] = 12'h  0;
rom[9076] = 12'h  0;
rom[9077] = 12'h  0;
rom[9078] = 12'h  0;
rom[9079] = 12'h  0;
rom[9080] = 12'h  0;
rom[9081] = 12'h  0;
rom[9082] = 12'h  0;
rom[9083] = 12'h  0;
rom[9084] = 12'h  0;
rom[9085] = 12'h  0;
rom[9086] = 12'h  0;
rom[9087] = 12'h  0;
rom[9088] = 12'h  0;
rom[9089] = 12'h  0;
rom[9090] = 12'h  0;
rom[9091] = 12'h  0;
rom[9092] = 12'h  0;
rom[9093] = 12'h  0;
rom[9094] = 12'h  0;
rom[9095] = 12'h  0;
rom[9096] = 12'h  0;
rom[9097] = 12'h  0;
rom[9098] = 12'h  0;
rom[9099] = 12'h  0;
rom[9100] = 12'h111;
rom[9101] = 12'h111;
rom[9102] = 12'h  0;
rom[9103] = 12'h  0;
rom[9104] = 12'h  0;
rom[9105] = 12'h  0;
rom[9106] = 12'h  0;
rom[9107] = 12'h  0;
rom[9108] = 12'h  0;
rom[9109] = 12'h  0;
rom[9110] = 12'h  0;
rom[9111] = 12'h  0;
rom[9112] = 12'h  0;
rom[9113] = 12'h  0;
rom[9114] = 12'h  0;
rom[9115] = 12'h111;
rom[9116] = 12'h111;
rom[9117] = 12'h111;
rom[9118] = 12'h333;
rom[9119] = 12'h555;
rom[9120] = 12'h555;
rom[9121] = 12'h777;
rom[9122] = 12'h777;
rom[9123] = 12'h666;
rom[9124] = 12'h444;
rom[9125] = 12'h444;
rom[9126] = 12'h444;
rom[9127] = 12'h444;
rom[9128] = 12'h333;
rom[9129] = 12'h333;
rom[9130] = 12'h222;
rom[9131] = 12'h111;
rom[9132] = 12'h111;
rom[9133] = 12'h111;
rom[9134] = 12'h111;
rom[9135] = 12'h  0;
rom[9136] = 12'h111;
rom[9137] = 12'h111;
rom[9138] = 12'h111;
rom[9139] = 12'h222;
rom[9140] = 12'h222;
rom[9141] = 12'h222;
rom[9142] = 12'h111;
rom[9143] = 12'h111;
rom[9144] = 12'h111;
rom[9145] = 12'h111;
rom[9146] = 12'h222;
rom[9147] = 12'h222;
rom[9148] = 12'h222;
rom[9149] = 12'h222;
rom[9150] = 12'h333;
rom[9151] = 12'h333;
rom[9152] = 12'h444;
rom[9153] = 12'h444;
rom[9154] = 12'h555;
rom[9155] = 12'h555;
rom[9156] = 12'h666;
rom[9157] = 12'h666;
rom[9158] = 12'h555;
rom[9159] = 12'h555;
rom[9160] = 12'h555;
rom[9161] = 12'h444;
rom[9162] = 12'h444;
rom[9163] = 12'h444;
rom[9164] = 12'h555;
rom[9165] = 12'h555;
rom[9166] = 12'h444;
rom[9167] = 12'h444;
rom[9168] = 12'h444;
rom[9169] = 12'h444;
rom[9170] = 12'h333;
rom[9171] = 12'h333;
rom[9172] = 12'h333;
rom[9173] = 12'h444;
rom[9174] = 12'h444;
rom[9175] = 12'h444;
rom[9176] = 12'h333;
rom[9177] = 12'h444;
rom[9178] = 12'h444;
rom[9179] = 12'h444;
rom[9180] = 12'h555;
rom[9181] = 12'h666;
rom[9182] = 12'h666;
rom[9183] = 12'h777;
rom[9184] = 12'h777;
rom[9185] = 12'h777;
rom[9186] = 12'h777;
rom[9187] = 12'h777;
rom[9188] = 12'h777;
rom[9189] = 12'h777;
rom[9190] = 12'h777;
rom[9191] = 12'h777;
rom[9192] = 12'h777;
rom[9193] = 12'h888;
rom[9194] = 12'h999;
rom[9195] = 12'h999;
rom[9196] = 12'haaa;
rom[9197] = 12'haaa;
rom[9198] = 12'haaa;
rom[9199] = 12'h999;
rom[9200] = 12'h444;
rom[9201] = 12'h333;
rom[9202] = 12'h333;
rom[9203] = 12'h333;
rom[9204] = 12'h333;
rom[9205] = 12'h222;
rom[9206] = 12'h222;
rom[9207] = 12'h222;
rom[9208] = 12'h222;
rom[9209] = 12'h111;
rom[9210] = 12'h111;
rom[9211] = 12'h111;
rom[9212] = 12'h111;
rom[9213] = 12'h222;
rom[9214] = 12'h111;
rom[9215] = 12'h111;
rom[9216] = 12'h111;
rom[9217] = 12'h111;
rom[9218] = 12'h111;
rom[9219] = 12'h111;
rom[9220] = 12'h  0;
rom[9221] = 12'h  0;
rom[9222] = 12'h111;
rom[9223] = 12'h111;
rom[9224] = 12'h111;
rom[9225] = 12'h111;
rom[9226] = 12'h111;
rom[9227] = 12'h111;
rom[9228] = 12'h111;
rom[9229] = 12'h111;
rom[9230] = 12'h111;
rom[9231] = 12'h111;
rom[9232] = 12'h111;
rom[9233] = 12'h111;
rom[9234] = 12'h111;
rom[9235] = 12'h111;
rom[9236] = 12'h111;
rom[9237] = 12'h111;
rom[9238] = 12'h111;
rom[9239] = 12'h111;
rom[9240] = 12'h111;
rom[9241] = 12'h111;
rom[9242] = 12'h111;
rom[9243] = 12'h222;
rom[9244] = 12'h222;
rom[9245] = 12'h222;
rom[9246] = 12'h222;
rom[9247] = 12'h222;
rom[9248] = 12'h111;
rom[9249] = 12'h111;
rom[9250] = 12'h111;
rom[9251] = 12'h  0;
rom[9252] = 12'h  0;
rom[9253] = 12'h111;
rom[9254] = 12'h111;
rom[9255] = 12'h222;
rom[9256] = 12'h111;
rom[9257] = 12'h222;
rom[9258] = 12'h222;
rom[9259] = 12'h222;
rom[9260] = 12'h222;
rom[9261] = 12'h222;
rom[9262] = 12'h222;
rom[9263] = 12'h222;
rom[9264] = 12'h222;
rom[9265] = 12'h222;
rom[9266] = 12'h222;
rom[9267] = 12'h222;
rom[9268] = 12'h222;
rom[9269] = 12'h222;
rom[9270] = 12'h222;
rom[9271] = 12'h222;
rom[9272] = 12'h111;
rom[9273] = 12'h111;
rom[9274] = 12'h111;
rom[9275] = 12'h111;
rom[9276] = 12'h111;
rom[9277] = 12'h111;
rom[9278] = 12'h111;
rom[9279] = 12'h111;
rom[9280] = 12'h111;
rom[9281] = 12'h111;
rom[9282] = 12'h111;
rom[9283] = 12'h111;
rom[9284] = 12'h111;
rom[9285] = 12'h222;
rom[9286] = 12'h222;
rom[9287] = 12'h222;
rom[9288] = 12'h222;
rom[9289] = 12'h222;
rom[9290] = 12'h222;
rom[9291] = 12'h111;
rom[9292] = 12'h111;
rom[9293] = 12'h111;
rom[9294] = 12'h111;
rom[9295] = 12'h  0;
rom[9296] = 12'h111;
rom[9297] = 12'h111;
rom[9298] = 12'h111;
rom[9299] = 12'h111;
rom[9300] = 12'h222;
rom[9301] = 12'h222;
rom[9302] = 12'h233;
rom[9303] = 12'h333;
rom[9304] = 12'h333;
rom[9305] = 12'h333;
rom[9306] = 12'h333;
rom[9307] = 12'h322;
rom[9308] = 12'h322;
rom[9309] = 12'h322;
rom[9310] = 12'h322;
rom[9311] = 12'h211;
rom[9312] = 12'h310;
rom[9313] = 12'h310;
rom[9314] = 12'h310;
rom[9315] = 12'h410;
rom[9316] = 12'h510;
rom[9317] = 12'h620;
rom[9318] = 12'h841;
rom[9319] = 12'h941;
rom[9320] = 12'hb63;
rom[9321] = 12'hb63;
rom[9322] = 12'hb63;
rom[9323] = 12'ha42;
rom[9324] = 12'h830;
rom[9325] = 12'h720;
rom[9326] = 12'h710;
rom[9327] = 12'h610;
rom[9328] = 12'h500;
rom[9329] = 12'h500;
rom[9330] = 12'h500;
rom[9331] = 12'h400;
rom[9332] = 12'h400;
rom[9333] = 12'h500;
rom[9334] = 12'h500;
rom[9335] = 12'h500;
rom[9336] = 12'h500;
rom[9337] = 12'h500;
rom[9338] = 12'h500;
rom[9339] = 12'h500;
rom[9340] = 12'h500;
rom[9341] = 12'h500;
rom[9342] = 12'h500;
rom[9343] = 12'h500;
rom[9344] = 12'h510;
rom[9345] = 12'h510;
rom[9346] = 12'h500;
rom[9347] = 12'h500;
rom[9348] = 12'h500;
rom[9349] = 12'h410;
rom[9350] = 12'h410;
rom[9351] = 12'h410;
rom[9352] = 12'h410;
rom[9353] = 12'h410;
rom[9354] = 12'h410;
rom[9355] = 12'h410;
rom[9356] = 12'h410;
rom[9357] = 12'h410;
rom[9358] = 12'h410;
rom[9359] = 12'h410;
rom[9360] = 12'h410;
rom[9361] = 12'h410;
rom[9362] = 12'h410;
rom[9363] = 12'h410;
rom[9364] = 12'h410;
rom[9365] = 12'h300;
rom[9366] = 12'h400;
rom[9367] = 12'h410;
rom[9368] = 12'h410;
rom[9369] = 12'h410;
rom[9370] = 12'h410;
rom[9371] = 12'h410;
rom[9372] = 12'h411;
rom[9373] = 12'h521;
rom[9374] = 12'h632;
rom[9375] = 12'h643;
rom[9376] = 12'h654;
rom[9377] = 12'h665;
rom[9378] = 12'h776;
rom[9379] = 12'h876;
rom[9380] = 12'h887;
rom[9381] = 12'h998;
rom[9382] = 12'haa9;
rom[9383] = 12'hbba;
rom[9384] = 12'hbbb;
rom[9385] = 12'haaa;
rom[9386] = 12'h999;
rom[9387] = 12'h999;
rom[9388] = 12'h99a;
rom[9389] = 12'h99a;
rom[9390] = 12'h99a;
rom[9391] = 12'h889;
rom[9392] = 12'h777;
rom[9393] = 12'h777;
rom[9394] = 12'h777;
rom[9395] = 12'h777;
rom[9396] = 12'h777;
rom[9397] = 12'h777;
rom[9398] = 12'h888;
rom[9399] = 12'h888;
rom[9400] = 12'h999;
rom[9401] = 12'h888;
rom[9402] = 12'h888;
rom[9403] = 12'h999;
rom[9404] = 12'h999;
rom[9405] = 12'h777;
rom[9406] = 12'h666;
rom[9407] = 12'h555;
rom[9408] = 12'h666;
rom[9409] = 12'h555;
rom[9410] = 12'h555;
rom[9411] = 12'h444;
rom[9412] = 12'h333;
rom[9413] = 12'h333;
rom[9414] = 12'h444;
rom[9415] = 12'h333;
rom[9416] = 12'h222;
rom[9417] = 12'h222;
rom[9418] = 12'h111;
rom[9419] = 12'h111;
rom[9420] = 12'h111;
rom[9421] = 12'h111;
rom[9422] = 12'h111;
rom[9423] = 12'h111;
rom[9424] = 12'h222;
rom[9425] = 12'h111;
rom[9426] = 12'h111;
rom[9427] = 12'h111;
rom[9428] = 12'h111;
rom[9429] = 12'h111;
rom[9430] = 12'h111;
rom[9431] = 12'h111;
rom[9432] = 12'h222;
rom[9433] = 12'h222;
rom[9434] = 12'h222;
rom[9435] = 12'h111;
rom[9436] = 12'h222;
rom[9437] = 12'h222;
rom[9438] = 12'h222;
rom[9439] = 12'h222;
rom[9440] = 12'h333;
rom[9441] = 12'h333;
rom[9442] = 12'h333;
rom[9443] = 12'h333;
rom[9444] = 12'h333;
rom[9445] = 12'h333;
rom[9446] = 12'h333;
rom[9447] = 12'h444;
rom[9448] = 12'h333;
rom[9449] = 12'h333;
rom[9450] = 12'h444;
rom[9451] = 12'h333;
rom[9452] = 12'h333;
rom[9453] = 12'h333;
rom[9454] = 12'h333;
rom[9455] = 12'h333;
rom[9456] = 12'h333;
rom[9457] = 12'h222;
rom[9458] = 12'h222;
rom[9459] = 12'h222;
rom[9460] = 12'h222;
rom[9461] = 12'h222;
rom[9462] = 12'h222;
rom[9463] = 12'h222;
rom[9464] = 12'h222;
rom[9465] = 12'h111;
rom[9466] = 12'h111;
rom[9467] = 12'h  0;
rom[9468] = 12'h  0;
rom[9469] = 12'h  0;
rom[9470] = 12'h  0;
rom[9471] = 12'h  0;
rom[9472] = 12'h  0;
rom[9473] = 12'h  0;
rom[9474] = 12'h  0;
rom[9475] = 12'h  0;
rom[9476] = 12'h  0;
rom[9477] = 12'h  0;
rom[9478] = 12'h  0;
rom[9479] = 12'h  0;
rom[9480] = 12'h  0;
rom[9481] = 12'h  0;
rom[9482] = 12'h  0;
rom[9483] = 12'h  0;
rom[9484] = 12'h  0;
rom[9485] = 12'h  0;
rom[9486] = 12'h  0;
rom[9487] = 12'h  0;
rom[9488] = 12'h  0;
rom[9489] = 12'h  0;
rom[9490] = 12'h  0;
rom[9491] = 12'h  0;
rom[9492] = 12'h  0;
rom[9493] = 12'h  0;
rom[9494] = 12'h  0;
rom[9495] = 12'h  0;
rom[9496] = 12'h  0;
rom[9497] = 12'h  0;
rom[9498] = 12'h  0;
rom[9499] = 12'h  0;
rom[9500] = 12'h111;
rom[9501] = 12'h111;
rom[9502] = 12'h  0;
rom[9503] = 12'h  0;
rom[9504] = 12'h  0;
rom[9505] = 12'h  0;
rom[9506] = 12'h  0;
rom[9507] = 12'h  0;
rom[9508] = 12'h  0;
rom[9509] = 12'h  0;
rom[9510] = 12'h  0;
rom[9511] = 12'h  0;
rom[9512] = 12'h  0;
rom[9513] = 12'h  0;
rom[9514] = 12'h  0;
rom[9515] = 12'h111;
rom[9516] = 12'h111;
rom[9517] = 12'h222;
rom[9518] = 12'h333;
rom[9519] = 12'h555;
rom[9520] = 12'h555;
rom[9521] = 12'h777;
rom[9522] = 12'h777;
rom[9523] = 12'h555;
rom[9524] = 12'h444;
rom[9525] = 12'h444;
rom[9526] = 12'h444;
rom[9527] = 12'h444;
rom[9528] = 12'h333;
rom[9529] = 12'h222;
rom[9530] = 12'h111;
rom[9531] = 12'h111;
rom[9532] = 12'h111;
rom[9533] = 12'h111;
rom[9534] = 12'h111;
rom[9535] = 12'h111;
rom[9536] = 12'h111;
rom[9537] = 12'h111;
rom[9538] = 12'h111;
rom[9539] = 12'h222;
rom[9540] = 12'h222;
rom[9541] = 12'h222;
rom[9542] = 12'h111;
rom[9543] = 12'h111;
rom[9544] = 12'h111;
rom[9545] = 12'h111;
rom[9546] = 12'h111;
rom[9547] = 12'h222;
rom[9548] = 12'h222;
rom[9549] = 12'h222;
rom[9550] = 12'h222;
rom[9551] = 12'h333;
rom[9552] = 12'h444;
rom[9553] = 12'h444;
rom[9554] = 12'h555;
rom[9555] = 12'h555;
rom[9556] = 12'h666;
rom[9557] = 12'h666;
rom[9558] = 12'h555;
rom[9559] = 12'h555;
rom[9560] = 12'h555;
rom[9561] = 12'h444;
rom[9562] = 12'h444;
rom[9563] = 12'h444;
rom[9564] = 12'h444;
rom[9565] = 12'h444;
rom[9566] = 12'h444;
rom[9567] = 12'h333;
rom[9568] = 12'h333;
rom[9569] = 12'h333;
rom[9570] = 12'h444;
rom[9571] = 12'h444;
rom[9572] = 12'h444;
rom[9573] = 12'h444;
rom[9574] = 12'h444;
rom[9575] = 12'h444;
rom[9576] = 12'h333;
rom[9577] = 12'h444;
rom[9578] = 12'h444;
rom[9579] = 12'h555;
rom[9580] = 12'h666;
rom[9581] = 12'h666;
rom[9582] = 12'h777;
rom[9583] = 12'h777;
rom[9584] = 12'h777;
rom[9585] = 12'h777;
rom[9586] = 12'h777;
rom[9587] = 12'h777;
rom[9588] = 12'h666;
rom[9589] = 12'h666;
rom[9590] = 12'h777;
rom[9591] = 12'h777;
rom[9592] = 12'h777;
rom[9593] = 12'h888;
rom[9594] = 12'h888;
rom[9595] = 12'h999;
rom[9596] = 12'haaa;
rom[9597] = 12'haaa;
rom[9598] = 12'haaa;
rom[9599] = 12'h999;
rom[9600] = 12'h333;
rom[9601] = 12'h333;
rom[9602] = 12'h333;
rom[9603] = 12'h333;
rom[9604] = 12'h333;
rom[9605] = 12'h333;
rom[9606] = 12'h222;
rom[9607] = 12'h222;
rom[9608] = 12'h222;
rom[9609] = 12'h222;
rom[9610] = 12'h222;
rom[9611] = 12'h111;
rom[9612] = 12'h111;
rom[9613] = 12'h111;
rom[9614] = 12'h111;
rom[9615] = 12'h111;
rom[9616] = 12'h111;
rom[9617] = 12'h111;
rom[9618] = 12'h111;
rom[9619] = 12'h111;
rom[9620] = 12'h111;
rom[9621] = 12'h  0;
rom[9622] = 12'h  0;
rom[9623] = 12'h  0;
rom[9624] = 12'h111;
rom[9625] = 12'h111;
rom[9626] = 12'h111;
rom[9627] = 12'h111;
rom[9628] = 12'h111;
rom[9629] = 12'h111;
rom[9630] = 12'h111;
rom[9631] = 12'h111;
rom[9632] = 12'h  0;
rom[9633] = 12'h111;
rom[9634] = 12'h111;
rom[9635] = 12'h111;
rom[9636] = 12'h111;
rom[9637] = 12'h111;
rom[9638] = 12'h111;
rom[9639] = 12'h111;
rom[9640] = 12'h111;
rom[9641] = 12'h111;
rom[9642] = 12'h111;
rom[9643] = 12'h111;
rom[9644] = 12'h111;
rom[9645] = 12'h222;
rom[9646] = 12'h222;
rom[9647] = 12'h222;
rom[9648] = 12'h333;
rom[9649] = 12'h222;
rom[9650] = 12'h222;
rom[9651] = 12'h111;
rom[9652] = 12'h111;
rom[9653] = 12'h111;
rom[9654] = 12'h111;
rom[9655] = 12'h111;
rom[9656] = 12'h111;
rom[9657] = 12'h222;
rom[9658] = 12'h222;
rom[9659] = 12'h333;
rom[9660] = 12'h333;
rom[9661] = 12'h333;
rom[9662] = 12'h222;
rom[9663] = 12'h222;
rom[9664] = 12'h222;
rom[9665] = 12'h222;
rom[9666] = 12'h222;
rom[9667] = 12'h222;
rom[9668] = 12'h222;
rom[9669] = 12'h222;
rom[9670] = 12'h222;
rom[9671] = 12'h222;
rom[9672] = 12'h222;
rom[9673] = 12'h222;
rom[9674] = 12'h111;
rom[9675] = 12'h111;
rom[9676] = 12'h111;
rom[9677] = 12'h111;
rom[9678] = 12'h111;
rom[9679] = 12'h111;
rom[9680] = 12'h111;
rom[9681] = 12'h111;
rom[9682] = 12'h222;
rom[9683] = 12'h222;
rom[9684] = 12'h222;
rom[9685] = 12'h222;
rom[9686] = 12'h222;
rom[9687] = 12'h222;
rom[9688] = 12'h222;
rom[9689] = 12'h222;
rom[9690] = 12'h111;
rom[9691] = 12'h111;
rom[9692] = 12'h111;
rom[9693] = 12'h  0;
rom[9694] = 12'h  0;
rom[9695] = 12'h  0;
rom[9696] = 12'h111;
rom[9697] = 12'h111;
rom[9698] = 12'h111;
rom[9699] = 12'h111;
rom[9700] = 12'h122;
rom[9701] = 12'h222;
rom[9702] = 12'h222;
rom[9703] = 12'h222;
rom[9704] = 12'h222;
rom[9705] = 12'h222;
rom[9706] = 12'h222;
rom[9707] = 12'h222;
rom[9708] = 12'h222;
rom[9709] = 12'h211;
rom[9710] = 12'h211;
rom[9711] = 12'h211;
rom[9712] = 12'h200;
rom[9713] = 12'h200;
rom[9714] = 12'h310;
rom[9715] = 12'h410;
rom[9716] = 12'h510;
rom[9717] = 12'h620;
rom[9718] = 12'h720;
rom[9719] = 12'h830;
rom[9720] = 12'ha52;
rom[9721] = 12'hb52;
rom[9722] = 12'hb53;
rom[9723] = 12'ha42;
rom[9724] = 12'h830;
rom[9725] = 12'h720;
rom[9726] = 12'h710;
rom[9727] = 12'h610;
rom[9728] = 12'h500;
rom[9729] = 12'h400;
rom[9730] = 12'h400;
rom[9731] = 12'h400;
rom[9732] = 12'h400;
rom[9733] = 12'h400;
rom[9734] = 12'h400;
rom[9735] = 12'h400;
rom[9736] = 12'h400;
rom[9737] = 12'h400;
rom[9738] = 12'h500;
rom[9739] = 12'h400;
rom[9740] = 12'h500;
rom[9741] = 12'h500;
rom[9742] = 12'h500;
rom[9743] = 12'h510;
rom[9744] = 12'h500;
rom[9745] = 12'h500;
rom[9746] = 12'h500;
rom[9747] = 12'h500;
rom[9748] = 12'h400;
rom[9749] = 12'h400;
rom[9750] = 12'h400;
rom[9751] = 12'h400;
rom[9752] = 12'h400;
rom[9753] = 12'h400;
rom[9754] = 12'h400;
rom[9755] = 12'h400;
rom[9756] = 12'h400;
rom[9757] = 12'h410;
rom[9758] = 12'h410;
rom[9759] = 12'h410;
rom[9760] = 12'h400;
rom[9761] = 12'h400;
rom[9762] = 12'h400;
rom[9763] = 12'h400;
rom[9764] = 12'h400;
rom[9765] = 12'h400;
rom[9766] = 12'h400;
rom[9767] = 12'h300;
rom[9768] = 12'h400;
rom[9769] = 12'h400;
rom[9770] = 12'h400;
rom[9771] = 12'h400;
rom[9772] = 12'h410;
rom[9773] = 12'h410;
rom[9774] = 12'h411;
rom[9775] = 12'h411;
rom[9776] = 12'h432;
rom[9777] = 12'h543;
rom[9778] = 12'h654;
rom[9779] = 12'h765;
rom[9780] = 12'h766;
rom[9781] = 12'h876;
rom[9782] = 12'h988;
rom[9783] = 12'ha99;
rom[9784] = 12'hbbb;
rom[9785] = 12'hbbb;
rom[9786] = 12'haaa;
rom[9787] = 12'haaa;
rom[9788] = 12'haaa;
rom[9789] = 12'haab;
rom[9790] = 12'h99a;
rom[9791] = 12'h899;
rom[9792] = 12'h888;
rom[9793] = 12'h888;
rom[9794] = 12'h888;
rom[9795] = 12'h777;
rom[9796] = 12'h777;
rom[9797] = 12'h777;
rom[9798] = 12'h888;
rom[9799] = 12'h888;
rom[9800] = 12'h999;
rom[9801] = 12'h999;
rom[9802] = 12'h888;
rom[9803] = 12'h999;
rom[9804] = 12'h999;
rom[9805] = 12'h888;
rom[9806] = 12'h666;
rom[9807] = 12'h666;
rom[9808] = 12'h666;
rom[9809] = 12'h555;
rom[9810] = 12'h555;
rom[9811] = 12'h444;
rom[9812] = 12'h444;
rom[9813] = 12'h444;
rom[9814] = 12'h444;
rom[9815] = 12'h444;
rom[9816] = 12'h222;
rom[9817] = 12'h222;
rom[9818] = 12'h222;
rom[9819] = 12'h222;
rom[9820] = 12'h222;
rom[9821] = 12'h222;
rom[9822] = 12'h222;
rom[9823] = 12'h222;
rom[9824] = 12'h111;
rom[9825] = 12'h111;
rom[9826] = 12'h111;
rom[9827] = 12'h111;
rom[9828] = 12'h111;
rom[9829] = 12'h111;
rom[9830] = 12'h222;
rom[9831] = 12'h222;
rom[9832] = 12'h333;
rom[9833] = 12'h222;
rom[9834] = 12'h111;
rom[9835] = 12'h222;
rom[9836] = 12'h222;
rom[9837] = 12'h333;
rom[9838] = 12'h333;
rom[9839] = 12'h333;
rom[9840] = 12'h333;
rom[9841] = 12'h333;
rom[9842] = 12'h333;
rom[9843] = 12'h333;
rom[9844] = 12'h444;
rom[9845] = 12'h555;
rom[9846] = 12'h444;
rom[9847] = 12'h444;
rom[9848] = 12'h444;
rom[9849] = 12'h444;
rom[9850] = 12'h333;
rom[9851] = 12'h333;
rom[9852] = 12'h333;
rom[9853] = 12'h333;
rom[9854] = 12'h333;
rom[9855] = 12'h333;
rom[9856] = 12'h222;
rom[9857] = 12'h222;
rom[9858] = 12'h222;
rom[9859] = 12'h222;
rom[9860] = 12'h222;
rom[9861] = 12'h222;
rom[9862] = 12'h222;
rom[9863] = 12'h222;
rom[9864] = 12'h111;
rom[9865] = 12'h111;
rom[9866] = 12'h111;
rom[9867] = 12'h  0;
rom[9868] = 12'h  0;
rom[9869] = 12'h  0;
rom[9870] = 12'h  0;
rom[9871] = 12'h  0;
rom[9872] = 12'h  0;
rom[9873] = 12'h  0;
rom[9874] = 12'h  0;
rom[9875] = 12'h  0;
rom[9876] = 12'h  0;
rom[9877] = 12'h  0;
rom[9878] = 12'h  0;
rom[9879] = 12'h  0;
rom[9880] = 12'h  0;
rom[9881] = 12'h  0;
rom[9882] = 12'h  0;
rom[9883] = 12'h  0;
rom[9884] = 12'h  0;
rom[9885] = 12'h  0;
rom[9886] = 12'h  0;
rom[9887] = 12'h  0;
rom[9888] = 12'h  0;
rom[9889] = 12'h  0;
rom[9890] = 12'h  0;
rom[9891] = 12'h  0;
rom[9892] = 12'h  0;
rom[9893] = 12'h  0;
rom[9894] = 12'h  0;
rom[9895] = 12'h  0;
rom[9896] = 12'h  0;
rom[9897] = 12'h  0;
rom[9898] = 12'h  0;
rom[9899] = 12'h  0;
rom[9900] = 12'h111;
rom[9901] = 12'h111;
rom[9902] = 12'h  0;
rom[9903] = 12'h  0;
rom[9904] = 12'h  0;
rom[9905] = 12'h  0;
rom[9906] = 12'h  0;
rom[9907] = 12'h  0;
rom[9908] = 12'h  0;
rom[9909] = 12'h  0;
rom[9910] = 12'h  0;
rom[9911] = 12'h  0;
rom[9912] = 12'h  0;
rom[9913] = 12'h  0;
rom[9914] = 12'h  0;
rom[9915] = 12'h111;
rom[9916] = 12'h111;
rom[9917] = 12'h222;
rom[9918] = 12'h444;
rom[9919] = 12'h666;
rom[9920] = 12'h777;
rom[9921] = 12'h777;
rom[9922] = 12'h666;
rom[9923] = 12'h555;
rom[9924] = 12'h444;
rom[9925] = 12'h444;
rom[9926] = 12'h444;
rom[9927] = 12'h444;
rom[9928] = 12'h333;
rom[9929] = 12'h222;
rom[9930] = 12'h111;
rom[9931] = 12'h111;
rom[9932] = 12'h111;
rom[9933] = 12'h111;
rom[9934] = 12'h111;
rom[9935] = 12'h111;
rom[9936] = 12'h111;
rom[9937] = 12'h111;
rom[9938] = 12'h111;
rom[9939] = 12'h222;
rom[9940] = 12'h111;
rom[9941] = 12'h111;
rom[9942] = 12'h111;
rom[9943] = 12'h111;
rom[9944] = 12'h111;
rom[9945] = 12'h111;
rom[9946] = 12'h111;
rom[9947] = 12'h111;
rom[9948] = 12'h222;
rom[9949] = 12'h222;
rom[9950] = 12'h333;
rom[9951] = 12'h333;
rom[9952] = 12'h444;
rom[9953] = 12'h444;
rom[9954] = 12'h555;
rom[9955] = 12'h555;
rom[9956] = 12'h666;
rom[9957] = 12'h666;
rom[9958] = 12'h555;
rom[9959] = 12'h555;
rom[9960] = 12'h444;
rom[9961] = 12'h444;
rom[9962] = 12'h555;
rom[9963] = 12'h555;
rom[9964] = 12'h444;
rom[9965] = 12'h444;
rom[9966] = 12'h444;
rom[9967] = 12'h333;
rom[9968] = 12'h333;
rom[9969] = 12'h333;
rom[9970] = 12'h444;
rom[9971] = 12'h444;
rom[9972] = 12'h444;
rom[9973] = 12'h444;
rom[9974] = 12'h444;
rom[9975] = 12'h444;
rom[9976] = 12'h444;
rom[9977] = 12'h555;
rom[9978] = 12'h555;
rom[9979] = 12'h666;
rom[9980] = 12'h777;
rom[9981] = 12'h777;
rom[9982] = 12'h777;
rom[9983] = 12'h777;
rom[9984] = 12'h666;
rom[9985] = 12'h666;
rom[9986] = 12'h666;
rom[9987] = 12'h666;
rom[9988] = 12'h666;
rom[9989] = 12'h666;
rom[9990] = 12'h666;
rom[9991] = 12'h777;
rom[9992] = 12'h777;
rom[9993] = 12'h888;
rom[9994] = 12'h888;
rom[9995] = 12'h999;
rom[9996] = 12'haaa;
rom[9997] = 12'haaa;
rom[9998] = 12'haaa;
rom[9999] = 12'haaa;
rom[10000] = 12'h333;
rom[10001] = 12'h333;
rom[10002] = 12'h333;
rom[10003] = 12'h333;
rom[10004] = 12'h333;
rom[10005] = 12'h333;
rom[10006] = 12'h333;
rom[10007] = 12'h222;
rom[10008] = 12'h222;
rom[10009] = 12'h222;
rom[10010] = 12'h222;
rom[10011] = 12'h111;
rom[10012] = 12'h111;
rom[10013] = 12'h111;
rom[10014] = 12'h111;
rom[10015] = 12'h111;
rom[10016] = 12'h111;
rom[10017] = 12'h111;
rom[10018] = 12'h111;
rom[10019] = 12'h111;
rom[10020] = 12'h111;
rom[10021] = 12'h111;
rom[10022] = 12'h  0;
rom[10023] = 12'h  0;
rom[10024] = 12'h111;
rom[10025] = 12'h111;
rom[10026] = 12'h111;
rom[10027] = 12'h111;
rom[10028] = 12'h111;
rom[10029] = 12'h111;
rom[10030] = 12'h111;
rom[10031] = 12'h111;
rom[10032] = 12'h111;
rom[10033] = 12'h111;
rom[10034] = 12'h111;
rom[10035] = 12'h111;
rom[10036] = 12'h111;
rom[10037] = 12'h111;
rom[10038] = 12'h111;
rom[10039] = 12'h111;
rom[10040] = 12'h111;
rom[10041] = 12'h111;
rom[10042] = 12'h111;
rom[10043] = 12'h111;
rom[10044] = 12'h111;
rom[10045] = 12'h111;
rom[10046] = 12'h111;
rom[10047] = 12'h222;
rom[10048] = 12'h222;
rom[10049] = 12'h222;
rom[10050] = 12'h222;
rom[10051] = 12'h333;
rom[10052] = 12'h222;
rom[10053] = 12'h222;
rom[10054] = 12'h222;
rom[10055] = 12'h111;
rom[10056] = 12'h111;
rom[10057] = 12'h222;
rom[10058] = 12'h222;
rom[10059] = 12'h222;
rom[10060] = 12'h333;
rom[10061] = 12'h333;
rom[10062] = 12'h333;
rom[10063] = 12'h333;
rom[10064] = 12'h333;
rom[10065] = 12'h333;
rom[10066] = 12'h333;
rom[10067] = 12'h333;
rom[10068] = 12'h333;
rom[10069] = 12'h222;
rom[10070] = 12'h222;
rom[10071] = 12'h222;
rom[10072] = 12'h222;
rom[10073] = 12'h222;
rom[10074] = 12'h222;
rom[10075] = 12'h222;
rom[10076] = 12'h222;
rom[10077] = 12'h222;
rom[10078] = 12'h222;
rom[10079] = 12'h222;
rom[10080] = 12'h222;
rom[10081] = 12'h222;
rom[10082] = 12'h222;
rom[10083] = 12'h222;
rom[10084] = 12'h222;
rom[10085] = 12'h222;
rom[10086] = 12'h222;
rom[10087] = 12'h222;
rom[10088] = 12'h222;
rom[10089] = 12'h111;
rom[10090] = 12'h111;
rom[10091] = 12'h111;
rom[10092] = 12'h111;
rom[10093] = 12'h111;
rom[10094] = 12'h111;
rom[10095] = 12'h111;
rom[10096] = 12'h111;
rom[10097] = 12'h111;
rom[10098] = 12'h111;
rom[10099] = 12'h111;
rom[10100] = 12'h122;
rom[10101] = 12'h122;
rom[10102] = 12'h222;
rom[10103] = 12'h222;
rom[10104] = 12'h222;
rom[10105] = 12'h222;
rom[10106] = 12'h222;
rom[10107] = 12'h222;
rom[10108] = 12'h211;
rom[10109] = 12'h211;
rom[10110] = 12'h201;
rom[10111] = 12'h200;
rom[10112] = 12'h200;
rom[10113] = 12'h200;
rom[10114] = 12'h310;
rom[10115] = 12'h410;
rom[10116] = 12'h410;
rom[10117] = 12'h620;
rom[10118] = 12'h720;
rom[10119] = 12'h830;
rom[10120] = 12'ha42;
rom[10121] = 12'hb52;
rom[10122] = 12'hb52;
rom[10123] = 12'ha42;
rom[10124] = 12'h820;
rom[10125] = 12'h720;
rom[10126] = 12'h710;
rom[10127] = 12'h610;
rom[10128] = 12'h500;
rom[10129] = 12'h400;
rom[10130] = 12'h400;
rom[10131] = 12'h400;
rom[10132] = 12'h400;
rom[10133] = 12'h400;
rom[10134] = 12'h400;
rom[10135] = 12'h400;
rom[10136] = 12'h400;
rom[10137] = 12'h400;
rom[10138] = 12'h400;
rom[10139] = 12'h400;
rom[10140] = 12'h400;
rom[10141] = 12'h400;
rom[10142] = 12'h500;
rom[10143] = 12'h500;
rom[10144] = 12'h500;
rom[10145] = 12'h500;
rom[10146] = 12'h500;
rom[10147] = 12'h400;
rom[10148] = 12'h400;
rom[10149] = 12'h400;
rom[10150] = 12'h400;
rom[10151] = 12'h300;
rom[10152] = 12'h300;
rom[10153] = 12'h300;
rom[10154] = 12'h300;
rom[10155] = 12'h300;
rom[10156] = 12'h300;
rom[10157] = 12'h300;
rom[10158] = 12'h400;
rom[10159] = 12'h400;
rom[10160] = 12'h300;
rom[10161] = 12'h300;
rom[10162] = 12'h300;
rom[10163] = 12'h300;
rom[10164] = 12'h300;
rom[10165] = 12'h300;
rom[10166] = 12'h300;
rom[10167] = 12'h300;
rom[10168] = 12'h300;
rom[10169] = 12'h300;
rom[10170] = 12'h400;
rom[10171] = 12'h400;
rom[10172] = 12'h410;
rom[10173] = 12'h410;
rom[10174] = 12'h410;
rom[10175] = 12'h410;
rom[10176] = 12'h421;
rom[10177] = 12'h431;
rom[10178] = 12'h543;
rom[10179] = 12'h654;
rom[10180] = 12'h654;
rom[10181] = 12'h765;
rom[10182] = 12'h876;
rom[10183] = 12'h887;
rom[10184] = 12'ha99;
rom[10185] = 12'haaa;
rom[10186] = 12'hbaa;
rom[10187] = 12'hbbb;
rom[10188] = 12'hbbb;
rom[10189] = 12'haab;
rom[10190] = 12'h9aa;
rom[10191] = 12'h899;
rom[10192] = 12'h999;
rom[10193] = 12'h888;
rom[10194] = 12'h888;
rom[10195] = 12'h888;
rom[10196] = 12'h888;
rom[10197] = 12'h888;
rom[10198] = 12'h888;
rom[10199] = 12'h999;
rom[10200] = 12'h999;
rom[10201] = 12'h999;
rom[10202] = 12'h888;
rom[10203] = 12'h999;
rom[10204] = 12'h999;
rom[10205] = 12'h888;
rom[10206] = 12'h666;
rom[10207] = 12'h666;
rom[10208] = 12'h666;
rom[10209] = 12'h666;
rom[10210] = 12'h555;
rom[10211] = 12'h555;
rom[10212] = 12'h444;
rom[10213] = 12'h444;
rom[10214] = 12'h444;
rom[10215] = 12'h444;
rom[10216] = 12'h333;
rom[10217] = 12'h333;
rom[10218] = 12'h222;
rom[10219] = 12'h222;
rom[10220] = 12'h222;
rom[10221] = 12'h222;
rom[10222] = 12'h222;
rom[10223] = 12'h222;
rom[10224] = 12'h111;
rom[10225] = 12'h111;
rom[10226] = 12'h111;
rom[10227] = 12'h111;
rom[10228] = 12'h111;
rom[10229] = 12'h222;
rom[10230] = 12'h222;
rom[10231] = 12'h222;
rom[10232] = 12'h222;
rom[10233] = 12'h222;
rom[10234] = 12'h222;
rom[10235] = 12'h222;
rom[10236] = 12'h333;
rom[10237] = 12'h333;
rom[10238] = 12'h444;
rom[10239] = 12'h444;
rom[10240] = 12'h333;
rom[10241] = 12'h333;
rom[10242] = 12'h444;
rom[10243] = 12'h444;
rom[10244] = 12'h444;
rom[10245] = 12'h555;
rom[10246] = 12'h444;
rom[10247] = 12'h444;
rom[10248] = 12'h444;
rom[10249] = 12'h444;
rom[10250] = 12'h444;
rom[10251] = 12'h444;
rom[10252] = 12'h333;
rom[10253] = 12'h333;
rom[10254] = 12'h333;
rom[10255] = 12'h333;
rom[10256] = 12'h222;
rom[10257] = 12'h222;
rom[10258] = 12'h222;
rom[10259] = 12'h222;
rom[10260] = 12'h222;
rom[10261] = 12'h222;
rom[10262] = 12'h222;
rom[10263] = 12'h222;
rom[10264] = 12'h111;
rom[10265] = 12'h111;
rom[10266] = 12'h111;
rom[10267] = 12'h  0;
rom[10268] = 12'h  0;
rom[10269] = 12'h  0;
rom[10270] = 12'h  0;
rom[10271] = 12'h  0;
rom[10272] = 12'h  0;
rom[10273] = 12'h  0;
rom[10274] = 12'h  0;
rom[10275] = 12'h  0;
rom[10276] = 12'h  0;
rom[10277] = 12'h  0;
rom[10278] = 12'h  0;
rom[10279] = 12'h  0;
rom[10280] = 12'h  0;
rom[10281] = 12'h  0;
rom[10282] = 12'h  0;
rom[10283] = 12'h  0;
rom[10284] = 12'h  0;
rom[10285] = 12'h  0;
rom[10286] = 12'h  0;
rom[10287] = 12'h  0;
rom[10288] = 12'h  0;
rom[10289] = 12'h  0;
rom[10290] = 12'h  0;
rom[10291] = 12'h  0;
rom[10292] = 12'h  0;
rom[10293] = 12'h  0;
rom[10294] = 12'h  0;
rom[10295] = 12'h  0;
rom[10296] = 12'h  0;
rom[10297] = 12'h  0;
rom[10298] = 12'h  0;
rom[10299] = 12'h  0;
rom[10300] = 12'h111;
rom[10301] = 12'h111;
rom[10302] = 12'h  0;
rom[10303] = 12'h  0;
rom[10304] = 12'h  0;
rom[10305] = 12'h  0;
rom[10306] = 12'h  0;
rom[10307] = 12'h  0;
rom[10308] = 12'h  0;
rom[10309] = 12'h  0;
rom[10310] = 12'h  0;
rom[10311] = 12'h  0;
rom[10312] = 12'h  0;
rom[10313] = 12'h  0;
rom[10314] = 12'h111;
rom[10315] = 12'h111;
rom[10316] = 12'h222;
rom[10317] = 12'h333;
rom[10318] = 12'h555;
rom[10319] = 12'h666;
rom[10320] = 12'h777;
rom[10321] = 12'h666;
rom[10322] = 12'h666;
rom[10323] = 12'h444;
rom[10324] = 12'h444;
rom[10325] = 12'h444;
rom[10326] = 12'h444;
rom[10327] = 12'h444;
rom[10328] = 12'h333;
rom[10329] = 12'h222;
rom[10330] = 12'h111;
rom[10331] = 12'h111;
rom[10332] = 12'h111;
rom[10333] = 12'h111;
rom[10334] = 12'h111;
rom[10335] = 12'h111;
rom[10336] = 12'h111;
rom[10337] = 12'h111;
rom[10338] = 12'h111;
rom[10339] = 12'h111;
rom[10340] = 12'h111;
rom[10341] = 12'h111;
rom[10342] = 12'h111;
rom[10343] = 12'h111;
rom[10344] = 12'h111;
rom[10345] = 12'h111;
rom[10346] = 12'h111;
rom[10347] = 12'h111;
rom[10348] = 12'h222;
rom[10349] = 12'h222;
rom[10350] = 12'h222;
rom[10351] = 12'h333;
rom[10352] = 12'h444;
rom[10353] = 12'h444;
rom[10354] = 12'h555;
rom[10355] = 12'h555;
rom[10356] = 12'h666;
rom[10357] = 12'h666;
rom[10358] = 12'h555;
rom[10359] = 12'h555;
rom[10360] = 12'h555;
rom[10361] = 12'h555;
rom[10362] = 12'h444;
rom[10363] = 12'h444;
rom[10364] = 12'h444;
rom[10365] = 12'h444;
rom[10366] = 12'h444;
rom[10367] = 12'h333;
rom[10368] = 12'h333;
rom[10369] = 12'h333;
rom[10370] = 12'h333;
rom[10371] = 12'h333;
rom[10372] = 12'h333;
rom[10373] = 12'h444;
rom[10374] = 12'h444;
rom[10375] = 12'h555;
rom[10376] = 12'h555;
rom[10377] = 12'h666;
rom[10378] = 12'h666;
rom[10379] = 12'h777;
rom[10380] = 12'h777;
rom[10381] = 12'h666;
rom[10382] = 12'h666;
rom[10383] = 12'h666;
rom[10384] = 12'h666;
rom[10385] = 12'h666;
rom[10386] = 12'h666;
rom[10387] = 12'h555;
rom[10388] = 12'h555;
rom[10389] = 12'h666;
rom[10390] = 12'h666;
rom[10391] = 12'h666;
rom[10392] = 12'h777;
rom[10393] = 12'h888;
rom[10394] = 12'h888;
rom[10395] = 12'h999;
rom[10396] = 12'haaa;
rom[10397] = 12'haaa;
rom[10398] = 12'haaa;
rom[10399] = 12'haaa;
rom[10400] = 12'h333;
rom[10401] = 12'h333;
rom[10402] = 12'h222;
rom[10403] = 12'h222;
rom[10404] = 12'h222;
rom[10405] = 12'h222;
rom[10406] = 12'h222;
rom[10407] = 12'h222;
rom[10408] = 12'h222;
rom[10409] = 12'h222;
rom[10410] = 12'h222;
rom[10411] = 12'h111;
rom[10412] = 12'h111;
rom[10413] = 12'h111;
rom[10414] = 12'h111;
rom[10415] = 12'h111;
rom[10416] = 12'h111;
rom[10417] = 12'h111;
rom[10418] = 12'h111;
rom[10419] = 12'h111;
rom[10420] = 12'h111;
rom[10421] = 12'h111;
rom[10422] = 12'h111;
rom[10423] = 12'h111;
rom[10424] = 12'h111;
rom[10425] = 12'h111;
rom[10426] = 12'h111;
rom[10427] = 12'h111;
rom[10428] = 12'h111;
rom[10429] = 12'h111;
rom[10430] = 12'h111;
rom[10431] = 12'h111;
rom[10432] = 12'h111;
rom[10433] = 12'h111;
rom[10434] = 12'h111;
rom[10435] = 12'h111;
rom[10436] = 12'h111;
rom[10437] = 12'h111;
rom[10438] = 12'h111;
rom[10439] = 12'h111;
rom[10440] = 12'h111;
rom[10441] = 12'h111;
rom[10442] = 12'h111;
rom[10443] = 12'h111;
rom[10444] = 12'h111;
rom[10445] = 12'h111;
rom[10446] = 12'h111;
rom[10447] = 12'h111;
rom[10448] = 12'h222;
rom[10449] = 12'h222;
rom[10450] = 12'h333;
rom[10451] = 12'h333;
rom[10452] = 12'h444;
rom[10453] = 12'h333;
rom[10454] = 12'h333;
rom[10455] = 12'h222;
rom[10456] = 12'h222;
rom[10457] = 12'h222;
rom[10458] = 12'h222;
rom[10459] = 12'h222;
rom[10460] = 12'h333;
rom[10461] = 12'h333;
rom[10462] = 12'h444;
rom[10463] = 12'h444;
rom[10464] = 12'h444;
rom[10465] = 12'h444;
rom[10466] = 12'h333;
rom[10467] = 12'h333;
rom[10468] = 12'h333;
rom[10469] = 12'h333;
rom[10470] = 12'h222;
rom[10471] = 12'h222;
rom[10472] = 12'h222;
rom[10473] = 12'h222;
rom[10474] = 12'h222;
rom[10475] = 12'h222;
rom[10476] = 12'h222;
rom[10477] = 12'h222;
rom[10478] = 12'h222;
rom[10479] = 12'h222;
rom[10480] = 12'h222;
rom[10481] = 12'h222;
rom[10482] = 12'h222;
rom[10483] = 12'h222;
rom[10484] = 12'h222;
rom[10485] = 12'h222;
rom[10486] = 12'h222;
rom[10487] = 12'h222;
rom[10488] = 12'h111;
rom[10489] = 12'h111;
rom[10490] = 12'h111;
rom[10491] = 12'h111;
rom[10492] = 12'h111;
rom[10493] = 12'h111;
rom[10494] = 12'h111;
rom[10495] = 12'h111;
rom[10496] = 12'h111;
rom[10497] = 12'h111;
rom[10498] = 12'h111;
rom[10499] = 12'h111;
rom[10500] = 12'h111;
rom[10501] = 12'h121;
rom[10502] = 12'h122;
rom[10503] = 12'h122;
rom[10504] = 12'h111;
rom[10505] = 12'h211;
rom[10506] = 12'h211;
rom[10507] = 12'h211;
rom[10508] = 12'h111;
rom[10509] = 12'h100;
rom[10510] = 12'h100;
rom[10511] = 12'h100;
rom[10512] = 12'h100;
rom[10513] = 12'h200;
rom[10514] = 12'h300;
rom[10515] = 12'h310;
rom[10516] = 12'h410;
rom[10517] = 12'h510;
rom[10518] = 12'h720;
rom[10519] = 12'h820;
rom[10520] = 12'ha41;
rom[10521] = 12'hb52;
rom[10522] = 12'hb52;
rom[10523] = 12'ha41;
rom[10524] = 12'h820;
rom[10525] = 12'h710;
rom[10526] = 12'h710;
rom[10527] = 12'h610;
rom[10528] = 12'h500;
rom[10529] = 12'h400;
rom[10530] = 12'h400;
rom[10531] = 12'h400;
rom[10532] = 12'h400;
rom[10533] = 12'h400;
rom[10534] = 12'h400;
rom[10535] = 12'h400;
rom[10536] = 12'h400;
rom[10537] = 12'h400;
rom[10538] = 12'h400;
rom[10539] = 12'h400;
rom[10540] = 12'h400;
rom[10541] = 12'h400;
rom[10542] = 12'h400;
rom[10543] = 12'h400;
rom[10544] = 12'h400;
rom[10545] = 12'h400;
rom[10546] = 12'h400;
rom[10547] = 12'h400;
rom[10548] = 12'h400;
rom[10549] = 12'h300;
rom[10550] = 12'h300;
rom[10551] = 12'h300;
rom[10552] = 12'h200;
rom[10553] = 12'h200;
rom[10554] = 12'h300;
rom[10555] = 12'h300;
rom[10556] = 12'h300;
rom[10557] = 12'h300;
rom[10558] = 12'h300;
rom[10559] = 12'h300;
rom[10560] = 12'h300;
rom[10561] = 12'h300;
rom[10562] = 12'h300;
rom[10563] = 12'h300;
rom[10564] = 12'h300;
rom[10565] = 12'h300;
rom[10566] = 12'h300;
rom[10567] = 12'h300;
rom[10568] = 12'h300;
rom[10569] = 12'h300;
rom[10570] = 12'h300;
rom[10571] = 12'h300;
rom[10572] = 12'h410;
rom[10573] = 12'h410;
rom[10574] = 12'h410;
rom[10575] = 12'h410;
rom[10576] = 12'h300;
rom[10577] = 12'h310;
rom[10578] = 12'h321;
rom[10579] = 12'h432;
rom[10580] = 12'h543;
rom[10581] = 12'h654;
rom[10582] = 12'h755;
rom[10583] = 12'h765;
rom[10584] = 12'h877;
rom[10585] = 12'h988;
rom[10586] = 12'haaa;
rom[10587] = 12'hbbb;
rom[10588] = 12'hbbb;
rom[10589] = 12'hbbb;
rom[10590] = 12'haaa;
rom[10591] = 12'h999;
rom[10592] = 12'h999;
rom[10593] = 12'h999;
rom[10594] = 12'h888;
rom[10595] = 12'h888;
rom[10596] = 12'h888;
rom[10597] = 12'h888;
rom[10598] = 12'h888;
rom[10599] = 12'h999;
rom[10600] = 12'h999;
rom[10601] = 12'h999;
rom[10602] = 12'h999;
rom[10603] = 12'h999;
rom[10604] = 12'h999;
rom[10605] = 12'h888;
rom[10606] = 12'h777;
rom[10607] = 12'h666;
rom[10608] = 12'h666;
rom[10609] = 12'h666;
rom[10610] = 12'h555;
rom[10611] = 12'h555;
rom[10612] = 12'h555;
rom[10613] = 12'h555;
rom[10614] = 12'h444;
rom[10615] = 12'h444;
rom[10616] = 12'h333;
rom[10617] = 12'h333;
rom[10618] = 12'h333;
rom[10619] = 12'h333;
rom[10620] = 12'h333;
rom[10621] = 12'h333;
rom[10622] = 12'h222;
rom[10623] = 12'h222;
rom[10624] = 12'h222;
rom[10625] = 12'h222;
rom[10626] = 12'h222;
rom[10627] = 12'h222;
rom[10628] = 12'h222;
rom[10629] = 12'h222;
rom[10630] = 12'h222;
rom[10631] = 12'h222;
rom[10632] = 12'h222;
rom[10633] = 12'h222;
rom[10634] = 12'h333;
rom[10635] = 12'h333;
rom[10636] = 12'h333;
rom[10637] = 12'h333;
rom[10638] = 12'h333;
rom[10639] = 12'h444;
rom[10640] = 12'h444;
rom[10641] = 12'h444;
rom[10642] = 12'h555;
rom[10643] = 12'h555;
rom[10644] = 12'h555;
rom[10645] = 12'h444;
rom[10646] = 12'h444;
rom[10647] = 12'h555;
rom[10648] = 12'h444;
rom[10649] = 12'h444;
rom[10650] = 12'h444;
rom[10651] = 12'h444;
rom[10652] = 12'h444;
rom[10653] = 12'h333;
rom[10654] = 12'h333;
rom[10655] = 12'h222;
rom[10656] = 12'h333;
rom[10657] = 12'h222;
rom[10658] = 12'h222;
rom[10659] = 12'h222;
rom[10660] = 12'h222;
rom[10661] = 12'h222;
rom[10662] = 12'h222;
rom[10663] = 12'h222;
rom[10664] = 12'h222;
rom[10665] = 12'h111;
rom[10666] = 12'h111;
rom[10667] = 12'h  0;
rom[10668] = 12'h  0;
rom[10669] = 12'h  0;
rom[10670] = 12'h  0;
rom[10671] = 12'h  0;
rom[10672] = 12'h  0;
rom[10673] = 12'h  0;
rom[10674] = 12'h  0;
rom[10675] = 12'h  0;
rom[10676] = 12'h  0;
rom[10677] = 12'h  0;
rom[10678] = 12'h  0;
rom[10679] = 12'h  0;
rom[10680] = 12'h  0;
rom[10681] = 12'h  0;
rom[10682] = 12'h  0;
rom[10683] = 12'h  0;
rom[10684] = 12'h  0;
rom[10685] = 12'h  0;
rom[10686] = 12'h  0;
rom[10687] = 12'h  0;
rom[10688] = 12'h  0;
rom[10689] = 12'h  0;
rom[10690] = 12'h  0;
rom[10691] = 12'h  0;
rom[10692] = 12'h  0;
rom[10693] = 12'h  0;
rom[10694] = 12'h  0;
rom[10695] = 12'h  0;
rom[10696] = 12'h  0;
rom[10697] = 12'h  0;
rom[10698] = 12'h  0;
rom[10699] = 12'h  0;
rom[10700] = 12'h111;
rom[10701] = 12'h111;
rom[10702] = 12'h  0;
rom[10703] = 12'h  0;
rom[10704] = 12'h  0;
rom[10705] = 12'h  0;
rom[10706] = 12'h  0;
rom[10707] = 12'h  0;
rom[10708] = 12'h  0;
rom[10709] = 12'h  0;
rom[10710] = 12'h  0;
rom[10711] = 12'h  0;
rom[10712] = 12'h  0;
rom[10713] = 12'h  0;
rom[10714] = 12'h111;
rom[10715] = 12'h111;
rom[10716] = 12'h222;
rom[10717] = 12'h444;
rom[10718] = 12'h555;
rom[10719] = 12'h666;
rom[10720] = 12'h777;
rom[10721] = 12'h666;
rom[10722] = 12'h555;
rom[10723] = 12'h444;
rom[10724] = 12'h444;
rom[10725] = 12'h444;
rom[10726] = 12'h444;
rom[10727] = 12'h444;
rom[10728] = 12'h333;
rom[10729] = 12'h222;
rom[10730] = 12'h111;
rom[10731] = 12'h111;
rom[10732] = 12'h111;
rom[10733] = 12'h111;
rom[10734] = 12'h111;
rom[10735] = 12'h111;
rom[10736] = 12'h111;
rom[10737] = 12'h111;
rom[10738] = 12'h111;
rom[10739] = 12'h111;
rom[10740] = 12'h111;
rom[10741] = 12'h111;
rom[10742] = 12'h111;
rom[10743] = 12'h111;
rom[10744] = 12'h111;
rom[10745] = 12'h111;
rom[10746] = 12'h111;
rom[10747] = 12'h111;
rom[10748] = 12'h111;
rom[10749] = 12'h222;
rom[10750] = 12'h222;
rom[10751] = 12'h333;
rom[10752] = 12'h444;
rom[10753] = 12'h444;
rom[10754] = 12'h555;
rom[10755] = 12'h555;
rom[10756] = 12'h666;
rom[10757] = 12'h666;
rom[10758] = 12'h555;
rom[10759] = 12'h555;
rom[10760] = 12'h555;
rom[10761] = 12'h555;
rom[10762] = 12'h444;
rom[10763] = 12'h444;
rom[10764] = 12'h444;
rom[10765] = 12'h444;
rom[10766] = 12'h444;
rom[10767] = 12'h333;
rom[10768] = 12'h333;
rom[10769] = 12'h333;
rom[10770] = 12'h333;
rom[10771] = 12'h444;
rom[10772] = 12'h444;
rom[10773] = 12'h555;
rom[10774] = 12'h555;
rom[10775] = 12'h666;
rom[10776] = 12'h666;
rom[10777] = 12'h666;
rom[10778] = 12'h666;
rom[10779] = 12'h666;
rom[10780] = 12'h666;
rom[10781] = 12'h555;
rom[10782] = 12'h555;
rom[10783] = 12'h555;
rom[10784] = 12'h555;
rom[10785] = 12'h555;
rom[10786] = 12'h555;
rom[10787] = 12'h555;
rom[10788] = 12'h555;
rom[10789] = 12'h666;
rom[10790] = 12'h666;
rom[10791] = 12'h666;
rom[10792] = 12'h777;
rom[10793] = 12'h888;
rom[10794] = 12'h888;
rom[10795] = 12'h999;
rom[10796] = 12'haaa;
rom[10797] = 12'haaa;
rom[10798] = 12'haaa;
rom[10799] = 12'haaa;
rom[10800] = 12'h222;
rom[10801] = 12'h222;
rom[10802] = 12'h222;
rom[10803] = 12'h222;
rom[10804] = 12'h222;
rom[10805] = 12'h222;
rom[10806] = 12'h222;
rom[10807] = 12'h222;
rom[10808] = 12'h222;
rom[10809] = 12'h222;
rom[10810] = 12'h222;
rom[10811] = 12'h111;
rom[10812] = 12'h111;
rom[10813] = 12'h111;
rom[10814] = 12'h111;
rom[10815] = 12'h111;
rom[10816] = 12'h111;
rom[10817] = 12'h111;
rom[10818] = 12'h111;
rom[10819] = 12'h111;
rom[10820] = 12'h111;
rom[10821] = 12'h111;
rom[10822] = 12'h111;
rom[10823] = 12'h111;
rom[10824] = 12'h111;
rom[10825] = 12'h111;
rom[10826] = 12'h111;
rom[10827] = 12'h111;
rom[10828] = 12'h111;
rom[10829] = 12'h111;
rom[10830] = 12'h111;
rom[10831] = 12'h111;
rom[10832] = 12'h111;
rom[10833] = 12'h111;
rom[10834] = 12'h111;
rom[10835] = 12'h111;
rom[10836] = 12'h111;
rom[10837] = 12'h111;
rom[10838] = 12'h111;
rom[10839] = 12'h111;
rom[10840] = 12'h111;
rom[10841] = 12'h111;
rom[10842] = 12'h111;
rom[10843] = 12'h111;
rom[10844] = 12'h111;
rom[10845] = 12'h111;
rom[10846] = 12'h111;
rom[10847] = 12'h111;
rom[10848] = 12'h111;
rom[10849] = 12'h222;
rom[10850] = 12'h222;
rom[10851] = 12'h333;
rom[10852] = 12'h333;
rom[10853] = 12'h444;
rom[10854] = 12'h444;
rom[10855] = 12'h444;
rom[10856] = 12'h444;
rom[10857] = 12'h333;
rom[10858] = 12'h333;
rom[10859] = 12'h333;
rom[10860] = 12'h333;
rom[10861] = 12'h333;
rom[10862] = 12'h444;
rom[10863] = 12'h444;
rom[10864] = 12'h555;
rom[10865] = 12'h444;
rom[10866] = 12'h444;
rom[10867] = 12'h444;
rom[10868] = 12'h444;
rom[10869] = 12'h444;
rom[10870] = 12'h333;
rom[10871] = 12'h333;
rom[10872] = 12'h222;
rom[10873] = 12'h222;
rom[10874] = 12'h222;
rom[10875] = 12'h222;
rom[10876] = 12'h222;
rom[10877] = 12'h222;
rom[10878] = 12'h222;
rom[10879] = 12'h222;
rom[10880] = 12'h222;
rom[10881] = 12'h222;
rom[10882] = 12'h222;
rom[10883] = 12'h222;
rom[10884] = 12'h222;
rom[10885] = 12'h222;
rom[10886] = 12'h222;
rom[10887] = 12'h111;
rom[10888] = 12'h111;
rom[10889] = 12'h111;
rom[10890] = 12'h111;
rom[10891] = 12'h111;
rom[10892] = 12'h111;
rom[10893] = 12'h111;
rom[10894] = 12'h111;
rom[10895] = 12'h111;
rom[10896] = 12'h111;
rom[10897] = 12'h111;
rom[10898] = 12'h111;
rom[10899] = 12'h111;
rom[10900] = 12'h111;
rom[10901] = 12'h111;
rom[10902] = 12'h111;
rom[10903] = 12'h121;
rom[10904] = 12'h111;
rom[10905] = 12'h111;
rom[10906] = 12'h111;
rom[10907] = 12'h111;
rom[10908] = 12'h100;
rom[10909] = 12'h100;
rom[10910] = 12'h100;
rom[10911] = 12'h100;
rom[10912] = 12'h100;
rom[10913] = 12'h200;
rom[10914] = 12'h200;
rom[10915] = 12'h300;
rom[10916] = 12'h410;
rom[10917] = 12'h510;
rom[10918] = 12'h620;
rom[10919] = 12'h720;
rom[10920] = 12'h941;
rom[10921] = 12'ha42;
rom[10922] = 12'hb42;
rom[10923] = 12'ha41;
rom[10924] = 12'h820;
rom[10925] = 12'h710;
rom[10926] = 12'h710;
rom[10927] = 12'h610;
rom[10928] = 12'h500;
rom[10929] = 12'h400;
rom[10930] = 12'h400;
rom[10931] = 12'h400;
rom[10932] = 12'h400;
rom[10933] = 12'h400;
rom[10934] = 12'h400;
rom[10935] = 12'h400;
rom[10936] = 12'h400;
rom[10937] = 12'h400;
rom[10938] = 12'h400;
rom[10939] = 12'h400;
rom[10940] = 12'h400;
rom[10941] = 12'h400;
rom[10942] = 12'h400;
rom[10943] = 12'h400;
rom[10944] = 12'h400;
rom[10945] = 12'h400;
rom[10946] = 12'h400;
rom[10947] = 12'h300;
rom[10948] = 12'h300;
rom[10949] = 12'h300;
rom[10950] = 12'h300;
rom[10951] = 12'h200;
rom[10952] = 12'h200;
rom[10953] = 12'h200;
rom[10954] = 12'h200;
rom[10955] = 12'h200;
rom[10956] = 12'h200;
rom[10957] = 12'h200;
rom[10958] = 12'h200;
rom[10959] = 12'h300;
rom[10960] = 12'h300;
rom[10961] = 12'h200;
rom[10962] = 12'h300;
rom[10963] = 12'h300;
rom[10964] = 12'h300;
rom[10965] = 12'h300;
rom[10966] = 12'h300;
rom[10967] = 12'h300;
rom[10968] = 12'h300;
rom[10969] = 12'h300;
rom[10970] = 12'h300;
rom[10971] = 12'h300;
rom[10972] = 12'h300;
rom[10973] = 12'h400;
rom[10974] = 12'h410;
rom[10975] = 12'h310;
rom[10976] = 12'h300;
rom[10977] = 12'h300;
rom[10978] = 12'h310;
rom[10979] = 12'h411;
rom[10980] = 12'h421;
rom[10981] = 12'h532;
rom[10982] = 12'h644;
rom[10983] = 12'h654;
rom[10984] = 12'h655;
rom[10985] = 12'h766;
rom[10986] = 12'h988;
rom[10987] = 12'ha99;
rom[10988] = 12'hbaa;
rom[10989] = 12'hbbb;
rom[10990] = 12'hbbb;
rom[10991] = 12'haaa;
rom[10992] = 12'haaa;
rom[10993] = 12'h999;
rom[10994] = 12'h888;
rom[10995] = 12'h888;
rom[10996] = 12'h888;
rom[10997] = 12'h888;
rom[10998] = 12'h888;
rom[10999] = 12'h999;
rom[11000] = 12'h999;
rom[11001] = 12'h999;
rom[11002] = 12'h999;
rom[11003] = 12'h999;
rom[11004] = 12'h999;
rom[11005] = 12'h888;
rom[11006] = 12'h777;
rom[11007] = 12'h666;
rom[11008] = 12'h666;
rom[11009] = 12'h666;
rom[11010] = 12'h666;
rom[11011] = 12'h666;
rom[11012] = 12'h666;
rom[11013] = 12'h555;
rom[11014] = 12'h444;
rom[11015] = 12'h444;
rom[11016] = 12'h444;
rom[11017] = 12'h444;
rom[11018] = 12'h333;
rom[11019] = 12'h333;
rom[11020] = 12'h333;
rom[11021] = 12'h333;
rom[11022] = 12'h333;
rom[11023] = 12'h222;
rom[11024] = 12'h333;
rom[11025] = 12'h333;
rom[11026] = 12'h222;
rom[11027] = 12'h222;
rom[11028] = 12'h333;
rom[11029] = 12'h333;
rom[11030] = 12'h333;
rom[11031] = 12'h333;
rom[11032] = 12'h333;
rom[11033] = 12'h333;
rom[11034] = 12'h333;
rom[11035] = 12'h333;
rom[11036] = 12'h333;
rom[11037] = 12'h333;
rom[11038] = 12'h444;
rom[11039] = 12'h444;
rom[11040] = 12'h555;
rom[11041] = 12'h666;
rom[11042] = 12'h666;
rom[11043] = 12'h666;
rom[11044] = 12'h555;
rom[11045] = 12'h555;
rom[11046] = 12'h444;
rom[11047] = 12'h555;
rom[11048] = 12'h444;
rom[11049] = 12'h444;
rom[11050] = 12'h444;
rom[11051] = 12'h444;
rom[11052] = 12'h333;
rom[11053] = 12'h333;
rom[11054] = 12'h222;
rom[11055] = 12'h222;
rom[11056] = 12'h222;
rom[11057] = 12'h222;
rom[11058] = 12'h222;
rom[11059] = 12'h222;
rom[11060] = 12'h222;
rom[11061] = 12'h222;
rom[11062] = 12'h222;
rom[11063] = 12'h222;
rom[11064] = 12'h111;
rom[11065] = 12'h111;
rom[11066] = 12'h111;
rom[11067] = 12'h111;
rom[11068] = 12'h  0;
rom[11069] = 12'h  0;
rom[11070] = 12'h  0;
rom[11071] = 12'h  0;
rom[11072] = 12'h  0;
rom[11073] = 12'h  0;
rom[11074] = 12'h  0;
rom[11075] = 12'h  0;
rom[11076] = 12'h  0;
rom[11077] = 12'h  0;
rom[11078] = 12'h  0;
rom[11079] = 12'h  0;
rom[11080] = 12'h  0;
rom[11081] = 12'h  0;
rom[11082] = 12'h  0;
rom[11083] = 12'h  0;
rom[11084] = 12'h  0;
rom[11085] = 12'h  0;
rom[11086] = 12'h  0;
rom[11087] = 12'h  0;
rom[11088] = 12'h  0;
rom[11089] = 12'h  0;
rom[11090] = 12'h  0;
rom[11091] = 12'h  0;
rom[11092] = 12'h  0;
rom[11093] = 12'h  0;
rom[11094] = 12'h  0;
rom[11095] = 12'h  0;
rom[11096] = 12'h  0;
rom[11097] = 12'h  0;
rom[11098] = 12'h  0;
rom[11099] = 12'h  0;
rom[11100] = 12'h111;
rom[11101] = 12'h111;
rom[11102] = 12'h  0;
rom[11103] = 12'h  0;
rom[11104] = 12'h  0;
rom[11105] = 12'h  0;
rom[11106] = 12'h  0;
rom[11107] = 12'h  0;
rom[11108] = 12'h  0;
rom[11109] = 12'h  0;
rom[11110] = 12'h  0;
rom[11111] = 12'h  0;
rom[11112] = 12'h  0;
rom[11113] = 12'h111;
rom[11114] = 12'h111;
rom[11115] = 12'h111;
rom[11116] = 12'h222;
rom[11117] = 12'h444;
rom[11118] = 12'h666;
rom[11119] = 12'h777;
rom[11120] = 12'h777;
rom[11121] = 12'h666;
rom[11122] = 12'h444;
rom[11123] = 12'h444;
rom[11124] = 12'h444;
rom[11125] = 12'h444;
rom[11126] = 12'h444;
rom[11127] = 12'h444;
rom[11128] = 12'h333;
rom[11129] = 12'h222;
rom[11130] = 12'h111;
rom[11131] = 12'h111;
rom[11132] = 12'h111;
rom[11133] = 12'h111;
rom[11134] = 12'h111;
rom[11135] = 12'h111;
rom[11136] = 12'h111;
rom[11137] = 12'h111;
rom[11138] = 12'h111;
rom[11139] = 12'h111;
rom[11140] = 12'h111;
rom[11141] = 12'h111;
rom[11142] = 12'h111;
rom[11143] = 12'h111;
rom[11144] = 12'h  0;
rom[11145] = 12'h111;
rom[11146] = 12'h111;
rom[11147] = 12'h111;
rom[11148] = 12'h111;
rom[11149] = 12'h222;
rom[11150] = 12'h222;
rom[11151] = 12'h333;
rom[11152] = 12'h444;
rom[11153] = 12'h444;
rom[11154] = 12'h555;
rom[11155] = 12'h555;
rom[11156] = 12'h666;
rom[11157] = 12'h666;
rom[11158] = 12'h555;
rom[11159] = 12'h555;
rom[11160] = 12'h555;
rom[11161] = 12'h555;
rom[11162] = 12'h444;
rom[11163] = 12'h444;
rom[11164] = 12'h444;
rom[11165] = 12'h333;
rom[11166] = 12'h333;
rom[11167] = 12'h333;
rom[11168] = 12'h444;
rom[11169] = 12'h444;
rom[11170] = 12'h444;
rom[11171] = 12'h555;
rom[11172] = 12'h555;
rom[11173] = 12'h666;
rom[11174] = 12'h666;
rom[11175] = 12'h666;
rom[11176] = 12'h666;
rom[11177] = 12'h666;
rom[11178] = 12'h555;
rom[11179] = 12'h555;
rom[11180] = 12'h444;
rom[11181] = 12'h444;
rom[11182] = 12'h555;
rom[11183] = 12'h555;
rom[11184] = 12'h444;
rom[11185] = 12'h555;
rom[11186] = 12'h555;
rom[11187] = 12'h555;
rom[11188] = 12'h555;
rom[11189] = 12'h666;
rom[11190] = 12'h666;
rom[11191] = 12'h666;
rom[11192] = 12'h777;
rom[11193] = 12'h888;
rom[11194] = 12'h888;
rom[11195] = 12'h999;
rom[11196] = 12'haaa;
rom[11197] = 12'haaa;
rom[11198] = 12'haaa;
rom[11199] = 12'haaa;
rom[11200] = 12'h222;
rom[11201] = 12'h222;
rom[11202] = 12'h222;
rom[11203] = 12'h222;
rom[11204] = 12'h222;
rom[11205] = 12'h222;
rom[11206] = 12'h111;
rom[11207] = 12'h111;
rom[11208] = 12'h222;
rom[11209] = 12'h222;
rom[11210] = 12'h111;
rom[11211] = 12'h111;
rom[11212] = 12'h111;
rom[11213] = 12'h111;
rom[11214] = 12'h111;
rom[11215] = 12'h111;
rom[11216] = 12'h111;
rom[11217] = 12'h111;
rom[11218] = 12'h111;
rom[11219] = 12'h111;
rom[11220] = 12'h111;
rom[11221] = 12'h111;
rom[11222] = 12'h111;
rom[11223] = 12'h111;
rom[11224] = 12'h111;
rom[11225] = 12'h111;
rom[11226] = 12'h111;
rom[11227] = 12'h111;
rom[11228] = 12'h111;
rom[11229] = 12'h111;
rom[11230] = 12'h111;
rom[11231] = 12'h111;
rom[11232] = 12'h111;
rom[11233] = 12'h111;
rom[11234] = 12'h111;
rom[11235] = 12'h111;
rom[11236] = 12'h111;
rom[11237] = 12'h111;
rom[11238] = 12'h111;
rom[11239] = 12'h111;
rom[11240] = 12'h111;
rom[11241] = 12'h111;
rom[11242] = 12'h111;
rom[11243] = 12'h111;
rom[11244] = 12'h111;
rom[11245] = 12'h111;
rom[11246] = 12'h111;
rom[11247] = 12'h111;
rom[11248] = 12'h111;
rom[11249] = 12'h111;
rom[11250] = 12'h111;
rom[11251] = 12'h222;
rom[11252] = 12'h222;
rom[11253] = 12'h333;
rom[11254] = 12'h444;
rom[11255] = 12'h444;
rom[11256] = 12'h444;
rom[11257] = 12'h444;
rom[11258] = 12'h444;
rom[11259] = 12'h444;
rom[11260] = 12'h444;
rom[11261] = 12'h444;
rom[11262] = 12'h444;
rom[11263] = 12'h444;
rom[11264] = 12'h555;
rom[11265] = 12'h555;
rom[11266] = 12'h555;
rom[11267] = 12'h555;
rom[11268] = 12'h555;
rom[11269] = 12'h555;
rom[11270] = 12'h444;
rom[11271] = 12'h444;
rom[11272] = 12'h333;
rom[11273] = 12'h333;
rom[11274] = 12'h333;
rom[11275] = 12'h333;
rom[11276] = 12'h333;
rom[11277] = 12'h333;
rom[11278] = 12'h333;
rom[11279] = 12'h222;
rom[11280] = 12'h333;
rom[11281] = 12'h333;
rom[11282] = 12'h333;
rom[11283] = 12'h222;
rom[11284] = 12'h222;
rom[11285] = 12'h222;
rom[11286] = 12'h222;
rom[11287] = 12'h111;
rom[11288] = 12'h111;
rom[11289] = 12'h111;
rom[11290] = 12'h111;
rom[11291] = 12'h111;
rom[11292] = 12'h111;
rom[11293] = 12'h111;
rom[11294] = 12'h111;
rom[11295] = 12'h111;
rom[11296] = 12'h111;
rom[11297] = 12'h111;
rom[11298] = 12'h111;
rom[11299] = 12'h111;
rom[11300] = 12'h111;
rom[11301] = 12'h111;
rom[11302] = 12'h111;
rom[11303] = 12'h111;
rom[11304] = 12'h111;
rom[11305] = 12'h111;
rom[11306] = 12'h111;
rom[11307] = 12'h100;
rom[11308] = 12'h100;
rom[11309] = 12'h100;
rom[11310] = 12'h100;
rom[11311] = 12'h100;
rom[11312] = 12'h100;
rom[11313] = 12'h200;
rom[11314] = 12'h200;
rom[11315] = 12'h300;
rom[11316] = 12'h400;
rom[11317] = 12'h510;
rom[11318] = 12'h610;
rom[11319] = 12'h720;
rom[11320] = 12'h931;
rom[11321] = 12'ha41;
rom[11322] = 12'ha42;
rom[11323] = 12'ha31;
rom[11324] = 12'h820;
rom[11325] = 12'h710;
rom[11326] = 12'h710;
rom[11327] = 12'h600;
rom[11328] = 12'h500;
rom[11329] = 12'h400;
rom[11330] = 12'h400;
rom[11331] = 12'h400;
rom[11332] = 12'h400;
rom[11333] = 12'h400;
rom[11334] = 12'h400;
rom[11335] = 12'h400;
rom[11336] = 12'h400;
rom[11337] = 12'h400;
rom[11338] = 12'h400;
rom[11339] = 12'h400;
rom[11340] = 12'h400;
rom[11341] = 12'h400;
rom[11342] = 12'h400;
rom[11343] = 12'h400;
rom[11344] = 12'h400;
rom[11345] = 12'h400;
rom[11346] = 12'h300;
rom[11347] = 12'h300;
rom[11348] = 12'h300;
rom[11349] = 12'h200;
rom[11350] = 12'h200;
rom[11351] = 12'h200;
rom[11352] = 12'h200;
rom[11353] = 12'h200;
rom[11354] = 12'h200;
rom[11355] = 12'h200;
rom[11356] = 12'h200;
rom[11357] = 12'h200;
rom[11358] = 12'h200;
rom[11359] = 12'h200;
rom[11360] = 12'h200;
rom[11361] = 12'h200;
rom[11362] = 12'h200;
rom[11363] = 12'h200;
rom[11364] = 12'h200;
rom[11365] = 12'h200;
rom[11366] = 12'h200;
rom[11367] = 12'h200;
rom[11368] = 12'h200;
rom[11369] = 12'h300;
rom[11370] = 12'h300;
rom[11371] = 12'h300;
rom[11372] = 12'h300;
rom[11373] = 12'h300;
rom[11374] = 12'h300;
rom[11375] = 12'h300;
rom[11376] = 12'h300;
rom[11377] = 12'h310;
rom[11378] = 12'h410;
rom[11379] = 12'h310;
rom[11380] = 12'h310;
rom[11381] = 12'h421;
rom[11382] = 12'h533;
rom[11383] = 12'h544;
rom[11384] = 12'h654;
rom[11385] = 12'h655;
rom[11386] = 12'h766;
rom[11387] = 12'h877;
rom[11388] = 12'h999;
rom[11389] = 12'haba;
rom[11390] = 12'hbbb;
rom[11391] = 12'hbbb;
rom[11392] = 12'haaa;
rom[11393] = 12'h999;
rom[11394] = 12'h999;
rom[11395] = 12'h888;
rom[11396] = 12'h888;
rom[11397] = 12'h888;
rom[11398] = 12'h888;
rom[11399] = 12'h999;
rom[11400] = 12'h999;
rom[11401] = 12'h999;
rom[11402] = 12'h999;
rom[11403] = 12'h999;
rom[11404] = 12'h999;
rom[11405] = 12'h999;
rom[11406] = 12'h777;
rom[11407] = 12'h777;
rom[11408] = 12'h666;
rom[11409] = 12'h666;
rom[11410] = 12'h666;
rom[11411] = 12'h666;
rom[11412] = 12'h666;
rom[11413] = 12'h555;
rom[11414] = 12'h444;
rom[11415] = 12'h444;
rom[11416] = 12'h444;
rom[11417] = 12'h444;
rom[11418] = 12'h444;
rom[11419] = 12'h444;
rom[11420] = 12'h444;
rom[11421] = 12'h444;
rom[11422] = 12'h333;
rom[11423] = 12'h333;
rom[11424] = 12'h333;
rom[11425] = 12'h333;
rom[11426] = 12'h333;
rom[11427] = 12'h333;
rom[11428] = 12'h333;
rom[11429] = 12'h333;
rom[11430] = 12'h333;
rom[11431] = 12'h444;
rom[11432] = 12'h333;
rom[11433] = 12'h333;
rom[11434] = 12'h333;
rom[11435] = 12'h333;
rom[11436] = 12'h444;
rom[11437] = 12'h444;
rom[11438] = 12'h555;
rom[11439] = 12'h555;
rom[11440] = 12'h666;
rom[11441] = 12'h666;
rom[11442] = 12'h666;
rom[11443] = 12'h666;
rom[11444] = 12'h666;
rom[11445] = 12'h555;
rom[11446] = 12'h555;
rom[11447] = 12'h444;
rom[11448] = 12'h444;
rom[11449] = 12'h444;
rom[11450] = 12'h333;
rom[11451] = 12'h333;
rom[11452] = 12'h333;
rom[11453] = 12'h333;
rom[11454] = 12'h222;
rom[11455] = 12'h222;
rom[11456] = 12'h222;
rom[11457] = 12'h222;
rom[11458] = 12'h222;
rom[11459] = 12'h333;
rom[11460] = 12'h333;
rom[11461] = 12'h333;
rom[11462] = 12'h222;
rom[11463] = 12'h222;
rom[11464] = 12'h111;
rom[11465] = 12'h111;
rom[11466] = 12'h111;
rom[11467] = 12'h111;
rom[11468] = 12'h  0;
rom[11469] = 12'h  0;
rom[11470] = 12'h  0;
rom[11471] = 12'h  0;
rom[11472] = 12'h  0;
rom[11473] = 12'h  0;
rom[11474] = 12'h  0;
rom[11475] = 12'h  0;
rom[11476] = 12'h  0;
rom[11477] = 12'h  0;
rom[11478] = 12'h  0;
rom[11479] = 12'h  0;
rom[11480] = 12'h  0;
rom[11481] = 12'h  0;
rom[11482] = 12'h  0;
rom[11483] = 12'h  0;
rom[11484] = 12'h  0;
rom[11485] = 12'h  0;
rom[11486] = 12'h  0;
rom[11487] = 12'h  0;
rom[11488] = 12'h  0;
rom[11489] = 12'h  0;
rom[11490] = 12'h  0;
rom[11491] = 12'h  0;
rom[11492] = 12'h  0;
rom[11493] = 12'h  0;
rom[11494] = 12'h  0;
rom[11495] = 12'h  0;
rom[11496] = 12'h  0;
rom[11497] = 12'h  0;
rom[11498] = 12'h  0;
rom[11499] = 12'h  0;
rom[11500] = 12'h111;
rom[11501] = 12'h111;
rom[11502] = 12'h  0;
rom[11503] = 12'h  0;
rom[11504] = 12'h  0;
rom[11505] = 12'h  0;
rom[11506] = 12'h  0;
rom[11507] = 12'h  0;
rom[11508] = 12'h  0;
rom[11509] = 12'h  0;
rom[11510] = 12'h  0;
rom[11511] = 12'h  0;
rom[11512] = 12'h111;
rom[11513] = 12'h111;
rom[11514] = 12'h111;
rom[11515] = 12'h111;
rom[11516] = 12'h333;
rom[11517] = 12'h555;
rom[11518] = 12'h666;
rom[11519] = 12'h666;
rom[11520] = 12'h666;
rom[11521] = 12'h555;
rom[11522] = 12'h444;
rom[11523] = 12'h333;
rom[11524] = 12'h444;
rom[11525] = 12'h555;
rom[11526] = 12'h444;
rom[11527] = 12'h444;
rom[11528] = 12'h333;
rom[11529] = 12'h222;
rom[11530] = 12'h111;
rom[11531] = 12'h111;
rom[11532] = 12'h111;
rom[11533] = 12'h111;
rom[11534] = 12'h111;
rom[11535] = 12'h111;
rom[11536] = 12'h111;
rom[11537] = 12'h111;
rom[11538] = 12'h111;
rom[11539] = 12'h  0;
rom[11540] = 12'h  0;
rom[11541] = 12'h  0;
rom[11542] = 12'h  0;
rom[11543] = 12'h  0;
rom[11544] = 12'h  0;
rom[11545] = 12'h111;
rom[11546] = 12'h111;
rom[11547] = 12'h111;
rom[11548] = 12'h111;
rom[11549] = 12'h222;
rom[11550] = 12'h222;
rom[11551] = 12'h333;
rom[11552] = 12'h444;
rom[11553] = 12'h444;
rom[11554] = 12'h555;
rom[11555] = 12'h666;
rom[11556] = 12'h666;
rom[11557] = 12'h666;
rom[11558] = 12'h555;
rom[11559] = 12'h555;
rom[11560] = 12'h555;
rom[11561] = 12'h555;
rom[11562] = 12'h444;
rom[11563] = 12'h444;
rom[11564] = 12'h444;
rom[11565] = 12'h333;
rom[11566] = 12'h333;
rom[11567] = 12'h444;
rom[11568] = 12'h444;
rom[11569] = 12'h555;
rom[11570] = 12'h555;
rom[11571] = 12'h666;
rom[11572] = 12'h666;
rom[11573] = 12'h666;
rom[11574] = 12'h666;
rom[11575] = 12'h666;
rom[11576] = 12'h555;
rom[11577] = 12'h444;
rom[11578] = 12'h444;
rom[11579] = 12'h444;
rom[11580] = 12'h444;
rom[11581] = 12'h444;
rom[11582] = 12'h444;
rom[11583] = 12'h444;
rom[11584] = 12'h444;
rom[11585] = 12'h444;
rom[11586] = 12'h555;
rom[11587] = 12'h555;
rom[11588] = 12'h555;
rom[11589] = 12'h666;
rom[11590] = 12'h666;
rom[11591] = 12'h777;
rom[11592] = 12'h777;
rom[11593] = 12'h888;
rom[11594] = 12'h888;
rom[11595] = 12'h999;
rom[11596] = 12'haaa;
rom[11597] = 12'haaa;
rom[11598] = 12'haaa;
rom[11599] = 12'haaa;
rom[11600] = 12'h333;
rom[11601] = 12'h222;
rom[11602] = 12'h222;
rom[11603] = 12'h222;
rom[11604] = 12'h222;
rom[11605] = 12'h222;
rom[11606] = 12'h222;
rom[11607] = 12'h111;
rom[11608] = 12'h111;
rom[11609] = 12'h111;
rom[11610] = 12'h111;
rom[11611] = 12'h111;
rom[11612] = 12'h111;
rom[11613] = 12'h111;
rom[11614] = 12'h111;
rom[11615] = 12'h111;
rom[11616] = 12'h111;
rom[11617] = 12'h111;
rom[11618] = 12'h111;
rom[11619] = 12'h111;
rom[11620] = 12'h111;
rom[11621] = 12'h111;
rom[11622] = 12'h111;
rom[11623] = 12'h111;
rom[11624] = 12'h111;
rom[11625] = 12'h111;
rom[11626] = 12'h111;
rom[11627] = 12'h111;
rom[11628] = 12'h111;
rom[11629] = 12'h111;
rom[11630] = 12'h111;
rom[11631] = 12'h111;
rom[11632] = 12'h111;
rom[11633] = 12'h111;
rom[11634] = 12'h111;
rom[11635] = 12'h111;
rom[11636] = 12'h111;
rom[11637] = 12'h222;
rom[11638] = 12'h222;
rom[11639] = 12'h222;
rom[11640] = 12'h111;
rom[11641] = 12'h111;
rom[11642] = 12'h111;
rom[11643] = 12'h111;
rom[11644] = 12'h111;
rom[11645] = 12'h111;
rom[11646] = 12'h111;
rom[11647] = 12'h111;
rom[11648] = 12'h111;
rom[11649] = 12'h111;
rom[11650] = 12'h111;
rom[11651] = 12'h222;
rom[11652] = 12'h222;
rom[11653] = 12'h222;
rom[11654] = 12'h333;
rom[11655] = 12'h333;
rom[11656] = 12'h444;
rom[11657] = 12'h444;
rom[11658] = 12'h444;
rom[11659] = 12'h444;
rom[11660] = 12'h444;
rom[11661] = 12'h444;
rom[11662] = 12'h444;
rom[11663] = 12'h444;
rom[11664] = 12'h444;
rom[11665] = 12'h555;
rom[11666] = 12'h555;
rom[11667] = 12'h666;
rom[11668] = 12'h666;
rom[11669] = 12'h666;
rom[11670] = 12'h555;
rom[11671] = 12'h555;
rom[11672] = 12'h444;
rom[11673] = 12'h444;
rom[11674] = 12'h444;
rom[11675] = 12'h333;
rom[11676] = 12'h333;
rom[11677] = 12'h333;
rom[11678] = 12'h333;
rom[11679] = 12'h333;
rom[11680] = 12'h333;
rom[11681] = 12'h333;
rom[11682] = 12'h333;
rom[11683] = 12'h222;
rom[11684] = 12'h222;
rom[11685] = 12'h222;
rom[11686] = 12'h222;
rom[11687] = 12'h111;
rom[11688] = 12'h111;
rom[11689] = 12'h111;
rom[11690] = 12'h111;
rom[11691] = 12'h111;
rom[11692] = 12'h111;
rom[11693] = 12'h111;
rom[11694] = 12'h111;
rom[11695] = 12'h111;
rom[11696] = 12'h111;
rom[11697] = 12'h111;
rom[11698] = 12'h111;
rom[11699] = 12'h111;
rom[11700] = 12'h111;
rom[11701] = 12'h111;
rom[11702] = 12'h111;
rom[11703] = 12'h111;
rom[11704] = 12'h111;
rom[11705] = 12'h111;
rom[11706] = 12'h100;
rom[11707] = 12'h100;
rom[11708] = 12'h  0;
rom[11709] = 12'h  0;
rom[11710] = 12'h100;
rom[11711] = 12'h100;
rom[11712] = 12'h100;
rom[11713] = 12'h100;
rom[11714] = 12'h200;
rom[11715] = 12'h300;
rom[11716] = 12'h400;
rom[11717] = 12'h510;
rom[11718] = 12'h610;
rom[11719] = 12'h720;
rom[11720] = 12'h930;
rom[11721] = 12'ha31;
rom[11722] = 12'ha42;
rom[11723] = 12'ha31;
rom[11724] = 12'h921;
rom[11725] = 12'h820;
rom[11726] = 12'h710;
rom[11727] = 12'h600;
rom[11728] = 12'h500;
rom[11729] = 12'h500;
rom[11730] = 12'h500;
rom[11731] = 12'h500;
rom[11732] = 12'h400;
rom[11733] = 12'h400;
rom[11734] = 12'h400;
rom[11735] = 12'h400;
rom[11736] = 12'h400;
rom[11737] = 12'h400;
rom[11738] = 12'h400;
rom[11739] = 12'h400;
rom[11740] = 12'h400;
rom[11741] = 12'h400;
rom[11742] = 12'h400;
rom[11743] = 12'h400;
rom[11744] = 12'h400;
rom[11745] = 12'h300;
rom[11746] = 12'h300;
rom[11747] = 12'h300;
rom[11748] = 12'h200;
rom[11749] = 12'h200;
rom[11750] = 12'h200;
rom[11751] = 12'h100;
rom[11752] = 12'h100;
rom[11753] = 12'h100;
rom[11754] = 12'h100;
rom[11755] = 12'h200;
rom[11756] = 12'h200;
rom[11757] = 12'h200;
rom[11758] = 12'h200;
rom[11759] = 12'h200;
rom[11760] = 12'h200;
rom[11761] = 12'h200;
rom[11762] = 12'h200;
rom[11763] = 12'h200;
rom[11764] = 12'h200;
rom[11765] = 12'h200;
rom[11766] = 12'h200;
rom[11767] = 12'h200;
rom[11768] = 12'h200;
rom[11769] = 12'h200;
rom[11770] = 12'h200;
rom[11771] = 12'h300;
rom[11772] = 12'h300;
rom[11773] = 12'h300;
rom[11774] = 12'h300;
rom[11775] = 12'h300;
rom[11776] = 12'h400;
rom[11777] = 12'h410;
rom[11778] = 12'h410;
rom[11779] = 12'h310;
rom[11780] = 12'h310;
rom[11781] = 12'h310;
rom[11782] = 12'h421;
rom[11783] = 12'h532;
rom[11784] = 12'h644;
rom[11785] = 12'h544;
rom[11786] = 12'h655;
rom[11787] = 12'h665;
rom[11788] = 12'h777;
rom[11789] = 12'h999;
rom[11790] = 12'haaa;
rom[11791] = 12'hbbb;
rom[11792] = 12'hbbb;
rom[11793] = 12'haaa;
rom[11794] = 12'haaa;
rom[11795] = 12'haaa;
rom[11796] = 12'h999;
rom[11797] = 12'h999;
rom[11798] = 12'h999;
rom[11799] = 12'h999;
rom[11800] = 12'h999;
rom[11801] = 12'haaa;
rom[11802] = 12'h999;
rom[11803] = 12'h999;
rom[11804] = 12'h999;
rom[11805] = 12'h999;
rom[11806] = 12'h888;
rom[11807] = 12'h777;
rom[11808] = 12'h777;
rom[11809] = 12'h666;
rom[11810] = 12'h666;
rom[11811] = 12'h777;
rom[11812] = 12'h666;
rom[11813] = 12'h666;
rom[11814] = 12'h555;
rom[11815] = 12'h555;
rom[11816] = 12'h555;
rom[11817] = 12'h555;
rom[11818] = 12'h444;
rom[11819] = 12'h444;
rom[11820] = 12'h444;
rom[11821] = 12'h444;
rom[11822] = 12'h444;
rom[11823] = 12'h444;
rom[11824] = 12'h444;
rom[11825] = 12'h444;
rom[11826] = 12'h333;
rom[11827] = 12'h444;
rom[11828] = 12'h444;
rom[11829] = 12'h444;
rom[11830] = 12'h444;
rom[11831] = 12'h444;
rom[11832] = 12'h444;
rom[11833] = 12'h444;
rom[11834] = 12'h444;
rom[11835] = 12'h444;
rom[11836] = 12'h555;
rom[11837] = 12'h666;
rom[11838] = 12'h777;
rom[11839] = 12'h777;
rom[11840] = 12'h666;
rom[11841] = 12'h666;
rom[11842] = 12'h555;
rom[11843] = 12'h555;
rom[11844] = 12'h555;
rom[11845] = 12'h555;
rom[11846] = 12'h555;
rom[11847] = 12'h444;
rom[11848] = 12'h444;
rom[11849] = 12'h333;
rom[11850] = 12'h333;
rom[11851] = 12'h333;
rom[11852] = 12'h333;
rom[11853] = 12'h333;
rom[11854] = 12'h333;
rom[11855] = 12'h333;
rom[11856] = 12'h222;
rom[11857] = 12'h222;
rom[11858] = 12'h333;
rom[11859] = 12'h333;
rom[11860] = 12'h333;
rom[11861] = 12'h333;
rom[11862] = 12'h222;
rom[11863] = 12'h222;
rom[11864] = 12'h111;
rom[11865] = 12'h111;
rom[11866] = 12'h111;
rom[11867] = 12'h111;
rom[11868] = 12'h  0;
rom[11869] = 12'h  0;
rom[11870] = 12'h  0;
rom[11871] = 12'h  0;
rom[11872] = 12'h  0;
rom[11873] = 12'h  0;
rom[11874] = 12'h  0;
rom[11875] = 12'h  0;
rom[11876] = 12'h  0;
rom[11877] = 12'h  0;
rom[11878] = 12'h  0;
rom[11879] = 12'h  0;
rom[11880] = 12'h  0;
rom[11881] = 12'h  0;
rom[11882] = 12'h  0;
rom[11883] = 12'h  0;
rom[11884] = 12'h  0;
rom[11885] = 12'h  0;
rom[11886] = 12'h  0;
rom[11887] = 12'h  0;
rom[11888] = 12'h  0;
rom[11889] = 12'h  0;
rom[11890] = 12'h  0;
rom[11891] = 12'h  0;
rom[11892] = 12'h  0;
rom[11893] = 12'h  0;
rom[11894] = 12'h  0;
rom[11895] = 12'h  0;
rom[11896] = 12'h  0;
rom[11897] = 12'h  0;
rom[11898] = 12'h  0;
rom[11899] = 12'h111;
rom[11900] = 12'h111;
rom[11901] = 12'h111;
rom[11902] = 12'h  0;
rom[11903] = 12'h  0;
rom[11904] = 12'h  0;
rom[11905] = 12'h  0;
rom[11906] = 12'h  0;
rom[11907] = 12'h  0;
rom[11908] = 12'h  0;
rom[11909] = 12'h  0;
rom[11910] = 12'h  0;
rom[11911] = 12'h  0;
rom[11912] = 12'h111;
rom[11913] = 12'h111;
rom[11914] = 12'h111;
rom[11915] = 12'h222;
rom[11916] = 12'h333;
rom[11917] = 12'h555;
rom[11918] = 12'h666;
rom[11919] = 12'h666;
rom[11920] = 12'h666;
rom[11921] = 12'h555;
rom[11922] = 12'h333;
rom[11923] = 12'h333;
rom[11924] = 12'h444;
rom[11925] = 12'h444;
rom[11926] = 12'h444;
rom[11927] = 12'h444;
rom[11928] = 12'h333;
rom[11929] = 12'h222;
rom[11930] = 12'h111;
rom[11931] = 12'h111;
rom[11932] = 12'h111;
rom[11933] = 12'h111;
rom[11934] = 12'h111;
rom[11935] = 12'h111;
rom[11936] = 12'h111;
rom[11937] = 12'h  0;
rom[11938] = 12'h  0;
rom[11939] = 12'h  0;
rom[11940] = 12'h  0;
rom[11941] = 12'h  0;
rom[11942] = 12'h  0;
rom[11943] = 12'h  0;
rom[11944] = 12'h  0;
rom[11945] = 12'h111;
rom[11946] = 12'h111;
rom[11947] = 12'h111;
rom[11948] = 12'h111;
rom[11949] = 12'h111;
rom[11950] = 12'h222;
rom[11951] = 12'h333;
rom[11952] = 12'h444;
rom[11953] = 12'h444;
rom[11954] = 12'h555;
rom[11955] = 12'h666;
rom[11956] = 12'h666;
rom[11957] = 12'h666;
rom[11958] = 12'h555;
rom[11959] = 12'h555;
rom[11960] = 12'h555;
rom[11961] = 12'h555;
rom[11962] = 12'h444;
rom[11963] = 12'h444;
rom[11964] = 12'h444;
rom[11965] = 12'h444;
rom[11966] = 12'h444;
rom[11967] = 12'h444;
rom[11968] = 12'h555;
rom[11969] = 12'h555;
rom[11970] = 12'h666;
rom[11971] = 12'h666;
rom[11972] = 12'h666;
rom[11973] = 12'h555;
rom[11974] = 12'h555;
rom[11975] = 12'h444;
rom[11976] = 12'h444;
rom[11977] = 12'h444;
rom[11978] = 12'h444;
rom[11979] = 12'h444;
rom[11980] = 12'h444;
rom[11981] = 12'h444;
rom[11982] = 12'h444;
rom[11983] = 12'h444;
rom[11984] = 12'h444;
rom[11985] = 12'h444;
rom[11986] = 12'h555;
rom[11987] = 12'h555;
rom[11988] = 12'h555;
rom[11989] = 12'h666;
rom[11990] = 12'h666;
rom[11991] = 12'h666;
rom[11992] = 12'h777;
rom[11993] = 12'h888;
rom[11994] = 12'h888;
rom[11995] = 12'h999;
rom[11996] = 12'haaa;
rom[11997] = 12'haaa;
rom[11998] = 12'haaa;
rom[11999] = 12'haaa;
rom[12000] = 12'h222;
rom[12001] = 12'h222;
rom[12002] = 12'h222;
rom[12003] = 12'h222;
rom[12004] = 12'h222;
rom[12005] = 12'h222;
rom[12006] = 12'h222;
rom[12007] = 12'h111;
rom[12008] = 12'h111;
rom[12009] = 12'h111;
rom[12010] = 12'h111;
rom[12011] = 12'h111;
rom[12012] = 12'h111;
rom[12013] = 12'h111;
rom[12014] = 12'h111;
rom[12015] = 12'h111;
rom[12016] = 12'h111;
rom[12017] = 12'h111;
rom[12018] = 12'h111;
rom[12019] = 12'h111;
rom[12020] = 12'h111;
rom[12021] = 12'h111;
rom[12022] = 12'h111;
rom[12023] = 12'h111;
rom[12024] = 12'h111;
rom[12025] = 12'h111;
rom[12026] = 12'h111;
rom[12027] = 12'h111;
rom[12028] = 12'h111;
rom[12029] = 12'h111;
rom[12030] = 12'h111;
rom[12031] = 12'h111;
rom[12032] = 12'h222;
rom[12033] = 12'h222;
rom[12034] = 12'h111;
rom[12035] = 12'h111;
rom[12036] = 12'h222;
rom[12037] = 12'h222;
rom[12038] = 12'h222;
rom[12039] = 12'h222;
rom[12040] = 12'h222;
rom[12041] = 12'h222;
rom[12042] = 12'h222;
rom[12043] = 12'h222;
rom[12044] = 12'h222;
rom[12045] = 12'h222;
rom[12046] = 12'h222;
rom[12047] = 12'h222;
rom[12048] = 12'h222;
rom[12049] = 12'h222;
rom[12050] = 12'h222;
rom[12051] = 12'h222;
rom[12052] = 12'h222;
rom[12053] = 12'h222;
rom[12054] = 12'h222;
rom[12055] = 12'h222;
rom[12056] = 12'h444;
rom[12057] = 12'h444;
rom[12058] = 12'h444;
rom[12059] = 12'h555;
rom[12060] = 12'h555;
rom[12061] = 12'h555;
rom[12062] = 12'h444;
rom[12063] = 12'h444;
rom[12064] = 12'h444;
rom[12065] = 12'h444;
rom[12066] = 12'h555;
rom[12067] = 12'h555;
rom[12068] = 12'h666;
rom[12069] = 12'h666;
rom[12070] = 12'h666;
rom[12071] = 12'h666;
rom[12072] = 12'h666;
rom[12073] = 12'h555;
rom[12074] = 12'h555;
rom[12075] = 12'h444;
rom[12076] = 12'h444;
rom[12077] = 12'h333;
rom[12078] = 12'h333;
rom[12079] = 12'h333;
rom[12080] = 12'h333;
rom[12081] = 12'h333;
rom[12082] = 12'h333;
rom[12083] = 12'h333;
rom[12084] = 12'h222;
rom[12085] = 12'h222;
rom[12086] = 12'h222;
rom[12087] = 12'h111;
rom[12088] = 12'h111;
rom[12089] = 12'h111;
rom[12090] = 12'h111;
rom[12091] = 12'h111;
rom[12092] = 12'h111;
rom[12093] = 12'h111;
rom[12094] = 12'h111;
rom[12095] = 12'h111;
rom[12096] = 12'h111;
rom[12097] = 12'h111;
rom[12098] = 12'h111;
rom[12099] = 12'h111;
rom[12100] = 12'h 11;
rom[12101] = 12'h 11;
rom[12102] = 12'h111;
rom[12103] = 12'h111;
rom[12104] = 12'h111;
rom[12105] = 12'h111;
rom[12106] = 12'h  0;
rom[12107] = 12'h  0;
rom[12108] = 12'h  0;
rom[12109] = 12'h  0;
rom[12110] = 12'h100;
rom[12111] = 12'h100;
rom[12112] = 12'h100;
rom[12113] = 12'h100;
rom[12114] = 12'h200;
rom[12115] = 12'h300;
rom[12116] = 12'h400;
rom[12117] = 12'h510;
rom[12118] = 12'h610;
rom[12119] = 12'h720;
rom[12120] = 12'h820;
rom[12121] = 12'h931;
rom[12122] = 12'ha41;
rom[12123] = 12'ha31;
rom[12124] = 12'h921;
rom[12125] = 12'h820;
rom[12126] = 12'h710;
rom[12127] = 12'h600;
rom[12128] = 12'h500;
rom[12129] = 12'h500;
rom[12130] = 12'h500;
rom[12131] = 12'h500;
rom[12132] = 12'h500;
rom[12133] = 12'h500;
rom[12134] = 12'h500;
rom[12135] = 12'h500;
rom[12136] = 12'h400;
rom[12137] = 12'h400;
rom[12138] = 12'h500;
rom[12139] = 12'h500;
rom[12140] = 12'h400;
rom[12141] = 12'h400;
rom[12142] = 12'h400;
rom[12143] = 12'h400;
rom[12144] = 12'h300;
rom[12145] = 12'h300;
rom[12146] = 12'h300;
rom[12147] = 12'h200;
rom[12148] = 12'h200;
rom[12149] = 12'h200;
rom[12150] = 12'h100;
rom[12151] = 12'h100;
rom[12152] = 12'h100;
rom[12153] = 12'h100;
rom[12154] = 12'h100;
rom[12155] = 12'h100;
rom[12156] = 12'h200;
rom[12157] = 12'h200;
rom[12158] = 12'h200;
rom[12159] = 12'h200;
rom[12160] = 12'h200;
rom[12161] = 12'h100;
rom[12162] = 12'h200;
rom[12163] = 12'h200;
rom[12164] = 12'h200;
rom[12165] = 12'h200;
rom[12166] = 12'h200;
rom[12167] = 12'h200;
rom[12168] = 12'h200;
rom[12169] = 12'h200;
rom[12170] = 12'h200;
rom[12171] = 12'h200;
rom[12172] = 12'h300;
rom[12173] = 12'h300;
rom[12174] = 12'h300;
rom[12175] = 12'h300;
rom[12176] = 12'h400;
rom[12177] = 12'h400;
rom[12178] = 12'h400;
rom[12179] = 12'h300;
rom[12180] = 12'h300;
rom[12181] = 12'h310;
rom[12182] = 12'h311;
rom[12183] = 12'h321;
rom[12184] = 12'h422;
rom[12185] = 12'h533;
rom[12186] = 12'h544;
rom[12187] = 12'h554;
rom[12188] = 12'h665;
rom[12189] = 12'h877;
rom[12190] = 12'h999;
rom[12191] = 12'haaa;
rom[12192] = 12'hbbb;
rom[12193] = 12'hbbb;
rom[12194] = 12'hbbb;
rom[12195] = 12'hbbb;
rom[12196] = 12'haaa;
rom[12197] = 12'h999;
rom[12198] = 12'h999;
rom[12199] = 12'h999;
rom[12200] = 12'haaa;
rom[12201] = 12'haaa;
rom[12202] = 12'h999;
rom[12203] = 12'h999;
rom[12204] = 12'haaa;
rom[12205] = 12'haaa;
rom[12206] = 12'h888;
rom[12207] = 12'h888;
rom[12208] = 12'h777;
rom[12209] = 12'h666;
rom[12210] = 12'h666;
rom[12211] = 12'h777;
rom[12212] = 12'h777;
rom[12213] = 12'h666;
rom[12214] = 12'h555;
rom[12215] = 12'h666;
rom[12216] = 12'h555;
rom[12217] = 12'h555;
rom[12218] = 12'h555;
rom[12219] = 12'h555;
rom[12220] = 12'h555;
rom[12221] = 12'h555;
rom[12222] = 12'h444;
rom[12223] = 12'h444;
rom[12224] = 12'h444;
rom[12225] = 12'h444;
rom[12226] = 12'h444;
rom[12227] = 12'h444;
rom[12228] = 12'h444;
rom[12229] = 12'h555;
rom[12230] = 12'h555;
rom[12231] = 12'h555;
rom[12232] = 12'h555;
rom[12233] = 12'h555;
rom[12234] = 12'h555;
rom[12235] = 12'h666;
rom[12236] = 12'h777;
rom[12237] = 12'h777;
rom[12238] = 12'h777;
rom[12239] = 12'h777;
rom[12240] = 12'h666;
rom[12241] = 12'h666;
rom[12242] = 12'h555;
rom[12243] = 12'h555;
rom[12244] = 12'h555;
rom[12245] = 12'h555;
rom[12246] = 12'h444;
rom[12247] = 12'h444;
rom[12248] = 12'h333;
rom[12249] = 12'h333;
rom[12250] = 12'h333;
rom[12251] = 12'h333;
rom[12252] = 12'h333;
rom[12253] = 12'h333;
rom[12254] = 12'h333;
rom[12255] = 12'h333;
rom[12256] = 12'h333;
rom[12257] = 12'h333;
rom[12258] = 12'h333;
rom[12259] = 12'h333;
rom[12260] = 12'h333;
rom[12261] = 12'h333;
rom[12262] = 12'h222;
rom[12263] = 12'h111;
rom[12264] = 12'h111;
rom[12265] = 12'h111;
rom[12266] = 12'h111;
rom[12267] = 12'h111;
rom[12268] = 12'h  0;
rom[12269] = 12'h  0;
rom[12270] = 12'h  0;
rom[12271] = 12'h  0;
rom[12272] = 12'h  0;
rom[12273] = 12'h  0;
rom[12274] = 12'h  0;
rom[12275] = 12'h  0;
rom[12276] = 12'h  0;
rom[12277] = 12'h  0;
rom[12278] = 12'h  0;
rom[12279] = 12'h  0;
rom[12280] = 12'h  0;
rom[12281] = 12'h  0;
rom[12282] = 12'h  0;
rom[12283] = 12'h  0;
rom[12284] = 12'h  0;
rom[12285] = 12'h  0;
rom[12286] = 12'h  0;
rom[12287] = 12'h  0;
rom[12288] = 12'h  0;
rom[12289] = 12'h  0;
rom[12290] = 12'h  0;
rom[12291] = 12'h  0;
rom[12292] = 12'h  0;
rom[12293] = 12'h  0;
rom[12294] = 12'h  0;
rom[12295] = 12'h  0;
rom[12296] = 12'h  0;
rom[12297] = 12'h  0;
rom[12298] = 12'h  0;
rom[12299] = 12'h111;
rom[12300] = 12'h111;
rom[12301] = 12'h111;
rom[12302] = 12'h  0;
rom[12303] = 12'h  0;
rom[12304] = 12'h  0;
rom[12305] = 12'h  0;
rom[12306] = 12'h  0;
rom[12307] = 12'h  0;
rom[12308] = 12'h  0;
rom[12309] = 12'h  0;
rom[12310] = 12'h  0;
rom[12311] = 12'h111;
rom[12312] = 12'h111;
rom[12313] = 12'h111;
rom[12314] = 12'h222;
rom[12315] = 12'h222;
rom[12316] = 12'h444;
rom[12317] = 12'h666;
rom[12318] = 12'h666;
rom[12319] = 12'h666;
rom[12320] = 12'h555;
rom[12321] = 12'h444;
rom[12322] = 12'h333;
rom[12323] = 12'h444;
rom[12324] = 12'h444;
rom[12325] = 12'h444;
rom[12326] = 12'h444;
rom[12327] = 12'h444;
rom[12328] = 12'h333;
rom[12329] = 12'h222;
rom[12330] = 12'h111;
rom[12331] = 12'h111;
rom[12332] = 12'h111;
rom[12333] = 12'h111;
rom[12334] = 12'h111;
rom[12335] = 12'h111;
rom[12336] = 12'h  0;
rom[12337] = 12'h  0;
rom[12338] = 12'h  0;
rom[12339] = 12'h  0;
rom[12340] = 12'h  0;
rom[12341] = 12'h  0;
rom[12342] = 12'h  0;
rom[12343] = 12'h  0;
rom[12344] = 12'h  0;
rom[12345] = 12'h  0;
rom[12346] = 12'h111;
rom[12347] = 12'h111;
rom[12348] = 12'h111;
rom[12349] = 12'h111;
rom[12350] = 12'h222;
rom[12351] = 12'h333;
rom[12352] = 12'h444;
rom[12353] = 12'h555;
rom[12354] = 12'h555;
rom[12355] = 12'h666;
rom[12356] = 12'h666;
rom[12357] = 12'h666;
rom[12358] = 12'h555;
rom[12359] = 12'h555;
rom[12360] = 12'h555;
rom[12361] = 12'h444;
rom[12362] = 12'h444;
rom[12363] = 12'h444;
rom[12364] = 12'h444;
rom[12365] = 12'h555;
rom[12366] = 12'h555;
rom[12367] = 12'h555;
rom[12368] = 12'h555;
rom[12369] = 12'h555;
rom[12370] = 12'h555;
rom[12371] = 12'h555;
rom[12372] = 12'h444;
rom[12373] = 12'h444;
rom[12374] = 12'h444;
rom[12375] = 12'h444;
rom[12376] = 12'h444;
rom[12377] = 12'h444;
rom[12378] = 12'h444;
rom[12379] = 12'h444;
rom[12380] = 12'h444;
rom[12381] = 12'h444;
rom[12382] = 12'h444;
rom[12383] = 12'h444;
rom[12384] = 12'h444;
rom[12385] = 12'h444;
rom[12386] = 12'h444;
rom[12387] = 12'h555;
rom[12388] = 12'h555;
rom[12389] = 12'h555;
rom[12390] = 12'h666;
rom[12391] = 12'h666;
rom[12392] = 12'h777;
rom[12393] = 12'h888;
rom[12394] = 12'h888;
rom[12395] = 12'h999;
rom[12396] = 12'haaa;
rom[12397] = 12'haaa;
rom[12398] = 12'haaa;
rom[12399] = 12'haaa;
rom[12400] = 12'h222;
rom[12401] = 12'h222;
rom[12402] = 12'h111;
rom[12403] = 12'h111;
rom[12404] = 12'h111;
rom[12405] = 12'h111;
rom[12406] = 12'h111;
rom[12407] = 12'h111;
rom[12408] = 12'h111;
rom[12409] = 12'h111;
rom[12410] = 12'h111;
rom[12411] = 12'h111;
rom[12412] = 12'h111;
rom[12413] = 12'h111;
rom[12414] = 12'h111;
rom[12415] = 12'h222;
rom[12416] = 12'h111;
rom[12417] = 12'h111;
rom[12418] = 12'h111;
rom[12419] = 12'h111;
rom[12420] = 12'h111;
rom[12421] = 12'h111;
rom[12422] = 12'h111;
rom[12423] = 12'h111;
rom[12424] = 12'h111;
rom[12425] = 12'h111;
rom[12426] = 12'h111;
rom[12427] = 12'h111;
rom[12428] = 12'h111;
rom[12429] = 12'h111;
rom[12430] = 12'h222;
rom[12431] = 12'h222;
rom[12432] = 12'h222;
rom[12433] = 12'h222;
rom[12434] = 12'h222;
rom[12435] = 12'h222;
rom[12436] = 12'h222;
rom[12437] = 12'h222;
rom[12438] = 12'h222;
rom[12439] = 12'h222;
rom[12440] = 12'h222;
rom[12441] = 12'h222;
rom[12442] = 12'h222;
rom[12443] = 12'h222;
rom[12444] = 12'h222;
rom[12445] = 12'h222;
rom[12446] = 12'h222;
rom[12447] = 12'h222;
rom[12448] = 12'h222;
rom[12449] = 12'h222;
rom[12450] = 12'h222;
rom[12451] = 12'h222;
rom[12452] = 12'h222;
rom[12453] = 12'h222;
rom[12454] = 12'h333;
rom[12455] = 12'h333;
rom[12456] = 12'h333;
rom[12457] = 12'h444;
rom[12458] = 12'h444;
rom[12459] = 12'h555;
rom[12460] = 12'h555;
rom[12461] = 12'h555;
rom[12462] = 12'h444;
rom[12463] = 12'h444;
rom[12464] = 12'h444;
rom[12465] = 12'h444;
rom[12466] = 12'h444;
rom[12467] = 12'h555;
rom[12468] = 12'h555;
rom[12469] = 12'h666;
rom[12470] = 12'h666;
rom[12471] = 12'h666;
rom[12472] = 12'h777;
rom[12473] = 12'h666;
rom[12474] = 12'h555;
rom[12475] = 12'h555;
rom[12476] = 12'h444;
rom[12477] = 12'h444;
rom[12478] = 12'h333;
rom[12479] = 12'h333;
rom[12480] = 12'h333;
rom[12481] = 12'h333;
rom[12482] = 12'h333;
rom[12483] = 12'h333;
rom[12484] = 12'h333;
rom[12485] = 12'h222;
rom[12486] = 12'h222;
rom[12487] = 12'h111;
rom[12488] = 12'h111;
rom[12489] = 12'h111;
rom[12490] = 12'h111;
rom[12491] = 12'h111;
rom[12492] = 12'h111;
rom[12493] = 12'h111;
rom[12494] = 12'h111;
rom[12495] = 12'h111;
rom[12496] = 12'h111;
rom[12497] = 12'h111;
rom[12498] = 12'h111;
rom[12499] = 12'h111;
rom[12500] = 12'h 11;
rom[12501] = 12'h 11;
rom[12502] = 12'h 11;
rom[12503] = 12'h 11;
rom[12504] = 12'h111;
rom[12505] = 12'h  0;
rom[12506] = 12'h  0;
rom[12507] = 12'h  0;
rom[12508] = 12'h  0;
rom[12509] = 12'h  0;
rom[12510] = 12'h  0;
rom[12511] = 12'h100;
rom[12512] = 12'h100;
rom[12513] = 12'h100;
rom[12514] = 12'h200;
rom[12515] = 12'h300;
rom[12516] = 12'h400;
rom[12517] = 12'h510;
rom[12518] = 12'h610;
rom[12519] = 12'h720;
rom[12520] = 12'h820;
rom[12521] = 12'h931;
rom[12522] = 12'ha41;
rom[12523] = 12'ha31;
rom[12524] = 12'h931;
rom[12525] = 12'h820;
rom[12526] = 12'h710;
rom[12527] = 12'h600;
rom[12528] = 12'h500;
rom[12529] = 12'h500;
rom[12530] = 12'h500;
rom[12531] = 12'h500;
rom[12532] = 12'h500;
rom[12533] = 12'h500;
rom[12534] = 12'h500;
rom[12535] = 12'h500;
rom[12536] = 12'h500;
rom[12537] = 12'h400;
rom[12538] = 12'h500;
rom[12539] = 12'h400;
rom[12540] = 12'h400;
rom[12541] = 12'h400;
rom[12542] = 12'h400;
rom[12543] = 12'h400;
rom[12544] = 12'h300;
rom[12545] = 12'h300;
rom[12546] = 12'h200;
rom[12547] = 12'h200;
rom[12548] = 12'h200;
rom[12549] = 12'h100;
rom[12550] = 12'h100;
rom[12551] = 12'h100;
rom[12552] = 12'h100;
rom[12553] = 12'h100;
rom[12554] = 12'h100;
rom[12555] = 12'h100;
rom[12556] = 12'h100;
rom[12557] = 12'h100;
rom[12558] = 12'h100;
rom[12559] = 12'h100;
rom[12560] = 12'h100;
rom[12561] = 12'h100;
rom[12562] = 12'h100;
rom[12563] = 12'h100;
rom[12564] = 12'h200;
rom[12565] = 12'h200;
rom[12566] = 12'h200;
rom[12567] = 12'h200;
rom[12568] = 12'h200;
rom[12569] = 12'h200;
rom[12570] = 12'h200;
rom[12571] = 12'h200;
rom[12572] = 12'h200;
rom[12573] = 12'h300;
rom[12574] = 12'h300;
rom[12575] = 12'h300;
rom[12576] = 12'h400;
rom[12577] = 12'h400;
rom[12578] = 12'h400;
rom[12579] = 12'h400;
rom[12580] = 12'h410;
rom[12581] = 12'h410;
rom[12582] = 12'h310;
rom[12583] = 12'h310;
rom[12584] = 12'h310;
rom[12585] = 12'h422;
rom[12586] = 12'h543;
rom[12587] = 12'h544;
rom[12588] = 12'h554;
rom[12589] = 12'h666;
rom[12590] = 12'h887;
rom[12591] = 12'h999;
rom[12592] = 12'hbbb;
rom[12593] = 12'hbbb;
rom[12594] = 12'hbbb;
rom[12595] = 12'hbbb;
rom[12596] = 12'hbaa;
rom[12597] = 12'haaa;
rom[12598] = 12'h999;
rom[12599] = 12'h999;
rom[12600] = 12'haaa;
rom[12601] = 12'haaa;
rom[12602] = 12'haaa;
rom[12603] = 12'h999;
rom[12604] = 12'haaa;
rom[12605] = 12'haaa;
rom[12606] = 12'h999;
rom[12607] = 12'h888;
rom[12608] = 12'h777;
rom[12609] = 12'h677;
rom[12610] = 12'h666;
rom[12611] = 12'h777;
rom[12612] = 12'h777;
rom[12613] = 12'h666;
rom[12614] = 12'h666;
rom[12615] = 12'h666;
rom[12616] = 12'h666;
rom[12617] = 12'h555;
rom[12618] = 12'h555;
rom[12619] = 12'h555;
rom[12620] = 12'h555;
rom[12621] = 12'h555;
rom[12622] = 12'h555;
rom[12623] = 12'h555;
rom[12624] = 12'h555;
rom[12625] = 12'h555;
rom[12626] = 12'h555;
rom[12627] = 12'h555;
rom[12628] = 12'h555;
rom[12629] = 12'h555;
rom[12630] = 12'h555;
rom[12631] = 12'h666;
rom[12632] = 12'h666;
rom[12633] = 12'h666;
rom[12634] = 12'h777;
rom[12635] = 12'h777;
rom[12636] = 12'h777;
rom[12637] = 12'h777;
rom[12638] = 12'h777;
rom[12639] = 12'h666;
rom[12640] = 12'h666;
rom[12641] = 12'h666;
rom[12642] = 12'h555;
rom[12643] = 12'h444;
rom[12644] = 12'h444;
rom[12645] = 12'h444;
rom[12646] = 12'h333;
rom[12647] = 12'h333;
rom[12648] = 12'h333;
rom[12649] = 12'h333;
rom[12650] = 12'h333;
rom[12651] = 12'h333;
rom[12652] = 12'h333;
rom[12653] = 12'h333;
rom[12654] = 12'h333;
rom[12655] = 12'h222;
rom[12656] = 12'h444;
rom[12657] = 12'h444;
rom[12658] = 12'h333;
rom[12659] = 12'h333;
rom[12660] = 12'h333;
rom[12661] = 12'h222;
rom[12662] = 12'h222;
rom[12663] = 12'h111;
rom[12664] = 12'h111;
rom[12665] = 12'h111;
rom[12666] = 12'h111;
rom[12667] = 12'h  0;
rom[12668] = 12'h  0;
rom[12669] = 12'h  0;
rom[12670] = 12'h  0;
rom[12671] = 12'h  0;
rom[12672] = 12'h  0;
rom[12673] = 12'h  0;
rom[12674] = 12'h  0;
rom[12675] = 12'h  0;
rom[12676] = 12'h  0;
rom[12677] = 12'h  0;
rom[12678] = 12'h  0;
rom[12679] = 12'h  0;
rom[12680] = 12'h  0;
rom[12681] = 12'h  0;
rom[12682] = 12'h  0;
rom[12683] = 12'h  0;
rom[12684] = 12'h  0;
rom[12685] = 12'h  0;
rom[12686] = 12'h  0;
rom[12687] = 12'h  0;
rom[12688] = 12'h  0;
rom[12689] = 12'h  0;
rom[12690] = 12'h  0;
rom[12691] = 12'h  0;
rom[12692] = 12'h  0;
rom[12693] = 12'h  0;
rom[12694] = 12'h  0;
rom[12695] = 12'h  0;
rom[12696] = 12'h  0;
rom[12697] = 12'h  0;
rom[12698] = 12'h  0;
rom[12699] = 12'h111;
rom[12700] = 12'h111;
rom[12701] = 12'h111;
rom[12702] = 12'h  0;
rom[12703] = 12'h  0;
rom[12704] = 12'h  0;
rom[12705] = 12'h  0;
rom[12706] = 12'h  0;
rom[12707] = 12'h  0;
rom[12708] = 12'h  0;
rom[12709] = 12'h  0;
rom[12710] = 12'h  0;
rom[12711] = 12'h111;
rom[12712] = 12'h111;
rom[12713] = 12'h222;
rom[12714] = 12'h222;
rom[12715] = 12'h333;
rom[12716] = 12'h444;
rom[12717] = 12'h666;
rom[12718] = 12'h666;
rom[12719] = 12'h555;
rom[12720] = 12'h555;
rom[12721] = 12'h444;
rom[12722] = 12'h333;
rom[12723] = 12'h444;
rom[12724] = 12'h444;
rom[12725] = 12'h444;
rom[12726] = 12'h444;
rom[12727] = 12'h444;
rom[12728] = 12'h333;
rom[12729] = 12'h222;
rom[12730] = 12'h111;
rom[12731] = 12'h111;
rom[12732] = 12'h111;
rom[12733] = 12'h111;
rom[12734] = 12'h111;
rom[12735] = 12'h  0;
rom[12736] = 12'h  0;
rom[12737] = 12'h  0;
rom[12738] = 12'h  0;
rom[12739] = 12'h  0;
rom[12740] = 12'h  0;
rom[12741] = 12'h  0;
rom[12742] = 12'h  0;
rom[12743] = 12'h  0;
rom[12744] = 12'h  0;
rom[12745] = 12'h  0;
rom[12746] = 12'h111;
rom[12747] = 12'h111;
rom[12748] = 12'h111;
rom[12749] = 12'h111;
rom[12750] = 12'h222;
rom[12751] = 12'h333;
rom[12752] = 12'h444;
rom[12753] = 12'h555;
rom[12754] = 12'h666;
rom[12755] = 12'h666;
rom[12756] = 12'h666;
rom[12757] = 12'h666;
rom[12758] = 12'h555;
rom[12759] = 12'h555;
rom[12760] = 12'h444;
rom[12761] = 12'h444;
rom[12762] = 12'h444;
rom[12763] = 12'h555;
rom[12764] = 12'h555;
rom[12765] = 12'h555;
rom[12766] = 12'h666;
rom[12767] = 12'h666;
rom[12768] = 12'h666;
rom[12769] = 12'h666;
rom[12770] = 12'h555;
rom[12771] = 12'h444;
rom[12772] = 12'h444;
rom[12773] = 12'h333;
rom[12774] = 12'h333;
rom[12775] = 12'h333;
rom[12776] = 12'h444;
rom[12777] = 12'h444;
rom[12778] = 12'h444;
rom[12779] = 12'h333;
rom[12780] = 12'h444;
rom[12781] = 12'h444;
rom[12782] = 12'h444;
rom[12783] = 12'h444;
rom[12784] = 12'h444;
rom[12785] = 12'h555;
rom[12786] = 12'h555;
rom[12787] = 12'h555;
rom[12788] = 12'h555;
rom[12789] = 12'h555;
rom[12790] = 12'h666;
rom[12791] = 12'h777;
rom[12792] = 12'h777;
rom[12793] = 12'h888;
rom[12794] = 12'h888;
rom[12795] = 12'h999;
rom[12796] = 12'haaa;
rom[12797] = 12'haaa;
rom[12798] = 12'haaa;
rom[12799] = 12'haaa;
rom[12800] = 12'h222;
rom[12801] = 12'h222;
rom[12802] = 12'h222;
rom[12803] = 12'h222;
rom[12804] = 12'h222;
rom[12805] = 12'h111;
rom[12806] = 12'h111;
rom[12807] = 12'h111;
rom[12808] = 12'h111;
rom[12809] = 12'h111;
rom[12810] = 12'h111;
rom[12811] = 12'h111;
rom[12812] = 12'h111;
rom[12813] = 12'h111;
rom[12814] = 12'h111;
rom[12815] = 12'h111;
rom[12816] = 12'h111;
rom[12817] = 12'h111;
rom[12818] = 12'h111;
rom[12819] = 12'h222;
rom[12820] = 12'h222;
rom[12821] = 12'h111;
rom[12822] = 12'h111;
rom[12823] = 12'h111;
rom[12824] = 12'h111;
rom[12825] = 12'h111;
rom[12826] = 12'h111;
rom[12827] = 12'h111;
rom[12828] = 12'h111;
rom[12829] = 12'h222;
rom[12830] = 12'h222;
rom[12831] = 12'h222;
rom[12832] = 12'h222;
rom[12833] = 12'h222;
rom[12834] = 12'h222;
rom[12835] = 12'h222;
rom[12836] = 12'h222;
rom[12837] = 12'h222;
rom[12838] = 12'h222;
rom[12839] = 12'h222;
rom[12840] = 12'h222;
rom[12841] = 12'h222;
rom[12842] = 12'h222;
rom[12843] = 12'h222;
rom[12844] = 12'h333;
rom[12845] = 12'h222;
rom[12846] = 12'h222;
rom[12847] = 12'h222;
rom[12848] = 12'h222;
rom[12849] = 12'h333;
rom[12850] = 12'h333;
rom[12851] = 12'h333;
rom[12852] = 12'h333;
rom[12853] = 12'h333;
rom[12854] = 12'h333;
rom[12855] = 12'h333;
rom[12856] = 12'h333;
rom[12857] = 12'h444;
rom[12858] = 12'h444;
rom[12859] = 12'h444;
rom[12860] = 12'h555;
rom[12861] = 12'h555;
rom[12862] = 12'h555;
rom[12863] = 12'h555;
rom[12864] = 12'h444;
rom[12865] = 12'h444;
rom[12866] = 12'h444;
rom[12867] = 12'h444;
rom[12868] = 12'h555;
rom[12869] = 12'h555;
rom[12870] = 12'h666;
rom[12871] = 12'h666;
rom[12872] = 12'h777;
rom[12873] = 12'h666;
rom[12874] = 12'h666;
rom[12875] = 12'h666;
rom[12876] = 12'h666;
rom[12877] = 12'h666;
rom[12878] = 12'h555;
rom[12879] = 12'h444;
rom[12880] = 12'h333;
rom[12881] = 12'h333;
rom[12882] = 12'h333;
rom[12883] = 12'h333;
rom[12884] = 12'h222;
rom[12885] = 12'h222;
rom[12886] = 12'h222;
rom[12887] = 12'h222;
rom[12888] = 12'h222;
rom[12889] = 12'h222;
rom[12890] = 12'h111;
rom[12891] = 12'h111;
rom[12892] = 12'h111;
rom[12893] = 12'h111;
rom[12894] = 12'h111;
rom[12895] = 12'h  0;
rom[12896] = 12'h111;
rom[12897] = 12'h111;
rom[12898] = 12'h111;
rom[12899] = 12'h111;
rom[12900] = 12'h111;
rom[12901] = 12'h  0;
rom[12902] = 12'h  0;
rom[12903] = 12'h  0;
rom[12904] = 12'h  0;
rom[12905] = 12'h  0;
rom[12906] = 12'h  0;
rom[12907] = 12'h  0;
rom[12908] = 12'h  0;
rom[12909] = 12'h  0;
rom[12910] = 12'h  0;
rom[12911] = 12'h  0;
rom[12912] = 12'h100;
rom[12913] = 12'h100;
rom[12914] = 12'h200;
rom[12915] = 12'h300;
rom[12916] = 12'h400;
rom[12917] = 12'h500;
rom[12918] = 12'h610;
rom[12919] = 12'h720;
rom[12920] = 12'h930;
rom[12921] = 12'h930;
rom[12922] = 12'h930;
rom[12923] = 12'h931;
rom[12924] = 12'ha31;
rom[12925] = 12'h920;
rom[12926] = 12'h810;
rom[12927] = 12'h710;
rom[12928] = 12'h500;
rom[12929] = 12'h500;
rom[12930] = 12'h400;
rom[12931] = 12'h500;
rom[12932] = 12'h500;
rom[12933] = 12'h500;
rom[12934] = 12'h500;
rom[12935] = 12'h400;
rom[12936] = 12'h400;
rom[12937] = 12'h400;
rom[12938] = 12'h400;
rom[12939] = 12'h400;
rom[12940] = 12'h400;
rom[12941] = 12'h300;
rom[12942] = 12'h300;
rom[12943] = 12'h300;
rom[12944] = 12'h200;
rom[12945] = 12'h200;
rom[12946] = 12'h200;
rom[12947] = 12'h200;
rom[12948] = 12'h100;
rom[12949] = 12'h100;
rom[12950] = 12'h100;
rom[12951] = 12'h100;
rom[12952] = 12'h100;
rom[12953] = 12'h100;
rom[12954] = 12'h  0;
rom[12955] = 12'h100;
rom[12956] = 12'h100;
rom[12957] = 12'h100;
rom[12958] = 12'h100;
rom[12959] = 12'h100;
rom[12960] = 12'h100;
rom[12961] = 12'h100;
rom[12962] = 12'h100;
rom[12963] = 12'h100;
rom[12964] = 12'h100;
rom[12965] = 12'h100;
rom[12966] = 12'h100;
rom[12967] = 12'h100;
rom[12968] = 12'h100;
rom[12969] = 12'h200;
rom[12970] = 12'h200;
rom[12971] = 12'h200;
rom[12972] = 12'h200;
rom[12973] = 12'h200;
rom[12974] = 12'h300;
rom[12975] = 12'h300;
rom[12976] = 12'h300;
rom[12977] = 12'h300;
rom[12978] = 12'h400;
rom[12979] = 12'h400;
rom[12980] = 12'h400;
rom[12981] = 12'h400;
rom[12982] = 12'h400;
rom[12983] = 12'h300;
rom[12984] = 12'h300;
rom[12985] = 12'h310;
rom[12986] = 12'h421;
rom[12987] = 12'h432;
rom[12988] = 12'h543;
rom[12989] = 12'h665;
rom[12990] = 12'h776;
rom[12991] = 12'h787;
rom[12992] = 12'h999;
rom[12993] = 12'haaa;
rom[12994] = 12'hbbb;
rom[12995] = 12'hccc;
rom[12996] = 12'hccc;
rom[12997] = 12'hbbb;
rom[12998] = 12'haaa;
rom[12999] = 12'ha99;
rom[13000] = 12'haaa;
rom[13001] = 12'haaa;
rom[13002] = 12'haaa;
rom[13003] = 12'haaa;
rom[13004] = 12'haaa;
rom[13005] = 12'haaa;
rom[13006] = 12'h999;
rom[13007] = 12'h888;
rom[13008] = 12'h777;
rom[13009] = 12'h777;
rom[13010] = 12'h777;
rom[13011] = 12'h777;
rom[13012] = 12'h777;
rom[13013] = 12'h777;
rom[13014] = 12'h677;
rom[13015] = 12'h666;
rom[13016] = 12'h666;
rom[13017] = 12'h666;
rom[13018] = 12'h666;
rom[13019] = 12'h666;
rom[13020] = 12'h666;
rom[13021] = 12'h666;
rom[13022] = 12'h666;
rom[13023] = 12'h666;
rom[13024] = 12'h666;
rom[13025] = 12'h666;
rom[13026] = 12'h666;
rom[13027] = 12'h666;
rom[13028] = 12'h666;
rom[13029] = 12'h666;
rom[13030] = 12'h666;
rom[13031] = 12'h666;
rom[13032] = 12'h777;
rom[13033] = 12'h777;
rom[13034] = 12'h888;
rom[13035] = 12'h888;
rom[13036] = 12'h888;
rom[13037] = 12'h777;
rom[13038] = 12'h777;
rom[13039] = 12'h666;
rom[13040] = 12'h666;
rom[13041] = 12'h555;
rom[13042] = 12'h444;
rom[13043] = 12'h444;
rom[13044] = 12'h444;
rom[13045] = 12'h444;
rom[13046] = 12'h444;
rom[13047] = 12'h444;
rom[13048] = 12'h333;
rom[13049] = 12'h333;
rom[13050] = 12'h333;
rom[13051] = 12'h333;
rom[13052] = 12'h333;
rom[13053] = 12'h444;
rom[13054] = 12'h444;
rom[13055] = 12'h555;
rom[13056] = 12'h444;
rom[13057] = 12'h444;
rom[13058] = 12'h333;
rom[13059] = 12'h333;
rom[13060] = 12'h222;
rom[13061] = 12'h222;
rom[13062] = 12'h111;
rom[13063] = 12'h111;
rom[13064] = 12'h111;
rom[13065] = 12'h111;
rom[13066] = 12'h  0;
rom[13067] = 12'h  0;
rom[13068] = 12'h  0;
rom[13069] = 12'h  0;
rom[13070] = 12'h  0;
rom[13071] = 12'h  0;
rom[13072] = 12'h  0;
rom[13073] = 12'h  0;
rom[13074] = 12'h  0;
rom[13075] = 12'h  0;
rom[13076] = 12'h  0;
rom[13077] = 12'h  0;
rom[13078] = 12'h  0;
rom[13079] = 12'h  0;
rom[13080] = 12'h  0;
rom[13081] = 12'h  0;
rom[13082] = 12'h  0;
rom[13083] = 12'h  0;
rom[13084] = 12'h  0;
rom[13085] = 12'h  0;
rom[13086] = 12'h  0;
rom[13087] = 12'h  0;
rom[13088] = 12'h  0;
rom[13089] = 12'h  0;
rom[13090] = 12'h  0;
rom[13091] = 12'h  0;
rom[13092] = 12'h  0;
rom[13093] = 12'h  0;
rom[13094] = 12'h  0;
rom[13095] = 12'h  0;
rom[13096] = 12'h  0;
rom[13097] = 12'h  0;
rom[13098] = 12'h111;
rom[13099] = 12'h111;
rom[13100] = 12'h111;
rom[13101] = 12'h  0;
rom[13102] = 12'h  0;
rom[13103] = 12'h  0;
rom[13104] = 12'h  0;
rom[13105] = 12'h  0;
rom[13106] = 12'h  0;
rom[13107] = 12'h  0;
rom[13108] = 12'h  0;
rom[13109] = 12'h  0;
rom[13110] = 12'h111;
rom[13111] = 12'h111;
rom[13112] = 12'h111;
rom[13113] = 12'h222;
rom[13114] = 12'h333;
rom[13115] = 12'h444;
rom[13116] = 12'h555;
rom[13117] = 12'h555;
rom[13118] = 12'h555;
rom[13119] = 12'h666;
rom[13120] = 12'h555;
rom[13121] = 12'h444;
rom[13122] = 12'h333;
rom[13123] = 12'h333;
rom[13124] = 12'h444;
rom[13125] = 12'h444;
rom[13126] = 12'h444;
rom[13127] = 12'h444;
rom[13128] = 12'h333;
rom[13129] = 12'h222;
rom[13130] = 12'h111;
rom[13131] = 12'h111;
rom[13132] = 12'h111;
rom[13133] = 12'h  0;
rom[13134] = 12'h  0;
rom[13135] = 12'h  0;
rom[13136] = 12'h  0;
rom[13137] = 12'h  0;
rom[13138] = 12'h  0;
rom[13139] = 12'h  0;
rom[13140] = 12'h  0;
rom[13141] = 12'h  0;
rom[13142] = 12'h  0;
rom[13143] = 12'h  0;
rom[13144] = 12'h  0;
rom[13145] = 12'h  0;
rom[13146] = 12'h111;
rom[13147] = 12'h111;
rom[13148] = 12'h111;
rom[13149] = 12'h111;
rom[13150] = 12'h222;
rom[13151] = 12'h333;
rom[13152] = 12'h555;
rom[13153] = 12'h555;
rom[13154] = 12'h666;
rom[13155] = 12'h666;
rom[13156] = 12'h666;
rom[13157] = 12'h666;
rom[13158] = 12'h555;
rom[13159] = 12'h555;
rom[13160] = 12'h444;
rom[13161] = 12'h555;
rom[13162] = 12'h555;
rom[13163] = 12'h555;
rom[13164] = 12'h555;
rom[13165] = 12'h555;
rom[13166] = 12'h555;
rom[13167] = 12'h555;
rom[13168] = 12'h555;
rom[13169] = 12'h555;
rom[13170] = 12'h444;
rom[13171] = 12'h444;
rom[13172] = 12'h444;
rom[13173] = 12'h444;
rom[13174] = 12'h444;
rom[13175] = 12'h444;
rom[13176] = 12'h444;
rom[13177] = 12'h444;
rom[13178] = 12'h444;
rom[13179] = 12'h444;
rom[13180] = 12'h444;
rom[13181] = 12'h444;
rom[13182] = 12'h444;
rom[13183] = 12'h444;
rom[13184] = 12'h444;
rom[13185] = 12'h444;
rom[13186] = 12'h555;
rom[13187] = 12'h555;
rom[13188] = 12'h555;
rom[13189] = 12'h666;
rom[13190] = 12'h666;
rom[13191] = 12'h777;
rom[13192] = 12'h888;
rom[13193] = 12'h888;
rom[13194] = 12'h999;
rom[13195] = 12'h999;
rom[13196] = 12'haaa;
rom[13197] = 12'haaa;
rom[13198] = 12'haaa;
rom[13199] = 12'haaa;
rom[13200] = 12'h222;
rom[13201] = 12'h222;
rom[13202] = 12'h222;
rom[13203] = 12'h222;
rom[13204] = 12'h222;
rom[13205] = 12'h111;
rom[13206] = 12'h111;
rom[13207] = 12'h111;
rom[13208] = 12'h111;
rom[13209] = 12'h111;
rom[13210] = 12'h111;
rom[13211] = 12'h111;
rom[13212] = 12'h111;
rom[13213] = 12'h111;
rom[13214] = 12'h111;
rom[13215] = 12'h111;
rom[13216] = 12'h111;
rom[13217] = 12'h111;
rom[13218] = 12'h111;
rom[13219] = 12'h222;
rom[13220] = 12'h222;
rom[13221] = 12'h222;
rom[13222] = 12'h222;
rom[13223] = 12'h222;
rom[13224] = 12'h111;
rom[13225] = 12'h111;
rom[13226] = 12'h111;
rom[13227] = 12'h111;
rom[13228] = 12'h111;
rom[13229] = 12'h222;
rom[13230] = 12'h222;
rom[13231] = 12'h222;
rom[13232] = 12'h222;
rom[13233] = 12'h222;
rom[13234] = 12'h222;
rom[13235] = 12'h222;
rom[13236] = 12'h222;
rom[13237] = 12'h222;
rom[13238] = 12'h222;
rom[13239] = 12'h222;
rom[13240] = 12'h222;
rom[13241] = 12'h222;
rom[13242] = 12'h222;
rom[13243] = 12'h333;
rom[13244] = 12'h333;
rom[13245] = 12'h333;
rom[13246] = 12'h333;
rom[13247] = 12'h333;
rom[13248] = 12'h333;
rom[13249] = 12'h333;
rom[13250] = 12'h333;
rom[13251] = 12'h333;
rom[13252] = 12'h333;
rom[13253] = 12'h444;
rom[13254] = 12'h444;
rom[13255] = 12'h444;
rom[13256] = 12'h444;
rom[13257] = 12'h444;
rom[13258] = 12'h444;
rom[13259] = 12'h444;
rom[13260] = 12'h555;
rom[13261] = 12'h555;
rom[13262] = 12'h555;
rom[13263] = 12'h555;
rom[13264] = 12'h555;
rom[13265] = 12'h555;
rom[13266] = 12'h555;
rom[13267] = 12'h444;
rom[13268] = 12'h444;
rom[13269] = 12'h555;
rom[13270] = 12'h555;
rom[13271] = 12'h666;
rom[13272] = 12'h777;
rom[13273] = 12'h666;
rom[13274] = 12'h666;
rom[13275] = 12'h666;
rom[13276] = 12'h666;
rom[13277] = 12'h666;
rom[13278] = 12'h555;
rom[13279] = 12'h555;
rom[13280] = 12'h444;
rom[13281] = 12'h444;
rom[13282] = 12'h333;
rom[13283] = 12'h333;
rom[13284] = 12'h333;
rom[13285] = 12'h222;
rom[13286] = 12'h222;
rom[13287] = 12'h222;
rom[13288] = 12'h222;
rom[13289] = 12'h222;
rom[13290] = 12'h111;
rom[13291] = 12'h111;
rom[13292] = 12'h111;
rom[13293] = 12'h111;
rom[13294] = 12'h111;
rom[13295] = 12'h111;
rom[13296] = 12'h111;
rom[13297] = 12'h111;
rom[13298] = 12'h111;
rom[13299] = 12'h111;
rom[13300] = 12'h111;
rom[13301] = 12'h  0;
rom[13302] = 12'h  0;
rom[13303] = 12'h  0;
rom[13304] = 12'h  0;
rom[13305] = 12'h  0;
rom[13306] = 12'h  0;
rom[13307] = 12'h  0;
rom[13308] = 12'h  0;
rom[13309] = 12'h  0;
rom[13310] = 12'h  0;
rom[13311] = 12'h  0;
rom[13312] = 12'h100;
rom[13313] = 12'h100;
rom[13314] = 12'h200;
rom[13315] = 12'h300;
rom[13316] = 12'h400;
rom[13317] = 12'h500;
rom[13318] = 12'h610;
rom[13319] = 12'h720;
rom[13320] = 12'h830;
rom[13321] = 12'h930;
rom[13322] = 12'h930;
rom[13323] = 12'ha31;
rom[13324] = 12'ha31;
rom[13325] = 12'h920;
rom[13326] = 12'h810;
rom[13327] = 12'h710;
rom[13328] = 12'h500;
rom[13329] = 12'h400;
rom[13330] = 12'h400;
rom[13331] = 12'h500;
rom[13332] = 12'h500;
rom[13333] = 12'h500;
rom[13334] = 12'h400;
rom[13335] = 12'h400;
rom[13336] = 12'h400;
rom[13337] = 12'h400;
rom[13338] = 12'h400;
rom[13339] = 12'h400;
rom[13340] = 12'h300;
rom[13341] = 12'h300;
rom[13342] = 12'h300;
rom[13343] = 12'h300;
rom[13344] = 12'h200;
rom[13345] = 12'h200;
rom[13346] = 12'h200;
rom[13347] = 12'h100;
rom[13348] = 12'h100;
rom[13349] = 12'h100;
rom[13350] = 12'h100;
rom[13351] = 12'h100;
rom[13352] = 12'h  0;
rom[13353] = 12'h  0;
rom[13354] = 12'h  0;
rom[13355] = 12'h  0;
rom[13356] = 12'h  0;
rom[13357] = 12'h  0;
rom[13358] = 12'h  0;
rom[13359] = 12'h100;
rom[13360] = 12'h100;
rom[13361] = 12'h100;
rom[13362] = 12'h100;
rom[13363] = 12'h100;
rom[13364] = 12'h100;
rom[13365] = 12'h100;
rom[13366] = 12'h100;
rom[13367] = 12'h100;
rom[13368] = 12'h100;
rom[13369] = 12'h100;
rom[13370] = 12'h200;
rom[13371] = 12'h200;
rom[13372] = 12'h200;
rom[13373] = 12'h200;
rom[13374] = 12'h300;
rom[13375] = 12'h300;
rom[13376] = 12'h300;
rom[13377] = 12'h300;
rom[13378] = 12'h400;
rom[13379] = 12'h400;
rom[13380] = 12'h400;
rom[13381] = 12'h400;
rom[13382] = 12'h400;
rom[13383] = 12'h400;
rom[13384] = 12'h300;
rom[13385] = 12'h310;
rom[13386] = 12'h311;
rom[13387] = 12'h422;
rom[13388] = 12'h433;
rom[13389] = 12'h554;
rom[13390] = 12'h665;
rom[13391] = 12'h776;
rom[13392] = 12'h998;
rom[13393] = 12'ha99;
rom[13394] = 12'hbbb;
rom[13395] = 12'hccc;
rom[13396] = 12'hccc;
rom[13397] = 12'hcbc;
rom[13398] = 12'hbbb;
rom[13399] = 12'haaa;
rom[13400] = 12'haaa;
rom[13401] = 12'haaa;
rom[13402] = 12'haaa;
rom[13403] = 12'haaa;
rom[13404] = 12'haaa;
rom[13405] = 12'haaa;
rom[13406] = 12'h999;
rom[13407] = 12'h888;
rom[13408] = 12'h788;
rom[13409] = 12'h777;
rom[13410] = 12'h777;
rom[13411] = 12'h777;
rom[13412] = 12'h777;
rom[13413] = 12'h777;
rom[13414] = 12'h677;
rom[13415] = 12'h676;
rom[13416] = 12'h666;
rom[13417] = 12'h666;
rom[13418] = 12'h666;
rom[13419] = 12'h666;
rom[13420] = 12'h666;
rom[13421] = 12'h666;
rom[13422] = 12'h666;
rom[13423] = 12'h666;
rom[13424] = 12'h666;
rom[13425] = 12'h666;
rom[13426] = 12'h666;
rom[13427] = 12'h666;
rom[13428] = 12'h666;
rom[13429] = 12'h666;
rom[13430] = 12'h666;
rom[13431] = 12'h666;
rom[13432] = 12'h888;
rom[13433] = 12'h888;
rom[13434] = 12'h888;
rom[13435] = 12'h888;
rom[13436] = 12'h777;
rom[13437] = 12'h777;
rom[13438] = 12'h666;
rom[13439] = 12'h666;
rom[13440] = 12'h555;
rom[13441] = 12'h555;
rom[13442] = 12'h444;
rom[13443] = 12'h444;
rom[13444] = 12'h444;
rom[13445] = 12'h444;
rom[13446] = 12'h444;
rom[13447] = 12'h444;
rom[13448] = 12'h444;
rom[13449] = 12'h444;
rom[13450] = 12'h444;
rom[13451] = 12'h444;
rom[13452] = 12'h444;
rom[13453] = 12'h444;
rom[13454] = 12'h444;
rom[13455] = 12'h444;
rom[13456] = 12'h444;
rom[13457] = 12'h444;
rom[13458] = 12'h333;
rom[13459] = 12'h333;
rom[13460] = 12'h222;
rom[13461] = 12'h222;
rom[13462] = 12'h111;
rom[13463] = 12'h111;
rom[13464] = 12'h111;
rom[13465] = 12'h111;
rom[13466] = 12'h  0;
rom[13467] = 12'h  0;
rom[13468] = 12'h  0;
rom[13469] = 12'h  0;
rom[13470] = 12'h  0;
rom[13471] = 12'h  0;
rom[13472] = 12'h  0;
rom[13473] = 12'h  0;
rom[13474] = 12'h  0;
rom[13475] = 12'h  0;
rom[13476] = 12'h  0;
rom[13477] = 12'h  0;
rom[13478] = 12'h  0;
rom[13479] = 12'h  0;
rom[13480] = 12'h  0;
rom[13481] = 12'h  0;
rom[13482] = 12'h  0;
rom[13483] = 12'h  0;
rom[13484] = 12'h  0;
rom[13485] = 12'h  0;
rom[13486] = 12'h  0;
rom[13487] = 12'h  0;
rom[13488] = 12'h  0;
rom[13489] = 12'h  0;
rom[13490] = 12'h  0;
rom[13491] = 12'h  0;
rom[13492] = 12'h  0;
rom[13493] = 12'h  0;
rom[13494] = 12'h  0;
rom[13495] = 12'h  0;
rom[13496] = 12'h  0;
rom[13497] = 12'h  0;
rom[13498] = 12'h111;
rom[13499] = 12'h111;
rom[13500] = 12'h111;
rom[13501] = 12'h  0;
rom[13502] = 12'h  0;
rom[13503] = 12'h  0;
rom[13504] = 12'h  0;
rom[13505] = 12'h  0;
rom[13506] = 12'h  0;
rom[13507] = 12'h  0;
rom[13508] = 12'h  0;
rom[13509] = 12'h111;
rom[13510] = 12'h111;
rom[13511] = 12'h111;
rom[13512] = 12'h111;
rom[13513] = 12'h222;
rom[13514] = 12'h333;
rom[13515] = 12'h444;
rom[13516] = 12'h555;
rom[13517] = 12'h555;
rom[13518] = 12'h555;
rom[13519] = 12'h555;
rom[13520] = 12'h444;
rom[13521] = 12'h333;
rom[13522] = 12'h333;
rom[13523] = 12'h444;
rom[13524] = 12'h444;
rom[13525] = 12'h444;
rom[13526] = 12'h444;
rom[13527] = 12'h444;
rom[13528] = 12'h333;
rom[13529] = 12'h222;
rom[13530] = 12'h111;
rom[13531] = 12'h111;
rom[13532] = 12'h111;
rom[13533] = 12'h  0;
rom[13534] = 12'h  0;
rom[13535] = 12'h  0;
rom[13536] = 12'h  0;
rom[13537] = 12'h  0;
rom[13538] = 12'h  0;
rom[13539] = 12'h  0;
rom[13540] = 12'h  0;
rom[13541] = 12'h  0;
rom[13542] = 12'h  0;
rom[13543] = 12'h  0;
rom[13544] = 12'h  0;
rom[13545] = 12'h  0;
rom[13546] = 12'h111;
rom[13547] = 12'h111;
rom[13548] = 12'h111;
rom[13549] = 12'h222;
rom[13550] = 12'h222;
rom[13551] = 12'h333;
rom[13552] = 12'h444;
rom[13553] = 12'h555;
rom[13554] = 12'h555;
rom[13555] = 12'h666;
rom[13556] = 12'h666;
rom[13557] = 12'h666;
rom[13558] = 12'h555;
rom[13559] = 12'h555;
rom[13560] = 12'h555;
rom[13561] = 12'h555;
rom[13562] = 12'h555;
rom[13563] = 12'h555;
rom[13564] = 12'h555;
rom[13565] = 12'h555;
rom[13566] = 12'h555;
rom[13567] = 12'h555;
rom[13568] = 12'h444;
rom[13569] = 12'h444;
rom[13570] = 12'h444;
rom[13571] = 12'h444;
rom[13572] = 12'h444;
rom[13573] = 12'h444;
rom[13574] = 12'h444;
rom[13575] = 12'h444;
rom[13576] = 12'h444;
rom[13577] = 12'h444;
rom[13578] = 12'h444;
rom[13579] = 12'h444;
rom[13580] = 12'h444;
rom[13581] = 12'h444;
rom[13582] = 12'h444;
rom[13583] = 12'h444;
rom[13584] = 12'h444;
rom[13585] = 12'h555;
rom[13586] = 12'h555;
rom[13587] = 12'h555;
rom[13588] = 12'h555;
rom[13589] = 12'h666;
rom[13590] = 12'h666;
rom[13591] = 12'h777;
rom[13592] = 12'h888;
rom[13593] = 12'h888;
rom[13594] = 12'h999;
rom[13595] = 12'h999;
rom[13596] = 12'haaa;
rom[13597] = 12'haaa;
rom[13598] = 12'haaa;
rom[13599] = 12'haaa;
rom[13600] = 12'h222;
rom[13601] = 12'h222;
rom[13602] = 12'h222;
rom[13603] = 12'h222;
rom[13604] = 12'h111;
rom[13605] = 12'h111;
rom[13606] = 12'h111;
rom[13607] = 12'h111;
rom[13608] = 12'h111;
rom[13609] = 12'h111;
rom[13610] = 12'h111;
rom[13611] = 12'h111;
rom[13612] = 12'h111;
rom[13613] = 12'h111;
rom[13614] = 12'h111;
rom[13615] = 12'h111;
rom[13616] = 12'h111;
rom[13617] = 12'h111;
rom[13618] = 12'h111;
rom[13619] = 12'h222;
rom[13620] = 12'h222;
rom[13621] = 12'h222;
rom[13622] = 12'h222;
rom[13623] = 12'h222;
rom[13624] = 12'h222;
rom[13625] = 12'h222;
rom[13626] = 12'h222;
rom[13627] = 12'h222;
rom[13628] = 12'h222;
rom[13629] = 12'h222;
rom[13630] = 12'h222;
rom[13631] = 12'h222;
rom[13632] = 12'h222;
rom[13633] = 12'h222;
rom[13634] = 12'h222;
rom[13635] = 12'h222;
rom[13636] = 12'h222;
rom[13637] = 12'h333;
rom[13638] = 12'h333;
rom[13639] = 12'h333;
rom[13640] = 12'h333;
rom[13641] = 12'h333;
rom[13642] = 12'h333;
rom[13643] = 12'h333;
rom[13644] = 12'h333;
rom[13645] = 12'h333;
rom[13646] = 12'h333;
rom[13647] = 12'h333;
rom[13648] = 12'h333;
rom[13649] = 12'h333;
rom[13650] = 12'h444;
rom[13651] = 12'h444;
rom[13652] = 12'h444;
rom[13653] = 12'h444;
rom[13654] = 12'h444;
rom[13655] = 12'h444;
rom[13656] = 12'h444;
rom[13657] = 12'h444;
rom[13658] = 12'h444;
rom[13659] = 12'h555;
rom[13660] = 12'h555;
rom[13661] = 12'h555;
rom[13662] = 12'h555;
rom[13663] = 12'h555;
rom[13664] = 12'h666;
rom[13665] = 12'h555;
rom[13666] = 12'h555;
rom[13667] = 12'h555;
rom[13668] = 12'h444;
rom[13669] = 12'h555;
rom[13670] = 12'h555;
rom[13671] = 12'h555;
rom[13672] = 12'h666;
rom[13673] = 12'h777;
rom[13674] = 12'h777;
rom[13675] = 12'h777;
rom[13676] = 12'h666;
rom[13677] = 12'h666;
rom[13678] = 12'h666;
rom[13679] = 12'h555;
rom[13680] = 12'h555;
rom[13681] = 12'h555;
rom[13682] = 12'h444;
rom[13683] = 12'h333;
rom[13684] = 12'h333;
rom[13685] = 12'h333;
rom[13686] = 12'h222;
rom[13687] = 12'h222;
rom[13688] = 12'h222;
rom[13689] = 12'h222;
rom[13690] = 12'h111;
rom[13691] = 12'h111;
rom[13692] = 12'h111;
rom[13693] = 12'h111;
rom[13694] = 12'h111;
rom[13695] = 12'h111;
rom[13696] = 12'h111;
rom[13697] = 12'h111;
rom[13698] = 12'h111;
rom[13699] = 12'h111;
rom[13700] = 12'h100;
rom[13701] = 12'h  0;
rom[13702] = 12'h  0;
rom[13703] = 12'h  0;
rom[13704] = 12'h  0;
rom[13705] = 12'h  0;
rom[13706] = 12'h  0;
rom[13707] = 12'h  0;
rom[13708] = 12'h  0;
rom[13709] = 12'h  0;
rom[13710] = 12'h  0;
rom[13711] = 12'h  0;
rom[13712] = 12'h100;
rom[13713] = 12'h100;
rom[13714] = 12'h200;
rom[13715] = 12'h300;
rom[13716] = 12'h300;
rom[13717] = 12'h400;
rom[13718] = 12'h610;
rom[13719] = 12'h720;
rom[13720] = 12'h820;
rom[13721] = 12'h930;
rom[13722] = 12'h930;
rom[13723] = 12'h931;
rom[13724] = 12'h931;
rom[13725] = 12'h920;
rom[13726] = 12'h810;
rom[13727] = 12'h710;
rom[13728] = 12'h500;
rom[13729] = 12'h500;
rom[13730] = 12'h400;
rom[13731] = 12'h500;
rom[13732] = 12'h500;
rom[13733] = 12'h500;
rom[13734] = 12'h400;
rom[13735] = 12'h400;
rom[13736] = 12'h400;
rom[13737] = 12'h400;
rom[13738] = 12'h400;
rom[13739] = 12'h400;
rom[13740] = 12'h300;
rom[13741] = 12'h300;
rom[13742] = 12'h300;
rom[13743] = 12'h300;
rom[13744] = 12'h200;
rom[13745] = 12'h100;
rom[13746] = 12'h100;
rom[13747] = 12'h100;
rom[13748] = 12'h100;
rom[13749] = 12'h100;
rom[13750] = 12'h100;
rom[13751] = 12'h  0;
rom[13752] = 12'h  0;
rom[13753] = 12'h  0;
rom[13754] = 12'h  0;
rom[13755] = 12'h  0;
rom[13756] = 12'h  0;
rom[13757] = 12'h  0;
rom[13758] = 12'h  0;
rom[13759] = 12'h100;
rom[13760] = 12'h100;
rom[13761] = 12'h100;
rom[13762] = 12'h100;
rom[13763] = 12'h100;
rom[13764] = 12'h100;
rom[13765] = 12'h100;
rom[13766] = 12'h100;
rom[13767] = 12'h100;
rom[13768] = 12'h100;
rom[13769] = 12'h100;
rom[13770] = 12'h200;
rom[13771] = 12'h200;
rom[13772] = 12'h200;
rom[13773] = 12'h200;
rom[13774] = 12'h300;
rom[13775] = 12'h300;
rom[13776] = 12'h300;
rom[13777] = 12'h300;
rom[13778] = 12'h300;
rom[13779] = 12'h400;
rom[13780] = 12'h400;
rom[13781] = 12'h400;
rom[13782] = 12'h400;
rom[13783] = 12'h400;
rom[13784] = 12'h300;
rom[13785] = 12'h300;
rom[13786] = 12'h310;
rom[13787] = 12'h311;
rom[13788] = 12'h321;
rom[13789] = 12'h432;
rom[13790] = 12'h544;
rom[13791] = 12'h555;
rom[13792] = 12'h877;
rom[13793] = 12'h988;
rom[13794] = 12'haaa;
rom[13795] = 12'hcbb;
rom[13796] = 12'hccc;
rom[13797] = 12'hccc;
rom[13798] = 12'hcbb;
rom[13799] = 12'hbbb;
rom[13800] = 12'hbaa;
rom[13801] = 12'hbaa;
rom[13802] = 12'haaa;
rom[13803] = 12'haaa;
rom[13804] = 12'haaa;
rom[13805] = 12'haaa;
rom[13806] = 12'h9aa;
rom[13807] = 12'h899;
rom[13808] = 12'h888;
rom[13809] = 12'h788;
rom[13810] = 12'h777;
rom[13811] = 12'h777;
rom[13812] = 12'h777;
rom[13813] = 12'h777;
rom[13814] = 12'h777;
rom[13815] = 12'h677;
rom[13816] = 12'h777;
rom[13817] = 12'h777;
rom[13818] = 12'h777;
rom[13819] = 12'h777;
rom[13820] = 12'h777;
rom[13821] = 12'h777;
rom[13822] = 12'h777;
rom[13823] = 12'h777;
rom[13824] = 12'h777;
rom[13825] = 12'h777;
rom[13826] = 12'h666;
rom[13827] = 12'h666;
rom[13828] = 12'h666;
rom[13829] = 12'h777;
rom[13830] = 12'h777;
rom[13831] = 12'h888;
rom[13832] = 12'h888;
rom[13833] = 12'h888;
rom[13834] = 12'h888;
rom[13835] = 12'h777;
rom[13836] = 12'h777;
rom[13837] = 12'h666;
rom[13838] = 12'h666;
rom[13839] = 12'h555;
rom[13840] = 12'h555;
rom[13841] = 12'h555;
rom[13842] = 12'h444;
rom[13843] = 12'h555;
rom[13844] = 12'h555;
rom[13845] = 12'h555;
rom[13846] = 12'h444;
rom[13847] = 12'h444;
rom[13848] = 12'h444;
rom[13849] = 12'h555;
rom[13850] = 12'h555;
rom[13851] = 12'h555;
rom[13852] = 12'h555;
rom[13853] = 12'h555;
rom[13854] = 12'h444;
rom[13855] = 12'h444;
rom[13856] = 12'h444;
rom[13857] = 12'h333;
rom[13858] = 12'h333;
rom[13859] = 12'h222;
rom[13860] = 12'h222;
rom[13861] = 12'h222;
rom[13862] = 12'h111;
rom[13863] = 12'h111;
rom[13864] = 12'h111;
rom[13865] = 12'h111;
rom[13866] = 12'h  0;
rom[13867] = 12'h  0;
rom[13868] = 12'h  0;
rom[13869] = 12'h  0;
rom[13870] = 12'h  0;
rom[13871] = 12'h  0;
rom[13872] = 12'h  0;
rom[13873] = 12'h  0;
rom[13874] = 12'h  0;
rom[13875] = 12'h  0;
rom[13876] = 12'h  0;
rom[13877] = 12'h  0;
rom[13878] = 12'h  0;
rom[13879] = 12'h  0;
rom[13880] = 12'h  0;
rom[13881] = 12'h  0;
rom[13882] = 12'h  0;
rom[13883] = 12'h  0;
rom[13884] = 12'h  0;
rom[13885] = 12'h  0;
rom[13886] = 12'h  0;
rom[13887] = 12'h  0;
rom[13888] = 12'h  0;
rom[13889] = 12'h  0;
rom[13890] = 12'h  0;
rom[13891] = 12'h  0;
rom[13892] = 12'h  0;
rom[13893] = 12'h  0;
rom[13894] = 12'h  0;
rom[13895] = 12'h  0;
rom[13896] = 12'h  0;
rom[13897] = 12'h  0;
rom[13898] = 12'h111;
rom[13899] = 12'h111;
rom[13900] = 12'h111;
rom[13901] = 12'h  0;
rom[13902] = 12'h  0;
rom[13903] = 12'h  0;
rom[13904] = 12'h  0;
rom[13905] = 12'h  0;
rom[13906] = 12'h  0;
rom[13907] = 12'h111;
rom[13908] = 12'h111;
rom[13909] = 12'h111;
rom[13910] = 12'h111;
rom[13911] = 12'h111;
rom[13912] = 12'h222;
rom[13913] = 12'h222;
rom[13914] = 12'h444;
rom[13915] = 12'h444;
rom[13916] = 12'h555;
rom[13917] = 12'h555;
rom[13918] = 12'h555;
rom[13919] = 12'h555;
rom[13920] = 12'h444;
rom[13921] = 12'h333;
rom[13922] = 12'h333;
rom[13923] = 12'h444;
rom[13924] = 12'h444;
rom[13925] = 12'h444;
rom[13926] = 12'h444;
rom[13927] = 12'h444;
rom[13928] = 12'h333;
rom[13929] = 12'h222;
rom[13930] = 12'h111;
rom[13931] = 12'h111;
rom[13932] = 12'h111;
rom[13933] = 12'h  0;
rom[13934] = 12'h  0;
rom[13935] = 12'h  0;
rom[13936] = 12'h  0;
rom[13937] = 12'h  0;
rom[13938] = 12'h  0;
rom[13939] = 12'h  0;
rom[13940] = 12'h  0;
rom[13941] = 12'h  0;
rom[13942] = 12'h  0;
rom[13943] = 12'h  0;
rom[13944] = 12'h  0;
rom[13945] = 12'h111;
rom[13946] = 12'h111;
rom[13947] = 12'h111;
rom[13948] = 12'h111;
rom[13949] = 12'h222;
rom[13950] = 12'h333;
rom[13951] = 12'h333;
rom[13952] = 12'h444;
rom[13953] = 12'h555;
rom[13954] = 12'h555;
rom[13955] = 12'h666;
rom[13956] = 12'h666;
rom[13957] = 12'h666;
rom[13958] = 12'h555;
rom[13959] = 12'h555;
rom[13960] = 12'h555;
rom[13961] = 12'h555;
rom[13962] = 12'h555;
rom[13963] = 12'h555;
rom[13964] = 12'h555;
rom[13965] = 12'h555;
rom[13966] = 12'h444;
rom[13967] = 12'h444;
rom[13968] = 12'h444;
rom[13969] = 12'h444;
rom[13970] = 12'h444;
rom[13971] = 12'h444;
rom[13972] = 12'h444;
rom[13973] = 12'h444;
rom[13974] = 12'h444;
rom[13975] = 12'h444;
rom[13976] = 12'h444;
rom[13977] = 12'h444;
rom[13978] = 12'h444;
rom[13979] = 12'h444;
rom[13980] = 12'h444;
rom[13981] = 12'h444;
rom[13982] = 12'h444;
rom[13983] = 12'h444;
rom[13984] = 12'h555;
rom[13985] = 12'h555;
rom[13986] = 12'h555;
rom[13987] = 12'h555;
rom[13988] = 12'h666;
rom[13989] = 12'h666;
rom[13990] = 12'h777;
rom[13991] = 12'h777;
rom[13992] = 12'h888;
rom[13993] = 12'h888;
rom[13994] = 12'h888;
rom[13995] = 12'h999;
rom[13996] = 12'haaa;
rom[13997] = 12'haaa;
rom[13998] = 12'haaa;
rom[13999] = 12'haaa;
rom[14000] = 12'h222;
rom[14001] = 12'h222;
rom[14002] = 12'h222;
rom[14003] = 12'h222;
rom[14004] = 12'h111;
rom[14005] = 12'h111;
rom[14006] = 12'h111;
rom[14007] = 12'h111;
rom[14008] = 12'h111;
rom[14009] = 12'h111;
rom[14010] = 12'h111;
rom[14011] = 12'h111;
rom[14012] = 12'h111;
rom[14013] = 12'h111;
rom[14014] = 12'h111;
rom[14015] = 12'h111;
rom[14016] = 12'h111;
rom[14017] = 12'h111;
rom[14018] = 12'h111;
rom[14019] = 12'h111;
rom[14020] = 12'h222;
rom[14021] = 12'h222;
rom[14022] = 12'h222;
rom[14023] = 12'h222;
rom[14024] = 12'h222;
rom[14025] = 12'h222;
rom[14026] = 12'h222;
rom[14027] = 12'h222;
rom[14028] = 12'h222;
rom[14029] = 12'h222;
rom[14030] = 12'h222;
rom[14031] = 12'h222;
rom[14032] = 12'h222;
rom[14033] = 12'h222;
rom[14034] = 12'h222;
rom[14035] = 12'h222;
rom[14036] = 12'h333;
rom[14037] = 12'h333;
rom[14038] = 12'h333;
rom[14039] = 12'h333;
rom[14040] = 12'h333;
rom[14041] = 12'h333;
rom[14042] = 12'h333;
rom[14043] = 12'h333;
rom[14044] = 12'h333;
rom[14045] = 12'h333;
rom[14046] = 12'h333;
rom[14047] = 12'h444;
rom[14048] = 12'h444;
rom[14049] = 12'h444;
rom[14050] = 12'h444;
rom[14051] = 12'h555;
rom[14052] = 12'h555;
rom[14053] = 12'h555;
rom[14054] = 12'h555;
rom[14055] = 12'h555;
rom[14056] = 12'h555;
rom[14057] = 12'h555;
rom[14058] = 12'h555;
rom[14059] = 12'h555;
rom[14060] = 12'h555;
rom[14061] = 12'h555;
rom[14062] = 12'h555;
rom[14063] = 12'h555;
rom[14064] = 12'h666;
rom[14065] = 12'h666;
rom[14066] = 12'h666;
rom[14067] = 12'h555;
rom[14068] = 12'h555;
rom[14069] = 12'h555;
rom[14070] = 12'h555;
rom[14071] = 12'h555;
rom[14072] = 12'h666;
rom[14073] = 12'h777;
rom[14074] = 12'h777;
rom[14075] = 12'h777;
rom[14076] = 12'h777;
rom[14077] = 12'h666;
rom[14078] = 12'h666;
rom[14079] = 12'h666;
rom[14080] = 12'h666;
rom[14081] = 12'h555;
rom[14082] = 12'h444;
rom[14083] = 12'h444;
rom[14084] = 12'h333;
rom[14085] = 12'h333;
rom[14086] = 12'h222;
rom[14087] = 12'h222;
rom[14088] = 12'h222;
rom[14089] = 12'h222;
rom[14090] = 12'h111;
rom[14091] = 12'h111;
rom[14092] = 12'h111;
rom[14093] = 12'h111;
rom[14094] = 12'h111;
rom[14095] = 12'h111;
rom[14096] = 12'h111;
rom[14097] = 12'h111;
rom[14098] = 12'h100;
rom[14099] = 12'h  0;
rom[14100] = 12'h  0;
rom[14101] = 12'h  0;
rom[14102] = 12'h  0;
rom[14103] = 12'h  0;
rom[14104] = 12'h  0;
rom[14105] = 12'h  0;
rom[14106] = 12'h  0;
rom[14107] = 12'h  0;
rom[14108] = 12'h  0;
rom[14109] = 12'h  0;
rom[14110] = 12'h  0;
rom[14111] = 12'h  0;
rom[14112] = 12'h100;
rom[14113] = 12'h100;
rom[14114] = 12'h100;
rom[14115] = 12'h200;
rom[14116] = 12'h300;
rom[14117] = 12'h400;
rom[14118] = 12'h610;
rom[14119] = 12'h720;
rom[14120] = 12'h820;
rom[14121] = 12'h820;
rom[14122] = 12'h920;
rom[14123] = 12'h931;
rom[14124] = 12'h931;
rom[14125] = 12'h920;
rom[14126] = 12'h820;
rom[14127] = 12'h710;
rom[14128] = 12'h600;
rom[14129] = 12'h500;
rom[14130] = 12'h500;
rom[14131] = 12'h500;
rom[14132] = 12'h500;
rom[14133] = 12'h500;
rom[14134] = 12'h500;
rom[14135] = 12'h400;
rom[14136] = 12'h400;
rom[14137] = 12'h400;
rom[14138] = 12'h400;
rom[14139] = 12'h400;
rom[14140] = 12'h300;
rom[14141] = 12'h300;
rom[14142] = 12'h300;
rom[14143] = 12'h200;
rom[14144] = 12'h100;
rom[14145] = 12'h100;
rom[14146] = 12'h100;
rom[14147] = 12'h100;
rom[14148] = 12'h100;
rom[14149] = 12'h  0;
rom[14150] = 12'h  0;
rom[14151] = 12'h  0;
rom[14152] = 12'h  0;
rom[14153] = 12'h  0;
rom[14154] = 12'h  0;
rom[14155] = 12'h  0;
rom[14156] = 12'h  0;
rom[14157] = 12'h  0;
rom[14158] = 12'h  0;
rom[14159] = 12'h100;
rom[14160] = 12'h100;
rom[14161] = 12'h100;
rom[14162] = 12'h100;
rom[14163] = 12'h100;
rom[14164] = 12'h100;
rom[14165] = 12'h100;
rom[14166] = 12'h100;
rom[14167] = 12'h100;
rom[14168] = 12'h100;
rom[14169] = 12'h100;
rom[14170] = 12'h200;
rom[14171] = 12'h200;
rom[14172] = 12'h200;
rom[14173] = 12'h200;
rom[14174] = 12'h300;
rom[14175] = 12'h300;
rom[14176] = 12'h300;
rom[14177] = 12'h300;
rom[14178] = 12'h300;
rom[14179] = 12'h300;
rom[14180] = 12'h400;
rom[14181] = 12'h400;
rom[14182] = 12'h400;
rom[14183] = 12'h400;
rom[14184] = 12'h300;
rom[14185] = 12'h300;
rom[14186] = 12'h300;
rom[14187] = 12'h210;
rom[14188] = 12'h210;
rom[14189] = 12'h321;
rom[14190] = 12'h432;
rom[14191] = 12'h443;
rom[14192] = 12'h665;
rom[14193] = 12'h777;
rom[14194] = 12'h999;
rom[14195] = 12'hbaa;
rom[14196] = 12'hcbb;
rom[14197] = 12'hccc;
rom[14198] = 12'hcbc;
rom[14199] = 12'hbbb;
rom[14200] = 12'hbbb;
rom[14201] = 12'hbbb;
rom[14202] = 12'hbbb;
rom[14203] = 12'haaa;
rom[14204] = 12'hbbb;
rom[14205] = 12'hbbb;
rom[14206] = 12'haaa;
rom[14207] = 12'h999;
rom[14208] = 12'h888;
rom[14209] = 12'h788;
rom[14210] = 12'h787;
rom[14211] = 12'h777;
rom[14212] = 12'h777;
rom[14213] = 12'h777;
rom[14214] = 12'h777;
rom[14215] = 12'h677;
rom[14216] = 12'h666;
rom[14217] = 12'h777;
rom[14218] = 12'h777;
rom[14219] = 12'h777;
rom[14220] = 12'h777;
rom[14221] = 12'h777;
rom[14222] = 12'h777;
rom[14223] = 12'h766;
rom[14224] = 12'h777;
rom[14225] = 12'h777;
rom[14226] = 12'h666;
rom[14227] = 12'h666;
rom[14228] = 12'h777;
rom[14229] = 12'h888;
rom[14230] = 12'h888;
rom[14231] = 12'h999;
rom[14232] = 12'h888;
rom[14233] = 12'h777;
rom[14234] = 12'h777;
rom[14235] = 12'h666;
rom[14236] = 12'h666;
rom[14237] = 12'h666;
rom[14238] = 12'h555;
rom[14239] = 12'h555;
rom[14240] = 12'h555;
rom[14241] = 12'h555;
rom[14242] = 12'h555;
rom[14243] = 12'h555;
rom[14244] = 12'h555;
rom[14245] = 12'h555;
rom[14246] = 12'h555;
rom[14247] = 12'h555;
rom[14248] = 12'h555;
rom[14249] = 12'h555;
rom[14250] = 12'h555;
rom[14251] = 12'h666;
rom[14252] = 12'h555;
rom[14253] = 12'h555;
rom[14254] = 12'h444;
rom[14255] = 12'h444;
rom[14256] = 12'h333;
rom[14257] = 12'h333;
rom[14258] = 12'h333;
rom[14259] = 12'h222;
rom[14260] = 12'h222;
rom[14261] = 12'h222;
rom[14262] = 12'h111;
rom[14263] = 12'h111;
rom[14264] = 12'h111;
rom[14265] = 12'h111;
rom[14266] = 12'h  0;
rom[14267] = 12'h  0;
rom[14268] = 12'h  0;
rom[14269] = 12'h  0;
rom[14270] = 12'h  0;
rom[14271] = 12'h  0;
rom[14272] = 12'h  0;
rom[14273] = 12'h  0;
rom[14274] = 12'h  0;
rom[14275] = 12'h  0;
rom[14276] = 12'h  0;
rom[14277] = 12'h  0;
rom[14278] = 12'h  0;
rom[14279] = 12'h  0;
rom[14280] = 12'h  0;
rom[14281] = 12'h  0;
rom[14282] = 12'h  0;
rom[14283] = 12'h  0;
rom[14284] = 12'h  0;
rom[14285] = 12'h  0;
rom[14286] = 12'h  0;
rom[14287] = 12'h  0;
rom[14288] = 12'h  0;
rom[14289] = 12'h  0;
rom[14290] = 12'h  0;
rom[14291] = 12'h  0;
rom[14292] = 12'h  0;
rom[14293] = 12'h  0;
rom[14294] = 12'h  0;
rom[14295] = 12'h  0;
rom[14296] = 12'h  0;
rom[14297] = 12'h  0;
rom[14298] = 12'h111;
rom[14299] = 12'h111;
rom[14300] = 12'h111;
rom[14301] = 12'h  0;
rom[14302] = 12'h  0;
rom[14303] = 12'h  0;
rom[14304] = 12'h  0;
rom[14305] = 12'h  0;
rom[14306] = 12'h  0;
rom[14307] = 12'h111;
rom[14308] = 12'h111;
rom[14309] = 12'h111;
rom[14310] = 12'h111;
rom[14311] = 12'h111;
rom[14312] = 12'h222;
rom[14313] = 12'h333;
rom[14314] = 12'h444;
rom[14315] = 12'h555;
rom[14316] = 12'h555;
rom[14317] = 12'h555;
rom[14318] = 12'h555;
rom[14319] = 12'h555;
rom[14320] = 12'h333;
rom[14321] = 12'h333;
rom[14322] = 12'h333;
rom[14323] = 12'h444;
rom[14324] = 12'h444;
rom[14325] = 12'h444;
rom[14326] = 12'h444;
rom[14327] = 12'h444;
rom[14328] = 12'h333;
rom[14329] = 12'h222;
rom[14330] = 12'h111;
rom[14331] = 12'h111;
rom[14332] = 12'h111;
rom[14333] = 12'h  0;
rom[14334] = 12'h  0;
rom[14335] = 12'h  0;
rom[14336] = 12'h  0;
rom[14337] = 12'h  0;
rom[14338] = 12'h  0;
rom[14339] = 12'h  0;
rom[14340] = 12'h  0;
rom[14341] = 12'h  0;
rom[14342] = 12'h  0;
rom[14343] = 12'h  0;
rom[14344] = 12'h  0;
rom[14345] = 12'h  0;
rom[14346] = 12'h111;
rom[14347] = 12'h111;
rom[14348] = 12'h111;
rom[14349] = 12'h222;
rom[14350] = 12'h333;
rom[14351] = 12'h444;
rom[14352] = 12'h555;
rom[14353] = 12'h555;
rom[14354] = 12'h555;
rom[14355] = 12'h666;
rom[14356] = 12'h666;
rom[14357] = 12'h555;
rom[14358] = 12'h555;
rom[14359] = 12'h555;
rom[14360] = 12'h555;
rom[14361] = 12'h555;
rom[14362] = 12'h555;
rom[14363] = 12'h555;
rom[14364] = 12'h555;
rom[14365] = 12'h555;
rom[14366] = 12'h555;
rom[14367] = 12'h444;
rom[14368] = 12'h444;
rom[14369] = 12'h555;
rom[14370] = 12'h555;
rom[14371] = 12'h555;
rom[14372] = 12'h555;
rom[14373] = 12'h444;
rom[14374] = 12'h444;
rom[14375] = 12'h444;
rom[14376] = 12'h444;
rom[14377] = 12'h444;
rom[14378] = 12'h444;
rom[14379] = 12'h444;
rom[14380] = 12'h444;
rom[14381] = 12'h444;
rom[14382] = 12'h444;
rom[14383] = 12'h444;
rom[14384] = 12'h555;
rom[14385] = 12'h555;
rom[14386] = 12'h555;
rom[14387] = 12'h555;
rom[14388] = 12'h666;
rom[14389] = 12'h666;
rom[14390] = 12'h777;
rom[14391] = 12'h777;
rom[14392] = 12'h777;
rom[14393] = 12'h888;
rom[14394] = 12'h888;
rom[14395] = 12'h999;
rom[14396] = 12'h999;
rom[14397] = 12'haaa;
rom[14398] = 12'haaa;
rom[14399] = 12'haaa;
rom[14400] = 12'h222;
rom[14401] = 12'h222;
rom[14402] = 12'h222;
rom[14403] = 12'h222;
rom[14404] = 12'h111;
rom[14405] = 12'h111;
rom[14406] = 12'h111;
rom[14407] = 12'h111;
rom[14408] = 12'h111;
rom[14409] = 12'h111;
rom[14410] = 12'h111;
rom[14411] = 12'h111;
rom[14412] = 12'h111;
rom[14413] = 12'h111;
rom[14414] = 12'h111;
rom[14415] = 12'h111;
rom[14416] = 12'h111;
rom[14417] = 12'h111;
rom[14418] = 12'h111;
rom[14419] = 12'h111;
rom[14420] = 12'h222;
rom[14421] = 12'h222;
rom[14422] = 12'h222;
rom[14423] = 12'h222;
rom[14424] = 12'h333;
rom[14425] = 12'h222;
rom[14426] = 12'h222;
rom[14427] = 12'h222;
rom[14428] = 12'h222;
rom[14429] = 12'h222;
rom[14430] = 12'h222;
rom[14431] = 12'h222;
rom[14432] = 12'h222;
rom[14433] = 12'h222;
rom[14434] = 12'h222;
rom[14435] = 12'h333;
rom[14436] = 12'h333;
rom[14437] = 12'h333;
rom[14438] = 12'h333;
rom[14439] = 12'h333;
rom[14440] = 12'h333;
rom[14441] = 12'h333;
rom[14442] = 12'h333;
rom[14443] = 12'h333;
rom[14444] = 12'h333;
rom[14445] = 12'h444;
rom[14446] = 12'h444;
rom[14447] = 12'h444;
rom[14448] = 12'h444;
rom[14449] = 12'h444;
rom[14450] = 12'h555;
rom[14451] = 12'h555;
rom[14452] = 12'h555;
rom[14453] = 12'h555;
rom[14454] = 12'h555;
rom[14455] = 12'h555;
rom[14456] = 12'h555;
rom[14457] = 12'h555;
rom[14458] = 12'h555;
rom[14459] = 12'h555;
rom[14460] = 12'h555;
rom[14461] = 12'h555;
rom[14462] = 12'h555;
rom[14463] = 12'h555;
rom[14464] = 12'h666;
rom[14465] = 12'h666;
rom[14466] = 12'h666;
rom[14467] = 12'h666;
rom[14468] = 12'h666;
rom[14469] = 12'h555;
rom[14470] = 12'h555;
rom[14471] = 12'h555;
rom[14472] = 12'h666;
rom[14473] = 12'h666;
rom[14474] = 12'h777;
rom[14475] = 12'h777;
rom[14476] = 12'h777;
rom[14477] = 12'h666;
rom[14478] = 12'h666;
rom[14479] = 12'h666;
rom[14480] = 12'h666;
rom[14481] = 12'h555;
rom[14482] = 12'h444;
rom[14483] = 12'h444;
rom[14484] = 12'h444;
rom[14485] = 12'h333;
rom[14486] = 12'h333;
rom[14487] = 12'h222;
rom[14488] = 12'h222;
rom[14489] = 12'h222;
rom[14490] = 12'h222;
rom[14491] = 12'h111;
rom[14492] = 12'h111;
rom[14493] = 12'h111;
rom[14494] = 12'h111;
rom[14495] = 12'h111;
rom[14496] = 12'h111;
rom[14497] = 12'h100;
rom[14498] = 12'h  0;
rom[14499] = 12'h  0;
rom[14500] = 12'h  0;
rom[14501] = 12'h  0;
rom[14502] = 12'h  0;
rom[14503] = 12'h  0;
rom[14504] = 12'h  0;
rom[14505] = 12'h  0;
rom[14506] = 12'h  0;
rom[14507] = 12'h  0;
rom[14508] = 12'h  0;
rom[14509] = 12'h  0;
rom[14510] = 12'h  0;
rom[14511] = 12'h  0;
rom[14512] = 12'h  0;
rom[14513] = 12'h100;
rom[14514] = 12'h100;
rom[14515] = 12'h200;
rom[14516] = 12'h300;
rom[14517] = 12'h400;
rom[14518] = 12'h510;
rom[14519] = 12'h710;
rom[14520] = 12'h820;
rom[14521] = 12'h820;
rom[14522] = 12'h920;
rom[14523] = 12'h921;
rom[14524] = 12'h931;
rom[14525] = 12'h921;
rom[14526] = 12'h820;
rom[14527] = 12'h710;
rom[14528] = 12'h610;
rom[14529] = 12'h500;
rom[14530] = 12'h500;
rom[14531] = 12'h500;
rom[14532] = 12'h500;
rom[14533] = 12'h500;
rom[14534] = 12'h500;
rom[14535] = 12'h400;
rom[14536] = 12'h400;
rom[14537] = 12'h400;
rom[14538] = 12'h400;
rom[14539] = 12'h300;
rom[14540] = 12'h300;
rom[14541] = 12'h300;
rom[14542] = 12'h200;
rom[14543] = 12'h200;
rom[14544] = 12'h100;
rom[14545] = 12'h100;
rom[14546] = 12'h100;
rom[14547] = 12'h  0;
rom[14548] = 12'h  0;
rom[14549] = 12'h  0;
rom[14550] = 12'h  0;
rom[14551] = 12'h  0;
rom[14552] = 12'h  0;
rom[14553] = 12'h  0;
rom[14554] = 12'h  0;
rom[14555] = 12'h  0;
rom[14556] = 12'h  0;
rom[14557] = 12'h  0;
rom[14558] = 12'h  0;
rom[14559] = 12'h100;
rom[14560] = 12'h100;
rom[14561] = 12'h100;
rom[14562] = 12'h100;
rom[14563] = 12'h100;
rom[14564] = 12'h100;
rom[14565] = 12'h100;
rom[14566] = 12'h100;
rom[14567] = 12'h100;
rom[14568] = 12'h100;
rom[14569] = 12'h100;
rom[14570] = 12'h200;
rom[14571] = 12'h200;
rom[14572] = 12'h200;
rom[14573] = 12'h200;
rom[14574] = 12'h200;
rom[14575] = 12'h300;
rom[14576] = 12'h300;
rom[14577] = 12'h300;
rom[14578] = 12'h300;
rom[14579] = 12'h300;
rom[14580] = 12'h300;
rom[14581] = 12'h300;
rom[14582] = 12'h300;
rom[14583] = 12'h300;
rom[14584] = 12'h300;
rom[14585] = 12'h300;
rom[14586] = 12'h300;
rom[14587] = 12'h200;
rom[14588] = 12'h200;
rom[14589] = 12'h210;
rom[14590] = 12'h321;
rom[14591] = 12'h422;
rom[14592] = 12'h544;
rom[14593] = 12'h655;
rom[14594] = 12'h777;
rom[14595] = 12'h999;
rom[14596] = 12'hbab;
rom[14597] = 12'hcbb;
rom[14598] = 12'hccc;
rom[14599] = 12'hccc;
rom[14600] = 12'hbbb;
rom[14601] = 12'hbbb;
rom[14602] = 12'hbbb;
rom[14603] = 12'hbbb;
rom[14604] = 12'hbbb;
rom[14605] = 12'hbbb;
rom[14606] = 12'haaa;
rom[14607] = 12'h999;
rom[14608] = 12'h888;
rom[14609] = 12'h888;
rom[14610] = 12'h788;
rom[14611] = 12'h777;
rom[14612] = 12'h777;
rom[14613] = 12'h777;
rom[14614] = 12'h777;
rom[14615] = 12'h777;
rom[14616] = 12'h666;
rom[14617] = 12'h666;
rom[14618] = 12'h777;
rom[14619] = 12'h777;
rom[14620] = 12'h777;
rom[14621] = 12'h777;
rom[14622] = 12'h777;
rom[14623] = 12'h766;
rom[14624] = 12'h777;
rom[14625] = 12'h777;
rom[14626] = 12'h777;
rom[14627] = 12'h777;
rom[14628] = 12'h888;
rom[14629] = 12'h888;
rom[14630] = 12'h888;
rom[14631] = 12'h888;
rom[14632] = 12'h777;
rom[14633] = 12'h666;
rom[14634] = 12'h666;
rom[14635] = 12'h666;
rom[14636] = 12'h666;
rom[14637] = 12'h666;
rom[14638] = 12'h666;
rom[14639] = 12'h555;
rom[14640] = 12'h666;
rom[14641] = 12'h555;
rom[14642] = 12'h555;
rom[14643] = 12'h555;
rom[14644] = 12'h555;
rom[14645] = 12'h555;
rom[14646] = 12'h555;
rom[14647] = 12'h555;
rom[14648] = 12'h555;
rom[14649] = 12'h555;
rom[14650] = 12'h555;
rom[14651] = 12'h555;
rom[14652] = 12'h555;
rom[14653] = 12'h555;
rom[14654] = 12'h444;
rom[14655] = 12'h444;
rom[14656] = 12'h333;
rom[14657] = 12'h333;
rom[14658] = 12'h222;
rom[14659] = 12'h222;
rom[14660] = 12'h222;
rom[14661] = 12'h111;
rom[14662] = 12'h111;
rom[14663] = 12'h111;
rom[14664] = 12'h111;
rom[14665] = 12'h111;
rom[14666] = 12'h  0;
rom[14667] = 12'h  0;
rom[14668] = 12'h  0;
rom[14669] = 12'h  0;
rom[14670] = 12'h  0;
rom[14671] = 12'h  0;
rom[14672] = 12'h  0;
rom[14673] = 12'h  0;
rom[14674] = 12'h  0;
rom[14675] = 12'h  0;
rom[14676] = 12'h  0;
rom[14677] = 12'h  0;
rom[14678] = 12'h  0;
rom[14679] = 12'h  0;
rom[14680] = 12'h  0;
rom[14681] = 12'h  0;
rom[14682] = 12'h  0;
rom[14683] = 12'h  0;
rom[14684] = 12'h  0;
rom[14685] = 12'h  0;
rom[14686] = 12'h  0;
rom[14687] = 12'h  0;
rom[14688] = 12'h  0;
rom[14689] = 12'h  0;
rom[14690] = 12'h  0;
rom[14691] = 12'h  0;
rom[14692] = 12'h  0;
rom[14693] = 12'h  0;
rom[14694] = 12'h  0;
rom[14695] = 12'h  0;
rom[14696] = 12'h  0;
rom[14697] = 12'h  0;
rom[14698] = 12'h111;
rom[14699] = 12'h111;
rom[14700] = 12'h111;
rom[14701] = 12'h  0;
rom[14702] = 12'h  0;
rom[14703] = 12'h  0;
rom[14704] = 12'h  0;
rom[14705] = 12'h  0;
rom[14706] = 12'h  0;
rom[14707] = 12'h111;
rom[14708] = 12'h111;
rom[14709] = 12'h111;
rom[14710] = 12'h111;
rom[14711] = 12'h222;
rom[14712] = 12'h333;
rom[14713] = 12'h333;
rom[14714] = 12'h444;
rom[14715] = 12'h555;
rom[14716] = 12'h555;
rom[14717] = 12'h444;
rom[14718] = 12'h444;
rom[14719] = 12'h444;
rom[14720] = 12'h333;
rom[14721] = 12'h333;
rom[14722] = 12'h444;
rom[14723] = 12'h444;
rom[14724] = 12'h444;
rom[14725] = 12'h444;
rom[14726] = 12'h444;
rom[14727] = 12'h444;
rom[14728] = 12'h333;
rom[14729] = 12'h222;
rom[14730] = 12'h111;
rom[14731] = 12'h111;
rom[14732] = 12'h111;
rom[14733] = 12'h  0;
rom[14734] = 12'h  0;
rom[14735] = 12'h  0;
rom[14736] = 12'h  0;
rom[14737] = 12'h  0;
rom[14738] = 12'h  0;
rom[14739] = 12'h  0;
rom[14740] = 12'h  0;
rom[14741] = 12'h  0;
rom[14742] = 12'h  0;
rom[14743] = 12'h  0;
rom[14744] = 12'h  0;
rom[14745] = 12'h  0;
rom[14746] = 12'h111;
rom[14747] = 12'h111;
rom[14748] = 12'h111;
rom[14749] = 12'h222;
rom[14750] = 12'h333;
rom[14751] = 12'h444;
rom[14752] = 12'h555;
rom[14753] = 12'h555;
rom[14754] = 12'h666;
rom[14755] = 12'h666;
rom[14756] = 12'h666;
rom[14757] = 12'h555;
rom[14758] = 12'h555;
rom[14759] = 12'h555;
rom[14760] = 12'h555;
rom[14761] = 12'h555;
rom[14762] = 12'h555;
rom[14763] = 12'h555;
rom[14764] = 12'h555;
rom[14765] = 12'h555;
rom[14766] = 12'h555;
rom[14767] = 12'h555;
rom[14768] = 12'h555;
rom[14769] = 12'h555;
rom[14770] = 12'h555;
rom[14771] = 12'h555;
rom[14772] = 12'h555;
rom[14773] = 12'h444;
rom[14774] = 12'h444;
rom[14775] = 12'h444;
rom[14776] = 12'h444;
rom[14777] = 12'h444;
rom[14778] = 12'h444;
rom[14779] = 12'h444;
rom[14780] = 12'h444;
rom[14781] = 12'h444;
rom[14782] = 12'h444;
rom[14783] = 12'h555;
rom[14784] = 12'h555;
rom[14785] = 12'h555;
rom[14786] = 12'h555;
rom[14787] = 12'h666;
rom[14788] = 12'h666;
rom[14789] = 12'h666;
rom[14790] = 12'h777;
rom[14791] = 12'h777;
rom[14792] = 12'h777;
rom[14793] = 12'h888;
rom[14794] = 12'h888;
rom[14795] = 12'h999;
rom[14796] = 12'h999;
rom[14797] = 12'haaa;
rom[14798] = 12'haaa;
rom[14799] = 12'haaa;
rom[14800] = 12'h222;
rom[14801] = 12'h222;
rom[14802] = 12'h222;
rom[14803] = 12'h222;
rom[14804] = 12'h222;
rom[14805] = 12'h222;
rom[14806] = 12'h222;
rom[14807] = 12'h222;
rom[14808] = 12'h222;
rom[14809] = 12'h111;
rom[14810] = 12'h111;
rom[14811] = 12'h111;
rom[14812] = 12'h111;
rom[14813] = 12'h111;
rom[14814] = 12'h111;
rom[14815] = 12'h111;
rom[14816] = 12'h111;
rom[14817] = 12'h111;
rom[14818] = 12'h111;
rom[14819] = 12'h111;
rom[14820] = 12'h222;
rom[14821] = 12'h222;
rom[14822] = 12'h222;
rom[14823] = 12'h222;
rom[14824] = 12'h333;
rom[14825] = 12'h333;
rom[14826] = 12'h333;
rom[14827] = 12'h222;
rom[14828] = 12'h222;
rom[14829] = 12'h222;
rom[14830] = 12'h333;
rom[14831] = 12'h333;
rom[14832] = 12'h333;
rom[14833] = 12'h333;
rom[14834] = 12'h333;
rom[14835] = 12'h333;
rom[14836] = 12'h333;
rom[14837] = 12'h333;
rom[14838] = 12'h333;
rom[14839] = 12'h333;
rom[14840] = 12'h444;
rom[14841] = 12'h444;
rom[14842] = 12'h444;
rom[14843] = 12'h444;
rom[14844] = 12'h444;
rom[14845] = 12'h444;
rom[14846] = 12'h555;
rom[14847] = 12'h555;
rom[14848] = 12'h555;
rom[14849] = 12'h555;
rom[14850] = 12'h555;
rom[14851] = 12'h555;
rom[14852] = 12'h555;
rom[14853] = 12'h555;
rom[14854] = 12'h555;
rom[14855] = 12'h555;
rom[14856] = 12'h555;
rom[14857] = 12'h555;
rom[14858] = 12'h555;
rom[14859] = 12'h555;
rom[14860] = 12'h555;
rom[14861] = 12'h555;
rom[14862] = 12'h555;
rom[14863] = 12'h555;
rom[14864] = 12'h555;
rom[14865] = 12'h555;
rom[14866] = 12'h666;
rom[14867] = 12'h666;
rom[14868] = 12'h666;
rom[14869] = 12'h666;
rom[14870] = 12'h666;
rom[14871] = 12'h555;
rom[14872] = 12'h666;
rom[14873] = 12'h666;
rom[14874] = 12'h777;
rom[14875] = 12'h777;
rom[14876] = 12'h777;
rom[14877] = 12'h666;
rom[14878] = 12'h666;
rom[14879] = 12'h666;
rom[14880] = 12'h666;
rom[14881] = 12'h555;
rom[14882] = 12'h555;
rom[14883] = 12'h444;
rom[14884] = 12'h444;
rom[14885] = 12'h333;
rom[14886] = 12'h333;
rom[14887] = 12'h333;
rom[14888] = 12'h222;
rom[14889] = 12'h222;
rom[14890] = 12'h222;
rom[14891] = 12'h111;
rom[14892] = 12'h111;
rom[14893] = 12'h111;
rom[14894] = 12'h111;
rom[14895] = 12'h111;
rom[14896] = 12'h111;
rom[14897] = 12'h100;
rom[14898] = 12'h  0;
rom[14899] = 12'h  0;
rom[14900] = 12'h  0;
rom[14901] = 12'h  0;
rom[14902] = 12'h  0;
rom[14903] = 12'h  0;
rom[14904] = 12'h  0;
rom[14905] = 12'h  0;
rom[14906] = 12'h  0;
rom[14907] = 12'h  0;
rom[14908] = 12'h  0;
rom[14909] = 12'h  0;
rom[14910] = 12'h  0;
rom[14911] = 12'h  0;
rom[14912] = 12'h  0;
rom[14913] = 12'h100;
rom[14914] = 12'h100;
rom[14915] = 12'h200;
rom[14916] = 12'h300;
rom[14917] = 12'h400;
rom[14918] = 12'h510;
rom[14919] = 12'h710;
rom[14920] = 12'h820;
rom[14921] = 12'h820;
rom[14922] = 12'h920;
rom[14923] = 12'h920;
rom[14924] = 12'h931;
rom[14925] = 12'h921;
rom[14926] = 12'h820;
rom[14927] = 12'h710;
rom[14928] = 12'h610;
rom[14929] = 12'h500;
rom[14930] = 12'h500;
rom[14931] = 12'h500;
rom[14932] = 12'h500;
rom[14933] = 12'h500;
rom[14934] = 12'h500;
rom[14935] = 12'h400;
rom[14936] = 12'h400;
rom[14937] = 12'h400;
rom[14938] = 12'h400;
rom[14939] = 12'h300;
rom[14940] = 12'h300;
rom[14941] = 12'h300;
rom[14942] = 12'h200;
rom[14943] = 12'h200;
rom[14944] = 12'h100;
rom[14945] = 12'h  0;
rom[14946] = 12'h  0;
rom[14947] = 12'h  0;
rom[14948] = 12'h  0;
rom[14949] = 12'h  0;
rom[14950] = 12'h  0;
rom[14951] = 12'h  0;
rom[14952] = 12'h  0;
rom[14953] = 12'h  0;
rom[14954] = 12'h  0;
rom[14955] = 12'h  0;
rom[14956] = 12'h  0;
rom[14957] = 12'h  0;
rom[14958] = 12'h  0;
rom[14959] = 12'h  0;
rom[14960] = 12'h100;
rom[14961] = 12'h100;
rom[14962] = 12'h100;
rom[14963] = 12'h100;
rom[14964] = 12'h100;
rom[14965] = 12'h100;
rom[14966] = 12'h100;
rom[14967] = 12'h100;
rom[14968] = 12'h100;
rom[14969] = 12'h100;
rom[14970] = 12'h100;
rom[14971] = 12'h200;
rom[14972] = 12'h200;
rom[14973] = 12'h200;
rom[14974] = 12'h200;
rom[14975] = 12'h200;
rom[14976] = 12'h200;
rom[14977] = 12'h300;
rom[14978] = 12'h300;
rom[14979] = 12'h300;
rom[14980] = 12'h300;
rom[14981] = 12'h300;
rom[14982] = 12'h300;
rom[14983] = 12'h300;
rom[14984] = 12'h300;
rom[14985] = 12'h300;
rom[14986] = 12'h300;
rom[14987] = 12'h300;
rom[14988] = 12'h300;
rom[14989] = 12'h310;
rom[14990] = 12'h311;
rom[14991] = 12'h321;
rom[14992] = 12'h433;
rom[14993] = 12'h444;
rom[14994] = 12'h666;
rom[14995] = 12'h888;
rom[14996] = 12'ha99;
rom[14997] = 12'hbbb;
rom[14998] = 12'hcbb;
rom[14999] = 12'hccc;
rom[15000] = 12'hbbb;
rom[15001] = 12'hbbb;
rom[15002] = 12'hbbb;
rom[15003] = 12'hbbb;
rom[15004] = 12'hbbb;
rom[15005] = 12'hbbb;
rom[15006] = 12'haaa;
rom[15007] = 12'h999;
rom[15008] = 12'h888;
rom[15009] = 12'h888;
rom[15010] = 12'h788;
rom[15011] = 12'h788;
rom[15012] = 12'h777;
rom[15013] = 12'h777;
rom[15014] = 12'h777;
rom[15015] = 12'h777;
rom[15016] = 12'h777;
rom[15017] = 12'h777;
rom[15018] = 12'h777;
rom[15019] = 12'h777;
rom[15020] = 12'h777;
rom[15021] = 12'h777;
rom[15022] = 12'h777;
rom[15023] = 12'h777;
rom[15024] = 12'h777;
rom[15025] = 12'h777;
rom[15026] = 12'h888;
rom[15027] = 12'h999;
rom[15028] = 12'h999;
rom[15029] = 12'h888;
rom[15030] = 12'h777;
rom[15031] = 12'h777;
rom[15032] = 12'h666;
rom[15033] = 12'h666;
rom[15034] = 12'h666;
rom[15035] = 12'h666;
rom[15036] = 12'h666;
rom[15037] = 12'h666;
rom[15038] = 12'h666;
rom[15039] = 12'h666;
rom[15040] = 12'h666;
rom[15041] = 12'h666;
rom[15042] = 12'h666;
rom[15043] = 12'h555;
rom[15044] = 12'h555;
rom[15045] = 12'h555;
rom[15046] = 12'h555;
rom[15047] = 12'h666;
rom[15048] = 12'h555;
rom[15049] = 12'h555;
rom[15050] = 12'h555;
rom[15051] = 12'h555;
rom[15052] = 12'h555;
rom[15053] = 12'h444;
rom[15054] = 12'h444;
rom[15055] = 12'h333;
rom[15056] = 12'h333;
rom[15057] = 12'h222;
rom[15058] = 12'h222;
rom[15059] = 12'h222;
rom[15060] = 12'h111;
rom[15061] = 12'h111;
rom[15062] = 12'h111;
rom[15063] = 12'h111;
rom[15064] = 12'h111;
rom[15065] = 12'h111;
rom[15066] = 12'h  0;
rom[15067] = 12'h  0;
rom[15068] = 12'h  0;
rom[15069] = 12'h  0;
rom[15070] = 12'h  0;
rom[15071] = 12'h  0;
rom[15072] = 12'h  0;
rom[15073] = 12'h  0;
rom[15074] = 12'h  0;
rom[15075] = 12'h  0;
rom[15076] = 12'h  0;
rom[15077] = 12'h  0;
rom[15078] = 12'h  0;
rom[15079] = 12'h  0;
rom[15080] = 12'h  0;
rom[15081] = 12'h  0;
rom[15082] = 12'h  0;
rom[15083] = 12'h  0;
rom[15084] = 12'h  0;
rom[15085] = 12'h  0;
rom[15086] = 12'h  0;
rom[15087] = 12'h  0;
rom[15088] = 12'h  0;
rom[15089] = 12'h  0;
rom[15090] = 12'h  0;
rom[15091] = 12'h  0;
rom[15092] = 12'h  0;
rom[15093] = 12'h  0;
rom[15094] = 12'h  0;
rom[15095] = 12'h  0;
rom[15096] = 12'h  0;
rom[15097] = 12'h  0;
rom[15098] = 12'h111;
rom[15099] = 12'h111;
rom[15100] = 12'h111;
rom[15101] = 12'h  0;
rom[15102] = 12'h  0;
rom[15103] = 12'h  0;
rom[15104] = 12'h  0;
rom[15105] = 12'h  0;
rom[15106] = 12'h  0;
rom[15107] = 12'h111;
rom[15108] = 12'h111;
rom[15109] = 12'h111;
rom[15110] = 12'h111;
rom[15111] = 12'h222;
rom[15112] = 12'h333;
rom[15113] = 12'h444;
rom[15114] = 12'h444;
rom[15115] = 12'h444;
rom[15116] = 12'h444;
rom[15117] = 12'h444;
rom[15118] = 12'h444;
rom[15119] = 12'h444;
rom[15120] = 12'h333;
rom[15121] = 12'h333;
rom[15122] = 12'h444;
rom[15123] = 12'h444;
rom[15124] = 12'h444;
rom[15125] = 12'h333;
rom[15126] = 12'h333;
rom[15127] = 12'h444;
rom[15128] = 12'h333;
rom[15129] = 12'h222;
rom[15130] = 12'h111;
rom[15131] = 12'h111;
rom[15132] = 12'h111;
rom[15133] = 12'h  0;
rom[15134] = 12'h  0;
rom[15135] = 12'h  0;
rom[15136] = 12'h  0;
rom[15137] = 12'h  0;
rom[15138] = 12'h  0;
rom[15139] = 12'h  0;
rom[15140] = 12'h  0;
rom[15141] = 12'h  0;
rom[15142] = 12'h  0;
rom[15143] = 12'h  0;
rom[15144] = 12'h  0;
rom[15145] = 12'h  0;
rom[15146] = 12'h111;
rom[15147] = 12'h111;
rom[15148] = 12'h111;
rom[15149] = 12'h222;
rom[15150] = 12'h444;
rom[15151] = 12'h444;
rom[15152] = 12'h666;
rom[15153] = 12'h666;
rom[15154] = 12'h666;
rom[15155] = 12'h666;
rom[15156] = 12'h666;
rom[15157] = 12'h555;
rom[15158] = 12'h555;
rom[15159] = 12'h555;
rom[15160] = 12'h555;
rom[15161] = 12'h555;
rom[15162] = 12'h555;
rom[15163] = 12'h555;
rom[15164] = 12'h555;
rom[15165] = 12'h555;
rom[15166] = 12'h555;
rom[15167] = 12'h555;
rom[15168] = 12'h555;
rom[15169] = 12'h555;
rom[15170] = 12'h555;
rom[15171] = 12'h555;
rom[15172] = 12'h555;
rom[15173] = 12'h555;
rom[15174] = 12'h444;
rom[15175] = 12'h444;
rom[15176] = 12'h444;
rom[15177] = 12'h444;
rom[15178] = 12'h444;
rom[15179] = 12'h444;
rom[15180] = 12'h555;
rom[15181] = 12'h555;
rom[15182] = 12'h555;
rom[15183] = 12'h555;
rom[15184] = 12'h555;
rom[15185] = 12'h555;
rom[15186] = 12'h666;
rom[15187] = 12'h666;
rom[15188] = 12'h666;
rom[15189] = 12'h777;
rom[15190] = 12'h777;
rom[15191] = 12'h777;
rom[15192] = 12'h777;
rom[15193] = 12'h888;
rom[15194] = 12'h888;
rom[15195] = 12'h999;
rom[15196] = 12'haaa;
rom[15197] = 12'haaa;
rom[15198] = 12'haaa;
rom[15199] = 12'haaa;
rom[15200] = 12'h222;
rom[15201] = 12'h222;
rom[15202] = 12'h222;
rom[15203] = 12'h222;
rom[15204] = 12'h222;
rom[15205] = 12'h222;
rom[15206] = 12'h222;
rom[15207] = 12'h222;
rom[15208] = 12'h222;
rom[15209] = 12'h222;
rom[15210] = 12'h111;
rom[15211] = 12'h111;
rom[15212] = 12'h111;
rom[15213] = 12'h111;
rom[15214] = 12'h111;
rom[15215] = 12'h111;
rom[15216] = 12'h222;
rom[15217] = 12'h222;
rom[15218] = 12'h222;
rom[15219] = 12'h222;
rom[15220] = 12'h222;
rom[15221] = 12'h222;
rom[15222] = 12'h222;
rom[15223] = 12'h222;
rom[15224] = 12'h333;
rom[15225] = 12'h333;
rom[15226] = 12'h333;
rom[15227] = 12'h333;
rom[15228] = 12'h333;
rom[15229] = 12'h333;
rom[15230] = 12'h333;
rom[15231] = 12'h333;
rom[15232] = 12'h333;
rom[15233] = 12'h333;
rom[15234] = 12'h333;
rom[15235] = 12'h444;
rom[15236] = 12'h444;
rom[15237] = 12'h444;
rom[15238] = 12'h444;
rom[15239] = 12'h444;
rom[15240] = 12'h444;
rom[15241] = 12'h444;
rom[15242] = 12'h555;
rom[15243] = 12'h555;
rom[15244] = 12'h555;
rom[15245] = 12'h555;
rom[15246] = 12'h555;
rom[15247] = 12'h555;
rom[15248] = 12'h555;
rom[15249] = 12'h555;
rom[15250] = 12'h555;
rom[15251] = 12'h555;
rom[15252] = 12'h555;
rom[15253] = 12'h555;
rom[15254] = 12'h555;
rom[15255] = 12'h555;
rom[15256] = 12'h555;
rom[15257] = 12'h555;
rom[15258] = 12'h555;
rom[15259] = 12'h555;
rom[15260] = 12'h555;
rom[15261] = 12'h555;
rom[15262] = 12'h555;
rom[15263] = 12'h555;
rom[15264] = 12'h555;
rom[15265] = 12'h555;
rom[15266] = 12'h555;
rom[15267] = 12'h666;
rom[15268] = 12'h666;
rom[15269] = 12'h777;
rom[15270] = 12'h666;
rom[15271] = 12'h666;
rom[15272] = 12'h666;
rom[15273] = 12'h666;
rom[15274] = 12'h666;
rom[15275] = 12'h777;
rom[15276] = 12'h777;
rom[15277] = 12'h777;
rom[15278] = 12'h666;
rom[15279] = 12'h666;
rom[15280] = 12'h555;
rom[15281] = 12'h555;
rom[15282] = 12'h555;
rom[15283] = 12'h555;
rom[15284] = 12'h444;
rom[15285] = 12'h444;
rom[15286] = 12'h333;
rom[15287] = 12'h333;
rom[15288] = 12'h222;
rom[15289] = 12'h222;
rom[15290] = 12'h222;
rom[15291] = 12'h111;
rom[15292] = 12'h111;
rom[15293] = 12'h111;
rom[15294] = 12'h111;
rom[15295] = 12'h111;
rom[15296] = 12'h100;
rom[15297] = 12'h  0;
rom[15298] = 12'h  0;
rom[15299] = 12'h  0;
rom[15300] = 12'h  0;
rom[15301] = 12'h  0;
rom[15302] = 12'h  0;
rom[15303] = 12'h  0;
rom[15304] = 12'h  0;
rom[15305] = 12'h  0;
rom[15306] = 12'h  0;
rom[15307] = 12'h  0;
rom[15308] = 12'h  0;
rom[15309] = 12'h  0;
rom[15310] = 12'h  0;
rom[15311] = 12'h  0;
rom[15312] = 12'h  0;
rom[15313] = 12'h  0;
rom[15314] = 12'h100;
rom[15315] = 12'h200;
rom[15316] = 12'h300;
rom[15317] = 12'h400;
rom[15318] = 12'h510;
rom[15319] = 12'h610;
rom[15320] = 12'h820;
rom[15321] = 12'h820;
rom[15322] = 12'h820;
rom[15323] = 12'h921;
rom[15324] = 12'h931;
rom[15325] = 12'h920;
rom[15326] = 12'h920;
rom[15327] = 12'h810;
rom[15328] = 12'h610;
rom[15329] = 12'h600;
rom[15330] = 12'h500;
rom[15331] = 12'h500;
rom[15332] = 12'h500;
rom[15333] = 12'h500;
rom[15334] = 12'h500;
rom[15335] = 12'h400;
rom[15336] = 12'h400;
rom[15337] = 12'h400;
rom[15338] = 12'h400;
rom[15339] = 12'h300;
rom[15340] = 12'h300;
rom[15341] = 12'h200;
rom[15342] = 12'h200;
rom[15343] = 12'h100;
rom[15344] = 12'h100;
rom[15345] = 12'h  0;
rom[15346] = 12'h  0;
rom[15347] = 12'h  0;
rom[15348] = 12'h  0;
rom[15349] = 12'h  0;
rom[15350] = 12'h  0;
rom[15351] = 12'h  0;
rom[15352] = 12'h  0;
rom[15353] = 12'h  0;
rom[15354] = 12'h  0;
rom[15355] = 12'h  0;
rom[15356] = 12'h  0;
rom[15357] = 12'h  0;
rom[15358] = 12'h  0;
rom[15359] = 12'h  0;
rom[15360] = 12'h100;
rom[15361] = 12'h100;
rom[15362] = 12'h100;
rom[15363] = 12'h100;
rom[15364] = 12'h100;
rom[15365] = 12'h100;
rom[15366] = 12'h100;
rom[15367] = 12'h100;
rom[15368] = 12'h100;
rom[15369] = 12'h100;
rom[15370] = 12'h100;
rom[15371] = 12'h200;
rom[15372] = 12'h200;
rom[15373] = 12'h200;
rom[15374] = 12'h200;
rom[15375] = 12'h200;
rom[15376] = 12'h200;
rom[15377] = 12'h200;
rom[15378] = 12'h300;
rom[15379] = 12'h300;
rom[15380] = 12'h300;
rom[15381] = 12'h300;
rom[15382] = 12'h300;
rom[15383] = 12'h300;
rom[15384] = 12'h300;
rom[15385] = 12'h300;
rom[15386] = 12'h300;
rom[15387] = 12'h300;
rom[15388] = 12'h300;
rom[15389] = 12'h310;
rom[15390] = 12'h311;
rom[15391] = 12'h311;
rom[15392] = 12'h322;
rom[15393] = 12'h333;
rom[15394] = 12'h544;
rom[15395] = 12'h766;
rom[15396] = 12'h888;
rom[15397] = 12'haaa;
rom[15398] = 12'hbbb;
rom[15399] = 12'hccc;
rom[15400] = 12'hcbb;
rom[15401] = 12'hcbb;
rom[15402] = 12'hbbb;
rom[15403] = 12'hbbb;
rom[15404] = 12'hbbb;
rom[15405] = 12'hbbb;
rom[15406] = 12'haaa;
rom[15407] = 12'h999;
rom[15408] = 12'h999;
rom[15409] = 12'h898;
rom[15410] = 12'h888;
rom[15411] = 12'h888;
rom[15412] = 12'h788;
rom[15413] = 12'h788;
rom[15414] = 12'h787;
rom[15415] = 12'h777;
rom[15416] = 12'h777;
rom[15417] = 12'h777;
rom[15418] = 12'h777;
rom[15419] = 12'h777;
rom[15420] = 12'h777;
rom[15421] = 12'h777;
rom[15422] = 12'h777;
rom[15423] = 12'h777;
rom[15424] = 12'h777;
rom[15425] = 12'h888;
rom[15426] = 12'h888;
rom[15427] = 12'h888;
rom[15428] = 12'h888;
rom[15429] = 12'h777;
rom[15430] = 12'h666;
rom[15431] = 12'h666;
rom[15432] = 12'h666;
rom[15433] = 12'h666;
rom[15434] = 12'h777;
rom[15435] = 12'h777;
rom[15436] = 12'h666;
rom[15437] = 12'h666;
rom[15438] = 12'h666;
rom[15439] = 12'h666;
rom[15440] = 12'h666;
rom[15441] = 12'h666;
rom[15442] = 12'h666;
rom[15443] = 12'h555;
rom[15444] = 12'h555;
rom[15445] = 12'h555;
rom[15446] = 12'h555;
rom[15447] = 12'h555;
rom[15448] = 12'h555;
rom[15449] = 12'h555;
rom[15450] = 12'h555;
rom[15451] = 12'h444;
rom[15452] = 12'h444;
rom[15453] = 12'h444;
rom[15454] = 12'h333;
rom[15455] = 12'h333;
rom[15456] = 12'h222;
rom[15457] = 12'h222;
rom[15458] = 12'h222;
rom[15459] = 12'h111;
rom[15460] = 12'h111;
rom[15461] = 12'h111;
rom[15462] = 12'h111;
rom[15463] = 12'h111;
rom[15464] = 12'h111;
rom[15465] = 12'h111;
rom[15466] = 12'h  0;
rom[15467] = 12'h  0;
rom[15468] = 12'h  0;
rom[15469] = 12'h  0;
rom[15470] = 12'h  0;
rom[15471] = 12'h  0;
rom[15472] = 12'h  0;
rom[15473] = 12'h  0;
rom[15474] = 12'h  0;
rom[15475] = 12'h  0;
rom[15476] = 12'h  0;
rom[15477] = 12'h  0;
rom[15478] = 12'h  0;
rom[15479] = 12'h  0;
rom[15480] = 12'h  0;
rom[15481] = 12'h  0;
rom[15482] = 12'h  0;
rom[15483] = 12'h  0;
rom[15484] = 12'h  0;
rom[15485] = 12'h  0;
rom[15486] = 12'h  0;
rom[15487] = 12'h  0;
rom[15488] = 12'h  0;
rom[15489] = 12'h  0;
rom[15490] = 12'h  0;
rom[15491] = 12'h  0;
rom[15492] = 12'h  0;
rom[15493] = 12'h  0;
rom[15494] = 12'h  0;
rom[15495] = 12'h  0;
rom[15496] = 12'h  0;
rom[15497] = 12'h  0;
rom[15498] = 12'h111;
rom[15499] = 12'h111;
rom[15500] = 12'h111;
rom[15501] = 12'h  0;
rom[15502] = 12'h  0;
rom[15503] = 12'h  0;
rom[15504] = 12'h  0;
rom[15505] = 12'h  0;
rom[15506] = 12'h  0;
rom[15507] = 12'h111;
rom[15508] = 12'h111;
rom[15509] = 12'h111;
rom[15510] = 12'h222;
rom[15511] = 12'h333;
rom[15512] = 12'h333;
rom[15513] = 12'h444;
rom[15514] = 12'h444;
rom[15515] = 12'h444;
rom[15516] = 12'h444;
rom[15517] = 12'h444;
rom[15518] = 12'h444;
rom[15519] = 12'h444;
rom[15520] = 12'h333;
rom[15521] = 12'h333;
rom[15522] = 12'h444;
rom[15523] = 12'h444;
rom[15524] = 12'h444;
rom[15525] = 12'h333;
rom[15526] = 12'h333;
rom[15527] = 12'h333;
rom[15528] = 12'h333;
rom[15529] = 12'h222;
rom[15530] = 12'h111;
rom[15531] = 12'h111;
rom[15532] = 12'h111;
rom[15533] = 12'h  0;
rom[15534] = 12'h  0;
rom[15535] = 12'h  0;
rom[15536] = 12'h  0;
rom[15537] = 12'h  0;
rom[15538] = 12'h  0;
rom[15539] = 12'h  0;
rom[15540] = 12'h  0;
rom[15541] = 12'h  0;
rom[15542] = 12'h  0;
rom[15543] = 12'h  0;
rom[15544] = 12'h  0;
rom[15545] = 12'h111;
rom[15546] = 12'h111;
rom[15547] = 12'h111;
rom[15548] = 12'h222;
rom[15549] = 12'h333;
rom[15550] = 12'h444;
rom[15551] = 12'h555;
rom[15552] = 12'h666;
rom[15553] = 12'h666;
rom[15554] = 12'h666;
rom[15555] = 12'h666;
rom[15556] = 12'h666;
rom[15557] = 12'h555;
rom[15558] = 12'h555;
rom[15559] = 12'h555;
rom[15560] = 12'h555;
rom[15561] = 12'h555;
rom[15562] = 12'h555;
rom[15563] = 12'h555;
rom[15564] = 12'h555;
rom[15565] = 12'h555;
rom[15566] = 12'h666;
rom[15567] = 12'h666;
rom[15568] = 12'h666;
rom[15569] = 12'h666;
rom[15570] = 12'h666;
rom[15571] = 12'h666;
rom[15572] = 12'h555;
rom[15573] = 12'h555;
rom[15574] = 12'h555;
rom[15575] = 12'h555;
rom[15576] = 12'h555;
rom[15577] = 12'h555;
rom[15578] = 12'h555;
rom[15579] = 12'h555;
rom[15580] = 12'h555;
rom[15581] = 12'h555;
rom[15582] = 12'h555;
rom[15583] = 12'h555;
rom[15584] = 12'h555;
rom[15585] = 12'h666;
rom[15586] = 12'h666;
rom[15587] = 12'h666;
rom[15588] = 12'h777;
rom[15589] = 12'h777;
rom[15590] = 12'h777;
rom[15591] = 12'h777;
rom[15592] = 12'h777;
rom[15593] = 12'h888;
rom[15594] = 12'h888;
rom[15595] = 12'h999;
rom[15596] = 12'haaa;
rom[15597] = 12'haaa;
rom[15598] = 12'haaa;
rom[15599] = 12'haaa;
rom[15600] = 12'h222;
rom[15601] = 12'h222;
rom[15602] = 12'h222;
rom[15603] = 12'h222;
rom[15604] = 12'h222;
rom[15605] = 12'h222;
rom[15606] = 12'h222;
rom[15607] = 12'h222;
rom[15608] = 12'h222;
rom[15609] = 12'h222;
rom[15610] = 12'h111;
rom[15611] = 12'h111;
rom[15612] = 12'h111;
rom[15613] = 12'h111;
rom[15614] = 12'h111;
rom[15615] = 12'h111;
rom[15616] = 12'h222;
rom[15617] = 12'h222;
rom[15618] = 12'h222;
rom[15619] = 12'h222;
rom[15620] = 12'h222;
rom[15621] = 12'h222;
rom[15622] = 12'h222;
rom[15623] = 12'h222;
rom[15624] = 12'h333;
rom[15625] = 12'h333;
rom[15626] = 12'h333;
rom[15627] = 12'h333;
rom[15628] = 12'h333;
rom[15629] = 12'h333;
rom[15630] = 12'h444;
rom[15631] = 12'h444;
rom[15632] = 12'h444;
rom[15633] = 12'h444;
rom[15634] = 12'h444;
rom[15635] = 12'h444;
rom[15636] = 12'h444;
rom[15637] = 12'h444;
rom[15638] = 12'h555;
rom[15639] = 12'h555;
rom[15640] = 12'h555;
rom[15641] = 12'h555;
rom[15642] = 12'h555;
rom[15643] = 12'h555;
rom[15644] = 12'h555;
rom[15645] = 12'h666;
rom[15646] = 12'h666;
rom[15647] = 12'h666;
rom[15648] = 12'h666;
rom[15649] = 12'h666;
rom[15650] = 12'h666;
rom[15651] = 12'h666;
rom[15652] = 12'h555;
rom[15653] = 12'h555;
rom[15654] = 12'h555;
rom[15655] = 12'h555;
rom[15656] = 12'h555;
rom[15657] = 12'h555;
rom[15658] = 12'h555;
rom[15659] = 12'h555;
rom[15660] = 12'h555;
rom[15661] = 12'h555;
rom[15662] = 12'h555;
rom[15663] = 12'h555;
rom[15664] = 12'h444;
rom[15665] = 12'h444;
rom[15666] = 12'h555;
rom[15667] = 12'h666;
rom[15668] = 12'h666;
rom[15669] = 12'h777;
rom[15670] = 12'h777;
rom[15671] = 12'h666;
rom[15672] = 12'h666;
rom[15673] = 12'h666;
rom[15674] = 12'h666;
rom[15675] = 12'h777;
rom[15676] = 12'h777;
rom[15677] = 12'h777;
rom[15678] = 12'h777;
rom[15679] = 12'h666;
rom[15680] = 12'h666;
rom[15681] = 12'h666;
rom[15682] = 12'h555;
rom[15683] = 12'h555;
rom[15684] = 12'h444;
rom[15685] = 12'h444;
rom[15686] = 12'h333;
rom[15687] = 12'h333;
rom[15688] = 12'h222;
rom[15689] = 12'h222;
rom[15690] = 12'h222;
rom[15691] = 12'h111;
rom[15692] = 12'h111;
rom[15693] = 12'h111;
rom[15694] = 12'h111;
rom[15695] = 12'h111;
rom[15696] = 12'h100;
rom[15697] = 12'h  0;
rom[15698] = 12'h  0;
rom[15699] = 12'h  0;
rom[15700] = 12'h  0;
rom[15701] = 12'h  0;
rom[15702] = 12'h  0;
rom[15703] = 12'h  0;
rom[15704] = 12'h  0;
rom[15705] = 12'h  0;
rom[15706] = 12'h  0;
rom[15707] = 12'h  0;
rom[15708] = 12'h  0;
rom[15709] = 12'h  0;
rom[15710] = 12'h  0;
rom[15711] = 12'h  0;
rom[15712] = 12'h  0;
rom[15713] = 12'h  0;
rom[15714] = 12'h100;
rom[15715] = 12'h200;
rom[15716] = 12'h300;
rom[15717] = 12'h300;
rom[15718] = 12'h510;
rom[15719] = 12'h610;
rom[15720] = 12'h821;
rom[15721] = 12'h820;
rom[15722] = 12'h820;
rom[15723] = 12'h920;
rom[15724] = 12'h931;
rom[15725] = 12'h920;
rom[15726] = 12'h920;
rom[15727] = 12'h810;
rom[15728] = 12'h710;
rom[15729] = 12'h600;
rom[15730] = 12'h600;
rom[15731] = 12'h500;
rom[15732] = 12'h500;
rom[15733] = 12'h500;
rom[15734] = 12'h500;
rom[15735] = 12'h500;
rom[15736] = 12'h400;
rom[15737] = 12'h400;
rom[15738] = 12'h300;
rom[15739] = 12'h300;
rom[15740] = 12'h300;
rom[15741] = 12'h200;
rom[15742] = 12'h200;
rom[15743] = 12'h100;
rom[15744] = 12'h  0;
rom[15745] = 12'h  0;
rom[15746] = 12'h  0;
rom[15747] = 12'h  0;
rom[15748] = 12'h  0;
rom[15749] = 12'h  0;
rom[15750] = 12'h  0;
rom[15751] = 12'h  0;
rom[15752] = 12'h  0;
rom[15753] = 12'h  0;
rom[15754] = 12'h  0;
rom[15755] = 12'h  0;
rom[15756] = 12'h  0;
rom[15757] = 12'h  0;
rom[15758] = 12'h  0;
rom[15759] = 12'h  0;
rom[15760] = 12'h  0;
rom[15761] = 12'h100;
rom[15762] = 12'h100;
rom[15763] = 12'h100;
rom[15764] = 12'h100;
rom[15765] = 12'h100;
rom[15766] = 12'h100;
rom[15767] = 12'h100;
rom[15768] = 12'h100;
rom[15769] = 12'h100;
rom[15770] = 12'h100;
rom[15771] = 12'h200;
rom[15772] = 12'h200;
rom[15773] = 12'h200;
rom[15774] = 12'h200;
rom[15775] = 12'h200;
rom[15776] = 12'h200;
rom[15777] = 12'h200;
rom[15778] = 12'h300;
rom[15779] = 12'h300;
rom[15780] = 12'h300;
rom[15781] = 12'h300;
rom[15782] = 12'h300;
rom[15783] = 12'h300;
rom[15784] = 12'h300;
rom[15785] = 12'h300;
rom[15786] = 12'h400;
rom[15787] = 12'h410;
rom[15788] = 12'h410;
rom[15789] = 12'h410;
rom[15790] = 12'h411;
rom[15791] = 12'h311;
rom[15792] = 12'h211;
rom[15793] = 12'h222;
rom[15794] = 12'h433;
rom[15795] = 12'h655;
rom[15796] = 12'h877;
rom[15797] = 12'h999;
rom[15798] = 12'hbaa;
rom[15799] = 12'hcbb;
rom[15800] = 12'hcbc;
rom[15801] = 12'hcbb;
rom[15802] = 12'hbbb;
rom[15803] = 12'hbbb;
rom[15804] = 12'hbbb;
rom[15805] = 12'hbbb;
rom[15806] = 12'haaa;
rom[15807] = 12'h9aa;
rom[15808] = 12'h999;
rom[15809] = 12'h899;
rom[15810] = 12'h888;
rom[15811] = 12'h888;
rom[15812] = 12'h888;
rom[15813] = 12'h888;
rom[15814] = 12'h788;
rom[15815] = 12'h788;
rom[15816] = 12'h777;
rom[15817] = 12'h777;
rom[15818] = 12'h777;
rom[15819] = 12'h777;
rom[15820] = 12'h777;
rom[15821] = 12'h777;
rom[15822] = 12'h877;
rom[15823] = 12'h888;
rom[15824] = 12'h888;
rom[15825] = 12'h888;
rom[15826] = 12'h888;
rom[15827] = 12'h777;
rom[15828] = 12'h777;
rom[15829] = 12'h666;
rom[15830] = 12'h666;
rom[15831] = 12'h666;
rom[15832] = 12'h666;
rom[15833] = 12'h777;
rom[15834] = 12'h777;
rom[15835] = 12'h777;
rom[15836] = 12'h666;
rom[15837] = 12'h666;
rom[15838] = 12'h666;
rom[15839] = 12'h666;
rom[15840] = 12'h555;
rom[15841] = 12'h666;
rom[15842] = 12'h666;
rom[15843] = 12'h555;
rom[15844] = 12'h555;
rom[15845] = 12'h555;
rom[15846] = 12'h555;
rom[15847] = 12'h555;
rom[15848] = 12'h555;
rom[15849] = 12'h555;
rom[15850] = 12'h555;
rom[15851] = 12'h555;
rom[15852] = 12'h444;
rom[15853] = 12'h333;
rom[15854] = 12'h333;
rom[15855] = 12'h222;
rom[15856] = 12'h222;
rom[15857] = 12'h222;
rom[15858] = 12'h222;
rom[15859] = 12'h111;
rom[15860] = 12'h111;
rom[15861] = 12'h111;
rom[15862] = 12'h111;
rom[15863] = 12'h111;
rom[15864] = 12'h  0;
rom[15865] = 12'h  0;
rom[15866] = 12'h  0;
rom[15867] = 12'h  0;
rom[15868] = 12'h  0;
rom[15869] = 12'h  0;
rom[15870] = 12'h  0;
rom[15871] = 12'h  0;
rom[15872] = 12'h  0;
rom[15873] = 12'h  0;
rom[15874] = 12'h  0;
rom[15875] = 12'h  0;
rom[15876] = 12'h  0;
rom[15877] = 12'h  0;
rom[15878] = 12'h  0;
rom[15879] = 12'h  0;
rom[15880] = 12'h  0;
rom[15881] = 12'h  0;
rom[15882] = 12'h  0;
rom[15883] = 12'h  0;
rom[15884] = 12'h  0;
rom[15885] = 12'h  0;
rom[15886] = 12'h  0;
rom[15887] = 12'h  0;
rom[15888] = 12'h  0;
rom[15889] = 12'h  0;
rom[15890] = 12'h  0;
rom[15891] = 12'h  0;
rom[15892] = 12'h  0;
rom[15893] = 12'h  0;
rom[15894] = 12'h  0;
rom[15895] = 12'h  0;
rom[15896] = 12'h  0;
rom[15897] = 12'h  0;
rom[15898] = 12'h111;
rom[15899] = 12'h111;
rom[15900] = 12'h111;
rom[15901] = 12'h  0;
rom[15902] = 12'h  0;
rom[15903] = 12'h  0;
rom[15904] = 12'h  0;
rom[15905] = 12'h  0;
rom[15906] = 12'h111;
rom[15907] = 12'h111;
rom[15908] = 12'h111;
rom[15909] = 12'h111;
rom[15910] = 12'h222;
rom[15911] = 12'h333;
rom[15912] = 12'h444;
rom[15913] = 12'h444;
rom[15914] = 12'h444;
rom[15915] = 12'h444;
rom[15916] = 12'h444;
rom[15917] = 12'h444;
rom[15918] = 12'h444;
rom[15919] = 12'h444;
rom[15920] = 12'h444;
rom[15921] = 12'h333;
rom[15922] = 12'h444;
rom[15923] = 12'h444;
rom[15924] = 12'h444;
rom[15925] = 12'h333;
rom[15926] = 12'h333;
rom[15927] = 12'h333;
rom[15928] = 12'h333;
rom[15929] = 12'h222;
rom[15930] = 12'h111;
rom[15931] = 12'h111;
rom[15932] = 12'h111;
rom[15933] = 12'h  0;
rom[15934] = 12'h  0;
rom[15935] = 12'h  0;
rom[15936] = 12'h  0;
rom[15937] = 12'h  0;
rom[15938] = 12'h  0;
rom[15939] = 12'h  0;
rom[15940] = 12'h  0;
rom[15941] = 12'h  0;
rom[15942] = 12'h  0;
rom[15943] = 12'h  0;
rom[15944] = 12'h  0;
rom[15945] = 12'h111;
rom[15946] = 12'h111;
rom[15947] = 12'h222;
rom[15948] = 12'h222;
rom[15949] = 12'h333;
rom[15950] = 12'h444;
rom[15951] = 12'h555;
rom[15952] = 12'h666;
rom[15953] = 12'h666;
rom[15954] = 12'h666;
rom[15955] = 12'h666;
rom[15956] = 12'h555;
rom[15957] = 12'h555;
rom[15958] = 12'h555;
rom[15959] = 12'h555;
rom[15960] = 12'h555;
rom[15961] = 12'h555;
rom[15962] = 12'h555;
rom[15963] = 12'h555;
rom[15964] = 12'h555;
rom[15965] = 12'h666;
rom[15966] = 12'h666;
rom[15967] = 12'h666;
rom[15968] = 12'h777;
rom[15969] = 12'h666;
rom[15970] = 12'h666;
rom[15971] = 12'h666;
rom[15972] = 12'h666;
rom[15973] = 12'h666;
rom[15974] = 12'h666;
rom[15975] = 12'h666;
rom[15976] = 12'h666;
rom[15977] = 12'h666;
rom[15978] = 12'h666;
rom[15979] = 12'h555;
rom[15980] = 12'h555;
rom[15981] = 12'h555;
rom[15982] = 12'h555;
rom[15983] = 12'h555;
rom[15984] = 12'h555;
rom[15985] = 12'h555;
rom[15986] = 12'h666;
rom[15987] = 12'h666;
rom[15988] = 12'h666;
rom[15989] = 12'h777;
rom[15990] = 12'h777;
rom[15991] = 12'h777;
rom[15992] = 12'h777;
rom[15993] = 12'h888;
rom[15994] = 12'h888;
rom[15995] = 12'h999;
rom[15996] = 12'haaa;
rom[15997] = 12'haaa;
rom[15998] = 12'haaa;
rom[15999] = 12'haaa;
rom[16000] = 12'h222;
rom[16001] = 12'h222;
rom[16002] = 12'h222;
rom[16003] = 12'h222;
rom[16004] = 12'h222;
rom[16005] = 12'h222;
rom[16006] = 12'h222;
rom[16007] = 12'h222;
rom[16008] = 12'h222;
rom[16009] = 12'h222;
rom[16010] = 12'h222;
rom[16011] = 12'h222;
rom[16012] = 12'h222;
rom[16013] = 12'h222;
rom[16014] = 12'h222;
rom[16015] = 12'h222;
rom[16016] = 12'h222;
rom[16017] = 12'h222;
rom[16018] = 12'h222;
rom[16019] = 12'h222;
rom[16020] = 12'h222;
rom[16021] = 12'h222;
rom[16022] = 12'h222;
rom[16023] = 12'h333;
rom[16024] = 12'h222;
rom[16025] = 12'h333;
rom[16026] = 12'h333;
rom[16027] = 12'h444;
rom[16028] = 12'h444;
rom[16029] = 12'h444;
rom[16030] = 12'h444;
rom[16031] = 12'h444;
rom[16032] = 12'h444;
rom[16033] = 12'h444;
rom[16034] = 12'h444;
rom[16035] = 12'h444;
rom[16036] = 12'h555;
rom[16037] = 12'h555;
rom[16038] = 12'h555;
rom[16039] = 12'h555;
rom[16040] = 12'h555;
rom[16041] = 12'h555;
rom[16042] = 12'h666;
rom[16043] = 12'h666;
rom[16044] = 12'h666;
rom[16045] = 12'h666;
rom[16046] = 12'h666;
rom[16047] = 12'h666;
rom[16048] = 12'h666;
rom[16049] = 12'h666;
rom[16050] = 12'h666;
rom[16051] = 12'h666;
rom[16052] = 12'h666;
rom[16053] = 12'h555;
rom[16054] = 12'h555;
rom[16055] = 12'h555;
rom[16056] = 12'h555;
rom[16057] = 12'h555;
rom[16058] = 12'h555;
rom[16059] = 12'h555;
rom[16060] = 12'h555;
rom[16061] = 12'h555;
rom[16062] = 12'h555;
rom[16063] = 12'h555;
rom[16064] = 12'h555;
rom[16065] = 12'h555;
rom[16066] = 12'h555;
rom[16067] = 12'h555;
rom[16068] = 12'h666;
rom[16069] = 12'h666;
rom[16070] = 12'h777;
rom[16071] = 12'h777;
rom[16072] = 12'h666;
rom[16073] = 12'h666;
rom[16074] = 12'h666;
rom[16075] = 12'h777;
rom[16076] = 12'h777;
rom[16077] = 12'h777;
rom[16078] = 12'h777;
rom[16079] = 12'h777;
rom[16080] = 12'h666;
rom[16081] = 12'h555;
rom[16082] = 12'h555;
rom[16083] = 12'h555;
rom[16084] = 12'h555;
rom[16085] = 12'h444;
rom[16086] = 12'h333;
rom[16087] = 12'h333;
rom[16088] = 12'h333;
rom[16089] = 12'h333;
rom[16090] = 12'h222;
rom[16091] = 12'h222;
rom[16092] = 12'h111;
rom[16093] = 12'h111;
rom[16094] = 12'h111;
rom[16095] = 12'h111;
rom[16096] = 12'h  0;
rom[16097] = 12'h  0;
rom[16098] = 12'h  0;
rom[16099] = 12'h  0;
rom[16100] = 12'h  0;
rom[16101] = 12'h  0;
rom[16102] = 12'h  0;
rom[16103] = 12'h  0;
rom[16104] = 12'h  0;
rom[16105] = 12'h  0;
rom[16106] = 12'h  0;
rom[16107] = 12'h  0;
rom[16108] = 12'h  0;
rom[16109] = 12'h  0;
rom[16110] = 12'h  0;
rom[16111] = 12'h  0;
rom[16112] = 12'h  0;
rom[16113] = 12'h  0;
rom[16114] = 12'h100;
rom[16115] = 12'h200;
rom[16116] = 12'h300;
rom[16117] = 12'h300;
rom[16118] = 12'h510;
rom[16119] = 12'h610;
rom[16120] = 12'h720;
rom[16121] = 12'h820;
rom[16122] = 12'h920;
rom[16123] = 12'h921;
rom[16124] = 12'h931;
rom[16125] = 12'h920;
rom[16126] = 12'h920;
rom[16127] = 12'h810;
rom[16128] = 12'h710;
rom[16129] = 12'h610;
rom[16130] = 12'h600;
rom[16131] = 12'h600;
rom[16132] = 12'h500;
rom[16133] = 12'h500;
rom[16134] = 12'h500;
rom[16135] = 12'h500;
rom[16136] = 12'h400;
rom[16137] = 12'h400;
rom[16138] = 12'h300;
rom[16139] = 12'h300;
rom[16140] = 12'h200;
rom[16141] = 12'h200;
rom[16142] = 12'h200;
rom[16143] = 12'h100;
rom[16144] = 12'h  0;
rom[16145] = 12'h  0;
rom[16146] = 12'h  0;
rom[16147] = 12'h  0;
rom[16148] = 12'h  0;
rom[16149] = 12'h  0;
rom[16150] = 12'h  0;
rom[16151] = 12'h  0;
rom[16152] = 12'h  0;
rom[16153] = 12'h  0;
rom[16154] = 12'h  0;
rom[16155] = 12'h  0;
rom[16156] = 12'h  0;
rom[16157] = 12'h  0;
rom[16158] = 12'h  0;
rom[16159] = 12'h  0;
rom[16160] = 12'h  0;
rom[16161] = 12'h  0;
rom[16162] = 12'h  0;
rom[16163] = 12'h  0;
rom[16164] = 12'h  0;
rom[16165] = 12'h100;
rom[16166] = 12'h100;
rom[16167] = 12'h100;
rom[16168] = 12'h100;
rom[16169] = 12'h100;
rom[16170] = 12'h200;
rom[16171] = 12'h200;
rom[16172] = 12'h200;
rom[16173] = 12'h200;
rom[16174] = 12'h200;
rom[16175] = 12'h200;
rom[16176] = 12'h200;
rom[16177] = 12'h200;
rom[16178] = 12'h200;
rom[16179] = 12'h300;
rom[16180] = 12'h300;
rom[16181] = 12'h300;
rom[16182] = 12'h300;
rom[16183] = 12'h300;
rom[16184] = 12'h300;
rom[16185] = 12'h300;
rom[16186] = 12'h300;
rom[16187] = 12'h300;
rom[16188] = 12'h300;
rom[16189] = 12'h300;
rom[16190] = 12'h410;
rom[16191] = 12'h311;
rom[16192] = 12'h211;
rom[16193] = 12'h211;
rom[16194] = 12'h322;
rom[16195] = 12'h444;
rom[16196] = 12'h666;
rom[16197] = 12'h988;
rom[16198] = 12'haaa;
rom[16199] = 12'hbab;
rom[16200] = 12'hbbb;
rom[16201] = 12'hcbb;
rom[16202] = 12'hcbb;
rom[16203] = 12'hbbb;
rom[16204] = 12'hbbb;
rom[16205] = 12'hbbb;
rom[16206] = 12'hbaa;
rom[16207] = 12'haaa;
rom[16208] = 12'h999;
rom[16209] = 12'h999;
rom[16210] = 12'h899;
rom[16211] = 12'h899;
rom[16212] = 12'h888;
rom[16213] = 12'h888;
rom[16214] = 12'h788;
rom[16215] = 12'h777;
rom[16216] = 12'h777;
rom[16217] = 12'h777;
rom[16218] = 12'h777;
rom[16219] = 12'h777;
rom[16220] = 12'h888;
rom[16221] = 12'h888;
rom[16222] = 12'h888;
rom[16223] = 12'h888;
rom[16224] = 12'h999;
rom[16225] = 12'h888;
rom[16226] = 12'h777;
rom[16227] = 12'h666;
rom[16228] = 12'h666;
rom[16229] = 12'h666;
rom[16230] = 12'h777;
rom[16231] = 12'h777;
rom[16232] = 12'h777;
rom[16233] = 12'h777;
rom[16234] = 12'h666;
rom[16235] = 12'h666;
rom[16236] = 12'h666;
rom[16237] = 12'h666;
rom[16238] = 12'h555;
rom[16239] = 12'h555;
rom[16240] = 12'h555;
rom[16241] = 12'h555;
rom[16242] = 12'h555;
rom[16243] = 12'h555;
rom[16244] = 12'h555;
rom[16245] = 12'h555;
rom[16246] = 12'h555;
rom[16247] = 12'h555;
rom[16248] = 12'h555;
rom[16249] = 12'h555;
rom[16250] = 12'h555;
rom[16251] = 12'h444;
rom[16252] = 12'h333;
rom[16253] = 12'h333;
rom[16254] = 12'h222;
rom[16255] = 12'h222;
rom[16256] = 12'h222;
rom[16257] = 12'h222;
rom[16258] = 12'h111;
rom[16259] = 12'h111;
rom[16260] = 12'h111;
rom[16261] = 12'h111;
rom[16262] = 12'h111;
rom[16263] = 12'h111;
rom[16264] = 12'h111;
rom[16265] = 12'h111;
rom[16266] = 12'h  0;
rom[16267] = 12'h  0;
rom[16268] = 12'h  0;
rom[16269] = 12'h  0;
rom[16270] = 12'h  0;
rom[16271] = 12'h  0;
rom[16272] = 12'h  0;
rom[16273] = 12'h  0;
rom[16274] = 12'h  0;
rom[16275] = 12'h  0;
rom[16276] = 12'h  0;
rom[16277] = 12'h  0;
rom[16278] = 12'h  0;
rom[16279] = 12'h  0;
rom[16280] = 12'h  0;
rom[16281] = 12'h  0;
rom[16282] = 12'h  0;
rom[16283] = 12'h  0;
rom[16284] = 12'h  0;
rom[16285] = 12'h  0;
rom[16286] = 12'h  0;
rom[16287] = 12'h  0;
rom[16288] = 12'h  0;
rom[16289] = 12'h  0;
rom[16290] = 12'h  0;
rom[16291] = 12'h  0;
rom[16292] = 12'h  0;
rom[16293] = 12'h  0;
rom[16294] = 12'h  0;
rom[16295] = 12'h  0;
rom[16296] = 12'h  0;
rom[16297] = 12'h111;
rom[16298] = 12'h111;
rom[16299] = 12'h111;
rom[16300] = 12'h111;
rom[16301] = 12'h  0;
rom[16302] = 12'h  0;
rom[16303] = 12'h  0;
rom[16304] = 12'h  0;
rom[16305] = 12'h111;
rom[16306] = 12'h111;
rom[16307] = 12'h111;
rom[16308] = 12'h111;
rom[16309] = 12'h222;
rom[16310] = 12'h333;
rom[16311] = 12'h333;
rom[16312] = 12'h444;
rom[16313] = 12'h444;
rom[16314] = 12'h444;
rom[16315] = 12'h444;
rom[16316] = 12'h333;
rom[16317] = 12'h333;
rom[16318] = 12'h333;
rom[16319] = 12'h444;
rom[16320] = 12'h333;
rom[16321] = 12'h333;
rom[16322] = 12'h333;
rom[16323] = 12'h333;
rom[16324] = 12'h333;
rom[16325] = 12'h444;
rom[16326] = 12'h444;
rom[16327] = 12'h333;
rom[16328] = 12'h333;
rom[16329] = 12'h222;
rom[16330] = 12'h111;
rom[16331] = 12'h111;
rom[16332] = 12'h111;
rom[16333] = 12'h111;
rom[16334] = 12'h  0;
rom[16335] = 12'h  0;
rom[16336] = 12'h  0;
rom[16337] = 12'h  0;
rom[16338] = 12'h  0;
rom[16339] = 12'h  0;
rom[16340] = 12'h  0;
rom[16341] = 12'h  0;
rom[16342] = 12'h  0;
rom[16343] = 12'h  0;
rom[16344] = 12'h  0;
rom[16345] = 12'h111;
rom[16346] = 12'h111;
rom[16347] = 12'h222;
rom[16348] = 12'h333;
rom[16349] = 12'h444;
rom[16350] = 12'h555;
rom[16351] = 12'h555;
rom[16352] = 12'h666;
rom[16353] = 12'h666;
rom[16354] = 12'h666;
rom[16355] = 12'h666;
rom[16356] = 12'h555;
rom[16357] = 12'h555;
rom[16358] = 12'h555;
rom[16359] = 12'h555;
rom[16360] = 12'h555;
rom[16361] = 12'h555;
rom[16362] = 12'h555;
rom[16363] = 12'h555;
rom[16364] = 12'h555;
rom[16365] = 12'h666;
rom[16366] = 12'h666;
rom[16367] = 12'h666;
rom[16368] = 12'h666;
rom[16369] = 12'h777;
rom[16370] = 12'h777;
rom[16371] = 12'h777;
rom[16372] = 12'h777;
rom[16373] = 12'h777;
rom[16374] = 12'h777;
rom[16375] = 12'h777;
rom[16376] = 12'h777;
rom[16377] = 12'h777;
rom[16378] = 12'h777;
rom[16379] = 12'h777;
rom[16380] = 12'h666;
rom[16381] = 12'h666;
rom[16382] = 12'h666;
rom[16383] = 12'h666;
rom[16384] = 12'h666;
rom[16385] = 12'h666;
rom[16386] = 12'h666;
rom[16387] = 12'h666;
rom[16388] = 12'h777;
rom[16389] = 12'h777;
rom[16390] = 12'h777;
rom[16391] = 12'h777;
rom[16392] = 12'h777;
rom[16393] = 12'h888;
rom[16394] = 12'h888;
rom[16395] = 12'h999;
rom[16396] = 12'haaa;
rom[16397] = 12'haaa;
rom[16398] = 12'haaa;
rom[16399] = 12'haaa;
rom[16400] = 12'h222;
rom[16401] = 12'h222;
rom[16402] = 12'h222;
rom[16403] = 12'h222;
rom[16404] = 12'h222;
rom[16405] = 12'h222;
rom[16406] = 12'h222;
rom[16407] = 12'h222;
rom[16408] = 12'h222;
rom[16409] = 12'h222;
rom[16410] = 12'h222;
rom[16411] = 12'h222;
rom[16412] = 12'h222;
rom[16413] = 12'h222;
rom[16414] = 12'h222;
rom[16415] = 12'h222;
rom[16416] = 12'h222;
rom[16417] = 12'h222;
rom[16418] = 12'h222;
rom[16419] = 12'h222;
rom[16420] = 12'h222;
rom[16421] = 12'h222;
rom[16422] = 12'h333;
rom[16423] = 12'h333;
rom[16424] = 12'h333;
rom[16425] = 12'h333;
rom[16426] = 12'h333;
rom[16427] = 12'h444;
rom[16428] = 12'h444;
rom[16429] = 12'h444;
rom[16430] = 12'h444;
rom[16431] = 12'h444;
rom[16432] = 12'h444;
rom[16433] = 12'h444;
rom[16434] = 12'h555;
rom[16435] = 12'h555;
rom[16436] = 12'h555;
rom[16437] = 12'h555;
rom[16438] = 12'h555;
rom[16439] = 12'h666;
rom[16440] = 12'h666;
rom[16441] = 12'h666;
rom[16442] = 12'h666;
rom[16443] = 12'h666;
rom[16444] = 12'h666;
rom[16445] = 12'h666;
rom[16446] = 12'h666;
rom[16447] = 12'h666;
rom[16448] = 12'h666;
rom[16449] = 12'h666;
rom[16450] = 12'h666;
rom[16451] = 12'h666;
rom[16452] = 12'h555;
rom[16453] = 12'h555;
rom[16454] = 12'h555;
rom[16455] = 12'h555;
rom[16456] = 12'h555;
rom[16457] = 12'h555;
rom[16458] = 12'h555;
rom[16459] = 12'h555;
rom[16460] = 12'h555;
rom[16461] = 12'h666;
rom[16462] = 12'h666;
rom[16463] = 12'h666;
rom[16464] = 12'h666;
rom[16465] = 12'h666;
rom[16466] = 12'h666;
rom[16467] = 12'h555;
rom[16468] = 12'h555;
rom[16469] = 12'h666;
rom[16470] = 12'h666;
rom[16471] = 12'h777;
rom[16472] = 12'h666;
rom[16473] = 12'h666;
rom[16474] = 12'h666;
rom[16475] = 12'h777;
rom[16476] = 12'h777;
rom[16477] = 12'h777;
rom[16478] = 12'h777;
rom[16479] = 12'h777;
rom[16480] = 12'h777;
rom[16481] = 12'h666;
rom[16482] = 12'h555;
rom[16483] = 12'h555;
rom[16484] = 12'h555;
rom[16485] = 12'h444;
rom[16486] = 12'h333;
rom[16487] = 12'h333;
rom[16488] = 12'h333;
rom[16489] = 12'h222;
rom[16490] = 12'h222;
rom[16491] = 12'h222;
rom[16492] = 12'h111;
rom[16493] = 12'h111;
rom[16494] = 12'h111;
rom[16495] = 12'h111;
rom[16496] = 12'h  0;
rom[16497] = 12'h  0;
rom[16498] = 12'h  0;
rom[16499] = 12'h  0;
rom[16500] = 12'h  0;
rom[16501] = 12'h  0;
rom[16502] = 12'h  0;
rom[16503] = 12'h  0;
rom[16504] = 12'h  0;
rom[16505] = 12'h  0;
rom[16506] = 12'h  0;
rom[16507] = 12'h  0;
rom[16508] = 12'h  0;
rom[16509] = 12'h  0;
rom[16510] = 12'h  0;
rom[16511] = 12'h  0;
rom[16512] = 12'h  0;
rom[16513] = 12'h  0;
rom[16514] = 12'h100;
rom[16515] = 12'h200;
rom[16516] = 12'h200;
rom[16517] = 12'h300;
rom[16518] = 12'h500;
rom[16519] = 12'h610;
rom[16520] = 12'h821;
rom[16521] = 12'h820;
rom[16522] = 12'h920;
rom[16523] = 12'h920;
rom[16524] = 12'h931;
rom[16525] = 12'h920;
rom[16526] = 12'h920;
rom[16527] = 12'h810;
rom[16528] = 12'h810;
rom[16529] = 12'h710;
rom[16530] = 12'h600;
rom[16531] = 12'h600;
rom[16532] = 12'h600;
rom[16533] = 12'h500;
rom[16534] = 12'h500;
rom[16535] = 12'h500;
rom[16536] = 12'h400;
rom[16537] = 12'h400;
rom[16538] = 12'h300;
rom[16539] = 12'h300;
rom[16540] = 12'h200;
rom[16541] = 12'h200;
rom[16542] = 12'h200;
rom[16543] = 12'h100;
rom[16544] = 12'h  0;
rom[16545] = 12'h  0;
rom[16546] = 12'h  0;
rom[16547] = 12'h  0;
rom[16548] = 12'h  0;
rom[16549] = 12'h  0;
rom[16550] = 12'h  0;
rom[16551] = 12'h  0;
rom[16552] = 12'h  0;
rom[16553] = 12'h  0;
rom[16554] = 12'h  0;
rom[16555] = 12'h  0;
rom[16556] = 12'h  0;
rom[16557] = 12'h  0;
rom[16558] = 12'h  0;
rom[16559] = 12'h  0;
rom[16560] = 12'h  0;
rom[16561] = 12'h  0;
rom[16562] = 12'h  0;
rom[16563] = 12'h  0;
rom[16564] = 12'h  0;
rom[16565] = 12'h100;
rom[16566] = 12'h100;
rom[16567] = 12'h100;
rom[16568] = 12'h100;
rom[16569] = 12'h100;
rom[16570] = 12'h200;
rom[16571] = 12'h200;
rom[16572] = 12'h200;
rom[16573] = 12'h200;
rom[16574] = 12'h300;
rom[16575] = 12'h300;
rom[16576] = 12'h200;
rom[16577] = 12'h200;
rom[16578] = 12'h200;
rom[16579] = 12'h300;
rom[16580] = 12'h300;
rom[16581] = 12'h300;
rom[16582] = 12'h300;
rom[16583] = 12'h300;
rom[16584] = 12'h300;
rom[16585] = 12'h300;
rom[16586] = 12'h300;
rom[16587] = 12'h300;
rom[16588] = 12'h300;
rom[16589] = 12'h300;
rom[16590] = 12'h300;
rom[16591] = 12'h300;
rom[16592] = 12'h211;
rom[16593] = 12'h211;
rom[16594] = 12'h222;
rom[16595] = 12'h433;
rom[16596] = 12'h655;
rom[16597] = 12'h877;
rom[16598] = 12'ha99;
rom[16599] = 12'hbaa;
rom[16600] = 12'hbbb;
rom[16601] = 12'hcbb;
rom[16602] = 12'hcbb;
rom[16603] = 12'hbbb;
rom[16604] = 12'hbbb;
rom[16605] = 12'hbbb;
rom[16606] = 12'hbaa;
rom[16607] = 12'haaa;
rom[16608] = 12'h9aa;
rom[16609] = 12'h999;
rom[16610] = 12'h999;
rom[16611] = 12'h899;
rom[16612] = 12'h899;
rom[16613] = 12'h888;
rom[16614] = 12'h888;
rom[16615] = 12'h788;
rom[16616] = 12'h888;
rom[16617] = 12'h888;
rom[16618] = 12'h888;
rom[16619] = 12'h888;
rom[16620] = 12'h888;
rom[16621] = 12'h888;
rom[16622] = 12'h988;
rom[16623] = 12'h888;
rom[16624] = 12'h888;
rom[16625] = 12'h888;
rom[16626] = 12'h777;
rom[16627] = 12'h777;
rom[16628] = 12'h777;
rom[16629] = 12'h777;
rom[16630] = 12'h777;
rom[16631] = 12'h777;
rom[16632] = 12'h777;
rom[16633] = 12'h777;
rom[16634] = 12'h666;
rom[16635] = 12'h666;
rom[16636] = 12'h666;
rom[16637] = 12'h555;
rom[16638] = 12'h555;
rom[16639] = 12'h555;
rom[16640] = 12'h666;
rom[16641] = 12'h666;
rom[16642] = 12'h555;
rom[16643] = 12'h555;
rom[16644] = 12'h555;
rom[16645] = 12'h555;
rom[16646] = 12'h555;
rom[16647] = 12'h555;
rom[16648] = 12'h555;
rom[16649] = 12'h555;
rom[16650] = 12'h444;
rom[16651] = 12'h333;
rom[16652] = 12'h333;
rom[16653] = 12'h222;
rom[16654] = 12'h222;
rom[16655] = 12'h222;
rom[16656] = 12'h222;
rom[16657] = 12'h222;
rom[16658] = 12'h111;
rom[16659] = 12'h111;
rom[16660] = 12'h111;
rom[16661] = 12'h111;
rom[16662] = 12'h111;
rom[16663] = 12'h111;
rom[16664] = 12'h111;
rom[16665] = 12'h111;
rom[16666] = 12'h  0;
rom[16667] = 12'h  0;
rom[16668] = 12'h  0;
rom[16669] = 12'h  0;
rom[16670] = 12'h  0;
rom[16671] = 12'h  0;
rom[16672] = 12'h  0;
rom[16673] = 12'h  0;
rom[16674] = 12'h  0;
rom[16675] = 12'h  0;
rom[16676] = 12'h  0;
rom[16677] = 12'h  0;
rom[16678] = 12'h  0;
rom[16679] = 12'h  0;
rom[16680] = 12'h  0;
rom[16681] = 12'h  0;
rom[16682] = 12'h  0;
rom[16683] = 12'h  0;
rom[16684] = 12'h  0;
rom[16685] = 12'h  0;
rom[16686] = 12'h  0;
rom[16687] = 12'h  0;
rom[16688] = 12'h  0;
rom[16689] = 12'h  0;
rom[16690] = 12'h  0;
rom[16691] = 12'h  0;
rom[16692] = 12'h  0;
rom[16693] = 12'h  0;
rom[16694] = 12'h  0;
rom[16695] = 12'h  0;
rom[16696] = 12'h  0;
rom[16697] = 12'h111;
rom[16698] = 12'h111;
rom[16699] = 12'h111;
rom[16700] = 12'h111;
rom[16701] = 12'h  0;
rom[16702] = 12'h  0;
rom[16703] = 12'h  0;
rom[16704] = 12'h111;
rom[16705] = 12'h111;
rom[16706] = 12'h111;
rom[16707] = 12'h111;
rom[16708] = 12'h222;
rom[16709] = 12'h222;
rom[16710] = 12'h333;
rom[16711] = 12'h333;
rom[16712] = 12'h333;
rom[16713] = 12'h333;
rom[16714] = 12'h333;
rom[16715] = 12'h333;
rom[16716] = 12'h333;
rom[16717] = 12'h333;
rom[16718] = 12'h333;
rom[16719] = 12'h444;
rom[16720] = 12'h333;
rom[16721] = 12'h333;
rom[16722] = 12'h333;
rom[16723] = 12'h333;
rom[16724] = 12'h333;
rom[16725] = 12'h444;
rom[16726] = 12'h444;
rom[16727] = 12'h333;
rom[16728] = 12'h222;
rom[16729] = 12'h222;
rom[16730] = 12'h111;
rom[16731] = 12'h111;
rom[16732] = 12'h111;
rom[16733] = 12'h111;
rom[16734] = 12'h  0;
rom[16735] = 12'h  0;
rom[16736] = 12'h  0;
rom[16737] = 12'h  0;
rom[16738] = 12'h  0;
rom[16739] = 12'h  0;
rom[16740] = 12'h  0;
rom[16741] = 12'h  0;
rom[16742] = 12'h111;
rom[16743] = 12'h111;
rom[16744] = 12'h  0;
rom[16745] = 12'h111;
rom[16746] = 12'h222;
rom[16747] = 12'h222;
rom[16748] = 12'h333;
rom[16749] = 12'h444;
rom[16750] = 12'h555;
rom[16751] = 12'h555;
rom[16752] = 12'h666;
rom[16753] = 12'h666;
rom[16754] = 12'h666;
rom[16755] = 12'h666;
rom[16756] = 12'h666;
rom[16757] = 12'h555;
rom[16758] = 12'h555;
rom[16759] = 12'h555;
rom[16760] = 12'h555;
rom[16761] = 12'h555;
rom[16762] = 12'h555;
rom[16763] = 12'h555;
rom[16764] = 12'h555;
rom[16765] = 12'h555;
rom[16766] = 12'h555;
rom[16767] = 12'h555;
rom[16768] = 12'h555;
rom[16769] = 12'h555;
rom[16770] = 12'h666;
rom[16771] = 12'h666;
rom[16772] = 12'h666;
rom[16773] = 12'h666;
rom[16774] = 12'h777;
rom[16775] = 12'h777;
rom[16776] = 12'h888;
rom[16777] = 12'h888;
rom[16778] = 12'h888;
rom[16779] = 12'h888;
rom[16780] = 12'h888;
rom[16781] = 12'h777;
rom[16782] = 12'h777;
rom[16783] = 12'h777;
rom[16784] = 12'h777;
rom[16785] = 12'h777;
rom[16786] = 12'h777;
rom[16787] = 12'h777;
rom[16788] = 12'h777;
rom[16789] = 12'h777;
rom[16790] = 12'h777;
rom[16791] = 12'h777;
rom[16792] = 12'h888;
rom[16793] = 12'h888;
rom[16794] = 12'h888;
rom[16795] = 12'h999;
rom[16796] = 12'h999;
rom[16797] = 12'haaa;
rom[16798] = 12'haaa;
rom[16799] = 12'haaa;
rom[16800] = 12'h222;
rom[16801] = 12'h222;
rom[16802] = 12'h222;
rom[16803] = 12'h222;
rom[16804] = 12'h222;
rom[16805] = 12'h222;
rom[16806] = 12'h222;
rom[16807] = 12'h222;
rom[16808] = 12'h222;
rom[16809] = 12'h222;
rom[16810] = 12'h222;
rom[16811] = 12'h222;
rom[16812] = 12'h222;
rom[16813] = 12'h222;
rom[16814] = 12'h222;
rom[16815] = 12'h222;
rom[16816] = 12'h222;
rom[16817] = 12'h222;
rom[16818] = 12'h222;
rom[16819] = 12'h222;
rom[16820] = 12'h222;
rom[16821] = 12'h333;
rom[16822] = 12'h333;
rom[16823] = 12'h333;
rom[16824] = 12'h333;
rom[16825] = 12'h333;
rom[16826] = 12'h444;
rom[16827] = 12'h444;
rom[16828] = 12'h444;
rom[16829] = 12'h444;
rom[16830] = 12'h555;
rom[16831] = 12'h555;
rom[16832] = 12'h555;
rom[16833] = 12'h555;
rom[16834] = 12'h555;
rom[16835] = 12'h555;
rom[16836] = 12'h555;
rom[16837] = 12'h666;
rom[16838] = 12'h666;
rom[16839] = 12'h666;
rom[16840] = 12'h666;
rom[16841] = 12'h666;
rom[16842] = 12'h666;
rom[16843] = 12'h666;
rom[16844] = 12'h666;
rom[16845] = 12'h666;
rom[16846] = 12'h666;
rom[16847] = 12'h666;
rom[16848] = 12'h666;
rom[16849] = 12'h666;
rom[16850] = 12'h666;
rom[16851] = 12'h666;
rom[16852] = 12'h555;
rom[16853] = 12'h555;
rom[16854] = 12'h555;
rom[16855] = 12'h555;
rom[16856] = 12'h555;
rom[16857] = 12'h555;
rom[16858] = 12'h555;
rom[16859] = 12'h555;
rom[16860] = 12'h555;
rom[16861] = 12'h666;
rom[16862] = 12'h666;
rom[16863] = 12'h666;
rom[16864] = 12'h666;
rom[16865] = 12'h666;
rom[16866] = 12'h666;
rom[16867] = 12'h666;
rom[16868] = 12'h555;
rom[16869] = 12'h555;
rom[16870] = 12'h666;
rom[16871] = 12'h666;
rom[16872] = 12'h777;
rom[16873] = 12'h777;
rom[16874] = 12'h777;
rom[16875] = 12'h777;
rom[16876] = 12'h777;
rom[16877] = 12'h777;
rom[16878] = 12'h777;
rom[16879] = 12'h777;
rom[16880] = 12'h777;
rom[16881] = 12'h666;
rom[16882] = 12'h666;
rom[16883] = 12'h555;
rom[16884] = 12'h555;
rom[16885] = 12'h444;
rom[16886] = 12'h333;
rom[16887] = 12'h333;
rom[16888] = 12'h333;
rom[16889] = 12'h222;
rom[16890] = 12'h222;
rom[16891] = 12'h222;
rom[16892] = 12'h111;
rom[16893] = 12'h111;
rom[16894] = 12'h111;
rom[16895] = 12'h111;
rom[16896] = 12'h  0;
rom[16897] = 12'h  0;
rom[16898] = 12'h  0;
rom[16899] = 12'h  0;
rom[16900] = 12'h  0;
rom[16901] = 12'h  0;
rom[16902] = 12'h  0;
rom[16903] = 12'h  0;
rom[16904] = 12'h  0;
rom[16905] = 12'h  0;
rom[16906] = 12'h  0;
rom[16907] = 12'h  0;
rom[16908] = 12'h  0;
rom[16909] = 12'h  0;
rom[16910] = 12'h  0;
rom[16911] = 12'h  0;
rom[16912] = 12'h  0;
rom[16913] = 12'h  0;
rom[16914] = 12'h100;
rom[16915] = 12'h100;
rom[16916] = 12'h200;
rom[16917] = 12'h300;
rom[16918] = 12'h500;
rom[16919] = 12'h610;
rom[16920] = 12'h821;
rom[16921] = 12'h821;
rom[16922] = 12'h920;
rom[16923] = 12'h920;
rom[16924] = 12'ha20;
rom[16925] = 12'h920;
rom[16926] = 12'h920;
rom[16927] = 12'h820;
rom[16928] = 12'h820;
rom[16929] = 12'h710;
rom[16930] = 12'h600;
rom[16931] = 12'h600;
rom[16932] = 12'h600;
rom[16933] = 12'h600;
rom[16934] = 12'h500;
rom[16935] = 12'h500;
rom[16936] = 12'h400;
rom[16937] = 12'h400;
rom[16938] = 12'h300;
rom[16939] = 12'h300;
rom[16940] = 12'h200;
rom[16941] = 12'h200;
rom[16942] = 12'h100;
rom[16943] = 12'h100;
rom[16944] = 12'h  0;
rom[16945] = 12'h  0;
rom[16946] = 12'h  0;
rom[16947] = 12'h  0;
rom[16948] = 12'h  0;
rom[16949] = 12'h  0;
rom[16950] = 12'h  0;
rom[16951] = 12'h  0;
rom[16952] = 12'h  0;
rom[16953] = 12'h  0;
rom[16954] = 12'h  0;
rom[16955] = 12'h  0;
rom[16956] = 12'h  0;
rom[16957] = 12'h  0;
rom[16958] = 12'h  0;
rom[16959] = 12'h  0;
rom[16960] = 12'h  0;
rom[16961] = 12'h  0;
rom[16962] = 12'h  0;
rom[16963] = 12'h  0;
rom[16964] = 12'h100;
rom[16965] = 12'h100;
rom[16966] = 12'h100;
rom[16967] = 12'h100;
rom[16968] = 12'h100;
rom[16969] = 12'h100;
rom[16970] = 12'h200;
rom[16971] = 12'h200;
rom[16972] = 12'h200;
rom[16973] = 12'h300;
rom[16974] = 12'h300;
rom[16975] = 12'h300;
rom[16976] = 12'h300;
rom[16977] = 12'h300;
rom[16978] = 12'h300;
rom[16979] = 12'h300;
rom[16980] = 12'h300;
rom[16981] = 12'h300;
rom[16982] = 12'h300;
rom[16983] = 12'h300;
rom[16984] = 12'h300;
rom[16985] = 12'h300;
rom[16986] = 12'h300;
rom[16987] = 12'h300;
rom[16988] = 12'h300;
rom[16989] = 12'h300;
rom[16990] = 12'h300;
rom[16991] = 12'h200;
rom[16992] = 12'h200;
rom[16993] = 12'h111;
rom[16994] = 12'h211;
rom[16995] = 12'h322;
rom[16996] = 12'h444;
rom[16997] = 12'h766;
rom[16998] = 12'h988;
rom[16999] = 12'haaa;
rom[17000] = 12'hbbb;
rom[17001] = 12'hcbb;
rom[17002] = 12'hcbb;
rom[17003] = 12'hcbb;
rom[17004] = 12'hbbb;
rom[17005] = 12'hbbb;
rom[17006] = 12'hbbb;
rom[17007] = 12'haaa;
rom[17008] = 12'haaa;
rom[17009] = 12'h9aa;
rom[17010] = 12'h999;
rom[17011] = 12'h999;
rom[17012] = 12'h899;
rom[17013] = 12'h899;
rom[17014] = 12'h888;
rom[17015] = 12'h888;
rom[17016] = 12'h888;
rom[17017] = 12'h888;
rom[17018] = 12'h888;
rom[17019] = 12'h888;
rom[17020] = 12'h999;
rom[17021] = 12'h999;
rom[17022] = 12'h999;
rom[17023] = 12'h888;
rom[17024] = 12'h777;
rom[17025] = 12'h777;
rom[17026] = 12'h777;
rom[17027] = 12'h777;
rom[17028] = 12'h888;
rom[17029] = 12'h777;
rom[17030] = 12'h777;
rom[17031] = 12'h777;
rom[17032] = 12'h777;
rom[17033] = 12'h777;
rom[17034] = 12'h666;
rom[17035] = 12'h666;
rom[17036] = 12'h555;
rom[17037] = 12'h555;
rom[17038] = 12'h666;
rom[17039] = 12'h666;
rom[17040] = 12'h666;
rom[17041] = 12'h666;
rom[17042] = 12'h555;
rom[17043] = 12'h555;
rom[17044] = 12'h666;
rom[17045] = 12'h666;
rom[17046] = 12'h666;
rom[17047] = 12'h555;
rom[17048] = 12'h555;
rom[17049] = 12'h444;
rom[17050] = 12'h333;
rom[17051] = 12'h333;
rom[17052] = 12'h222;
rom[17053] = 12'h222;
rom[17054] = 12'h222;
rom[17055] = 12'h222;
rom[17056] = 12'h222;
rom[17057] = 12'h222;
rom[17058] = 12'h111;
rom[17059] = 12'h111;
rom[17060] = 12'h111;
rom[17061] = 12'h111;
rom[17062] = 12'h111;
rom[17063] = 12'h111;
rom[17064] = 12'h111;
rom[17065] = 12'h  0;
rom[17066] = 12'h  0;
rom[17067] = 12'h  0;
rom[17068] = 12'h  0;
rom[17069] = 12'h  0;
rom[17070] = 12'h  0;
rom[17071] = 12'h  0;
rom[17072] = 12'h  0;
rom[17073] = 12'h  0;
rom[17074] = 12'h  0;
rom[17075] = 12'h  0;
rom[17076] = 12'h  0;
rom[17077] = 12'h  0;
rom[17078] = 12'h  0;
rom[17079] = 12'h  0;
rom[17080] = 12'h  0;
rom[17081] = 12'h  0;
rom[17082] = 12'h  0;
rom[17083] = 12'h  0;
rom[17084] = 12'h  0;
rom[17085] = 12'h  0;
rom[17086] = 12'h  0;
rom[17087] = 12'h  0;
rom[17088] = 12'h  0;
rom[17089] = 12'h  0;
rom[17090] = 12'h  0;
rom[17091] = 12'h  0;
rom[17092] = 12'h  0;
rom[17093] = 12'h  0;
rom[17094] = 12'h  0;
rom[17095] = 12'h  0;
rom[17096] = 12'h  0;
rom[17097] = 12'h111;
rom[17098] = 12'h111;
rom[17099] = 12'h111;
rom[17100] = 12'h111;
rom[17101] = 12'h  0;
rom[17102] = 12'h  0;
rom[17103] = 12'h  0;
rom[17104] = 12'h111;
rom[17105] = 12'h111;
rom[17106] = 12'h111;
rom[17107] = 12'h111;
rom[17108] = 12'h222;
rom[17109] = 12'h333;
rom[17110] = 12'h333;
rom[17111] = 12'h333;
rom[17112] = 12'h333;
rom[17113] = 12'h333;
rom[17114] = 12'h333;
rom[17115] = 12'h333;
rom[17116] = 12'h333;
rom[17117] = 12'h333;
rom[17118] = 12'h333;
rom[17119] = 12'h333;
rom[17120] = 12'h333;
rom[17121] = 12'h333;
rom[17122] = 12'h333;
rom[17123] = 12'h333;
rom[17124] = 12'h333;
rom[17125] = 12'h444;
rom[17126] = 12'h444;
rom[17127] = 12'h444;
rom[17128] = 12'h333;
rom[17129] = 12'h222;
rom[17130] = 12'h111;
rom[17131] = 12'h111;
rom[17132] = 12'h111;
rom[17133] = 12'h111;
rom[17134] = 12'h111;
rom[17135] = 12'h111;
rom[17136] = 12'h  0;
rom[17137] = 12'h  0;
rom[17138] = 12'h111;
rom[17139] = 12'h111;
rom[17140] = 12'h111;
rom[17141] = 12'h111;
rom[17142] = 12'h111;
rom[17143] = 12'h111;
rom[17144] = 12'h  0;
rom[17145] = 12'h111;
rom[17146] = 12'h222;
rom[17147] = 12'h333;
rom[17148] = 12'h444;
rom[17149] = 12'h555;
rom[17150] = 12'h555;
rom[17151] = 12'h555;
rom[17152] = 12'h666;
rom[17153] = 12'h666;
rom[17154] = 12'h666;
rom[17155] = 12'h666;
rom[17156] = 12'h555;
rom[17157] = 12'h555;
rom[17158] = 12'h555;
rom[17159] = 12'h555;
rom[17160] = 12'h555;
rom[17161] = 12'h555;
rom[17162] = 12'h555;
rom[17163] = 12'h444;
rom[17164] = 12'h444;
rom[17165] = 12'h444;
rom[17166] = 12'h444;
rom[17167] = 12'h444;
rom[17168] = 12'h444;
rom[17169] = 12'h444;
rom[17170] = 12'h555;
rom[17171] = 12'h555;
rom[17172] = 12'h555;
rom[17173] = 12'h555;
rom[17174] = 12'h666;
rom[17175] = 12'h666;
rom[17176] = 12'h777;
rom[17177] = 12'h777;
rom[17178] = 12'h888;
rom[17179] = 12'h888;
rom[17180] = 12'h888;
rom[17181] = 12'h888;
rom[17182] = 12'h888;
rom[17183] = 12'h888;
rom[17184] = 12'h888;
rom[17185] = 12'h888;
rom[17186] = 12'h888;
rom[17187] = 12'h888;
rom[17188] = 12'h777;
rom[17189] = 12'h777;
rom[17190] = 12'h888;
rom[17191] = 12'h888;
rom[17192] = 12'h888;
rom[17193] = 12'h888;
rom[17194] = 12'h888;
rom[17195] = 12'h999;
rom[17196] = 12'h999;
rom[17197] = 12'haaa;
rom[17198] = 12'haaa;
rom[17199] = 12'haaa;
rom[17200] = 12'h222;
rom[17201] = 12'h222;
rom[17202] = 12'h222;
rom[17203] = 12'h222;
rom[17204] = 12'h222;
rom[17205] = 12'h222;
rom[17206] = 12'h222;
rom[17207] = 12'h222;
rom[17208] = 12'h222;
rom[17209] = 12'h222;
rom[17210] = 12'h222;
rom[17211] = 12'h222;
rom[17212] = 12'h222;
rom[17213] = 12'h222;
rom[17214] = 12'h222;
rom[17215] = 12'h222;
rom[17216] = 12'h222;
rom[17217] = 12'h222;
rom[17218] = 12'h222;
rom[17219] = 12'h333;
rom[17220] = 12'h333;
rom[17221] = 12'h333;
rom[17222] = 12'h333;
rom[17223] = 12'h333;
rom[17224] = 12'h333;
rom[17225] = 12'h444;
rom[17226] = 12'h444;
rom[17227] = 12'h444;
rom[17228] = 12'h444;
rom[17229] = 12'h555;
rom[17230] = 12'h555;
rom[17231] = 12'h555;
rom[17232] = 12'h555;
rom[17233] = 12'h555;
rom[17234] = 12'h555;
rom[17235] = 12'h666;
rom[17236] = 12'h666;
rom[17237] = 12'h666;
rom[17238] = 12'h666;
rom[17239] = 12'h666;
rom[17240] = 12'h666;
rom[17241] = 12'h666;
rom[17242] = 12'h777;
rom[17243] = 12'h777;
rom[17244] = 12'h666;
rom[17245] = 12'h666;
rom[17246] = 12'h666;
rom[17247] = 12'h666;
rom[17248] = 12'h666;
rom[17249] = 12'h555;
rom[17250] = 12'h555;
rom[17251] = 12'h555;
rom[17252] = 12'h555;
rom[17253] = 12'h555;
rom[17254] = 12'h555;
rom[17255] = 12'h555;
rom[17256] = 12'h555;
rom[17257] = 12'h555;
rom[17258] = 12'h555;
rom[17259] = 12'h555;
rom[17260] = 12'h555;
rom[17261] = 12'h555;
rom[17262] = 12'h555;
rom[17263] = 12'h555;
rom[17264] = 12'h555;
rom[17265] = 12'h666;
rom[17266] = 12'h777;
rom[17267] = 12'h777;
rom[17268] = 12'h666;
rom[17269] = 12'h666;
rom[17270] = 12'h666;
rom[17271] = 12'h666;
rom[17272] = 12'h777;
rom[17273] = 12'h777;
rom[17274] = 12'h777;
rom[17275] = 12'h777;
rom[17276] = 12'h777;
rom[17277] = 12'h777;
rom[17278] = 12'h777;
rom[17279] = 12'h777;
rom[17280] = 12'h777;
rom[17281] = 12'h777;
rom[17282] = 12'h666;
rom[17283] = 12'h555;
rom[17284] = 12'h555;
rom[17285] = 12'h444;
rom[17286] = 12'h444;
rom[17287] = 12'h333;
rom[17288] = 12'h333;
rom[17289] = 12'h222;
rom[17290] = 12'h222;
rom[17291] = 12'h222;
rom[17292] = 12'h111;
rom[17293] = 12'h111;
rom[17294] = 12'h111;
rom[17295] = 12'h111;
rom[17296] = 12'h  0;
rom[17297] = 12'h  0;
rom[17298] = 12'h  0;
rom[17299] = 12'h  0;
rom[17300] = 12'h  0;
rom[17301] = 12'h  0;
rom[17302] = 12'h  0;
rom[17303] = 12'h  0;
rom[17304] = 12'h  0;
rom[17305] = 12'h  0;
rom[17306] = 12'h  0;
rom[17307] = 12'h  0;
rom[17308] = 12'h  0;
rom[17309] = 12'h  0;
rom[17310] = 12'h  0;
rom[17311] = 12'h  0;
rom[17312] = 12'h  0;
rom[17313] = 12'h  0;
rom[17314] = 12'h100;
rom[17315] = 12'h100;
rom[17316] = 12'h200;
rom[17317] = 12'h300;
rom[17318] = 12'h510;
rom[17319] = 12'h710;
rom[17320] = 12'h821;
rom[17321] = 12'h921;
rom[17322] = 12'h920;
rom[17323] = 12'h920;
rom[17324] = 12'h920;
rom[17325] = 12'ha20;
rom[17326] = 12'ha20;
rom[17327] = 12'h920;
rom[17328] = 12'h820;
rom[17329] = 12'h710;
rom[17330] = 12'h710;
rom[17331] = 12'h600;
rom[17332] = 12'h600;
rom[17333] = 12'h600;
rom[17334] = 12'h500;
rom[17335] = 12'h500;
rom[17336] = 12'h400;
rom[17337] = 12'h400;
rom[17338] = 12'h300;
rom[17339] = 12'h200;
rom[17340] = 12'h200;
rom[17341] = 12'h100;
rom[17342] = 12'h100;
rom[17343] = 12'h100;
rom[17344] = 12'h  0;
rom[17345] = 12'h  0;
rom[17346] = 12'h  0;
rom[17347] = 12'h  0;
rom[17348] = 12'h  0;
rom[17349] = 12'h  0;
rom[17350] = 12'h  0;
rom[17351] = 12'h  0;
rom[17352] = 12'h  0;
rom[17353] = 12'h  0;
rom[17354] = 12'h  0;
rom[17355] = 12'h  0;
rom[17356] = 12'h  0;
rom[17357] = 12'h  0;
rom[17358] = 12'h  0;
rom[17359] = 12'h  0;
rom[17360] = 12'h  0;
rom[17361] = 12'h  0;
rom[17362] = 12'h  0;
rom[17363] = 12'h  0;
rom[17364] = 12'h100;
rom[17365] = 12'h100;
rom[17366] = 12'h100;
rom[17367] = 12'h100;
rom[17368] = 12'h100;
rom[17369] = 12'h200;
rom[17370] = 12'h200;
rom[17371] = 12'h200;
rom[17372] = 12'h300;
rom[17373] = 12'h300;
rom[17374] = 12'h300;
rom[17375] = 12'h300;
rom[17376] = 12'h300;
rom[17377] = 12'h300;
rom[17378] = 12'h300;
rom[17379] = 12'h300;
rom[17380] = 12'h300;
rom[17381] = 12'h300;
rom[17382] = 12'h300;
rom[17383] = 12'h200;
rom[17384] = 12'h200;
rom[17385] = 12'h200;
rom[17386] = 12'h200;
rom[17387] = 12'h200;
rom[17388] = 12'h200;
rom[17389] = 12'h200;
rom[17390] = 12'h200;
rom[17391] = 12'h200;
rom[17392] = 12'h100;
rom[17393] = 12'h100;
rom[17394] = 12'h111;
rom[17395] = 12'h212;
rom[17396] = 12'h333;
rom[17397] = 12'h555;
rom[17398] = 12'h877;
rom[17399] = 12'ha99;
rom[17400] = 12'hbaa;
rom[17401] = 12'hbbb;
rom[17402] = 12'hcbb;
rom[17403] = 12'hcbb;
rom[17404] = 12'hbbb;
rom[17405] = 12'hbbb;
rom[17406] = 12'hbbb;
rom[17407] = 12'hbaa;
rom[17408] = 12'haaa;
rom[17409] = 12'haaa;
rom[17410] = 12'h9a9;
rom[17411] = 12'h999;
rom[17412] = 12'h999;
rom[17413] = 12'h899;
rom[17414] = 12'h898;
rom[17415] = 12'h888;
rom[17416] = 12'h888;
rom[17417] = 12'h888;
rom[17418] = 12'h888;
rom[17419] = 12'h888;
rom[17420] = 12'h999;
rom[17421] = 12'h888;
rom[17422] = 12'h888;
rom[17423] = 12'h888;
rom[17424] = 12'h888;
rom[17425] = 12'h777;
rom[17426] = 12'h777;
rom[17427] = 12'h777;
rom[17428] = 12'h777;
rom[17429] = 12'h777;
rom[17430] = 12'h777;
rom[17431] = 12'h777;
rom[17432] = 12'h777;
rom[17433] = 12'h777;
rom[17434] = 12'h666;
rom[17435] = 12'h666;
rom[17436] = 12'h666;
rom[17437] = 12'h666;
rom[17438] = 12'h666;
rom[17439] = 12'h666;
rom[17440] = 12'h666;
rom[17441] = 12'h666;
rom[17442] = 12'h666;
rom[17443] = 12'h666;
rom[17444] = 12'h666;
rom[17445] = 12'h666;
rom[17446] = 12'h555;
rom[17447] = 12'h555;
rom[17448] = 12'h444;
rom[17449] = 12'h333;
rom[17450] = 12'h333;
rom[17451] = 12'h333;
rom[17452] = 12'h333;
rom[17453] = 12'h333;
rom[17454] = 12'h222;
rom[17455] = 12'h222;
rom[17456] = 12'h222;
rom[17457] = 12'h222;
rom[17458] = 12'h111;
rom[17459] = 12'h111;
rom[17460] = 12'h111;
rom[17461] = 12'h111;
rom[17462] = 12'h111;
rom[17463] = 12'h111;
rom[17464] = 12'h111;
rom[17465] = 12'h  0;
rom[17466] = 12'h  0;
rom[17467] = 12'h  0;
rom[17468] = 12'h  0;
rom[17469] = 12'h  0;
rom[17470] = 12'h  0;
rom[17471] = 12'h  0;
rom[17472] = 12'h  0;
rom[17473] = 12'h  0;
rom[17474] = 12'h  0;
rom[17475] = 12'h  0;
rom[17476] = 12'h  0;
rom[17477] = 12'h  0;
rom[17478] = 12'h  0;
rom[17479] = 12'h  0;
rom[17480] = 12'h  0;
rom[17481] = 12'h  0;
rom[17482] = 12'h  0;
rom[17483] = 12'h  0;
rom[17484] = 12'h  0;
rom[17485] = 12'h  0;
rom[17486] = 12'h  0;
rom[17487] = 12'h  0;
rom[17488] = 12'h  0;
rom[17489] = 12'h  0;
rom[17490] = 12'h  0;
rom[17491] = 12'h  0;
rom[17492] = 12'h  0;
rom[17493] = 12'h  0;
rom[17494] = 12'h  0;
rom[17495] = 12'h  0;
rom[17496] = 12'h111;
rom[17497] = 12'h111;
rom[17498] = 12'h111;
rom[17499] = 12'h111;
rom[17500] = 12'h111;
rom[17501] = 12'h  0;
rom[17502] = 12'h  0;
rom[17503] = 12'h111;
rom[17504] = 12'h111;
rom[17505] = 12'h111;
rom[17506] = 12'h111;
rom[17507] = 12'h222;
rom[17508] = 12'h222;
rom[17509] = 12'h333;
rom[17510] = 12'h333;
rom[17511] = 12'h333;
rom[17512] = 12'h333;
rom[17513] = 12'h333;
rom[17514] = 12'h333;
rom[17515] = 12'h333;
rom[17516] = 12'h333;
rom[17517] = 12'h444;
rom[17518] = 12'h444;
rom[17519] = 12'h333;
rom[17520] = 12'h333;
rom[17521] = 12'h333;
rom[17522] = 12'h333;
rom[17523] = 12'h333;
rom[17524] = 12'h333;
rom[17525] = 12'h444;
rom[17526] = 12'h444;
rom[17527] = 12'h444;
rom[17528] = 12'h333;
rom[17529] = 12'h222;
rom[17530] = 12'h222;
rom[17531] = 12'h111;
rom[17532] = 12'h111;
rom[17533] = 12'h111;
rom[17534] = 12'h111;
rom[17535] = 12'h111;
rom[17536] = 12'h111;
rom[17537] = 12'h111;
rom[17538] = 12'h111;
rom[17539] = 12'h111;
rom[17540] = 12'h111;
rom[17541] = 12'h111;
rom[17542] = 12'h111;
rom[17543] = 12'h111;
rom[17544] = 12'h222;
rom[17545] = 12'h222;
rom[17546] = 12'h333;
rom[17547] = 12'h444;
rom[17548] = 12'h444;
rom[17549] = 12'h555;
rom[17550] = 12'h555;
rom[17551] = 12'h555;
rom[17552] = 12'h666;
rom[17553] = 12'h666;
rom[17554] = 12'h555;
rom[17555] = 12'h555;
rom[17556] = 12'h555;
rom[17557] = 12'h555;
rom[17558] = 12'h555;
rom[17559] = 12'h555;
rom[17560] = 12'h555;
rom[17561] = 12'h555;
rom[17562] = 12'h444;
rom[17563] = 12'h444;
rom[17564] = 12'h444;
rom[17565] = 12'h444;
rom[17566] = 12'h444;
rom[17567] = 12'h444;
rom[17568] = 12'h444;
rom[17569] = 12'h444;
rom[17570] = 12'h555;
rom[17571] = 12'h555;
rom[17572] = 12'h555;
rom[17573] = 12'h555;
rom[17574] = 12'h555;
rom[17575] = 12'h555;
rom[17576] = 12'h555;
rom[17577] = 12'h555;
rom[17578] = 12'h666;
rom[17579] = 12'h777;
rom[17580] = 12'h777;
rom[17581] = 12'h888;
rom[17582] = 12'h888;
rom[17583] = 12'h888;
rom[17584] = 12'h888;
rom[17585] = 12'h888;
rom[17586] = 12'h888;
rom[17587] = 12'h888;
rom[17588] = 12'h888;
rom[17589] = 12'h777;
rom[17590] = 12'h777;
rom[17591] = 12'h777;
rom[17592] = 12'h888;
rom[17593] = 12'h888;
rom[17594] = 12'h888;
rom[17595] = 12'h999;
rom[17596] = 12'haaa;
rom[17597] = 12'haaa;
rom[17598] = 12'haaa;
rom[17599] = 12'haaa;
rom[17600] = 12'h222;
rom[17601] = 12'h222;
rom[17602] = 12'h222;
rom[17603] = 12'h222;
rom[17604] = 12'h222;
rom[17605] = 12'h222;
rom[17606] = 12'h222;
rom[17607] = 12'h222;
rom[17608] = 12'h222;
rom[17609] = 12'h222;
rom[17610] = 12'h222;
rom[17611] = 12'h222;
rom[17612] = 12'h222;
rom[17613] = 12'h222;
rom[17614] = 12'h333;
rom[17615] = 12'h333;
rom[17616] = 12'h333;
rom[17617] = 12'h333;
rom[17618] = 12'h333;
rom[17619] = 12'h333;
rom[17620] = 12'h333;
rom[17621] = 12'h444;
rom[17622] = 12'h444;
rom[17623] = 12'h444;
rom[17624] = 12'h444;
rom[17625] = 12'h444;
rom[17626] = 12'h444;
rom[17627] = 12'h444;
rom[17628] = 12'h555;
rom[17629] = 12'h555;
rom[17630] = 12'h555;
rom[17631] = 12'h555;
rom[17632] = 12'h666;
rom[17633] = 12'h666;
rom[17634] = 12'h666;
rom[17635] = 12'h666;
rom[17636] = 12'h666;
rom[17637] = 12'h666;
rom[17638] = 12'h666;
rom[17639] = 12'h666;
rom[17640] = 12'h666;
rom[17641] = 12'h666;
rom[17642] = 12'h666;
rom[17643] = 12'h666;
rom[17644] = 12'h666;
rom[17645] = 12'h666;
rom[17646] = 12'h666;
rom[17647] = 12'h666;
rom[17648] = 12'h555;
rom[17649] = 12'h555;
rom[17650] = 12'h555;
rom[17651] = 12'h555;
rom[17652] = 12'h555;
rom[17653] = 12'h555;
rom[17654] = 12'h555;
rom[17655] = 12'h555;
rom[17656] = 12'h555;
rom[17657] = 12'h555;
rom[17658] = 12'h555;
rom[17659] = 12'h555;
rom[17660] = 12'h555;
rom[17661] = 12'h555;
rom[17662] = 12'h555;
rom[17663] = 12'h555;
rom[17664] = 12'h555;
rom[17665] = 12'h555;
rom[17666] = 12'h666;
rom[17667] = 12'h777;
rom[17668] = 12'h777;
rom[17669] = 12'h777;
rom[17670] = 12'h777;
rom[17671] = 12'h666;
rom[17672] = 12'h666;
rom[17673] = 12'h777;
rom[17674] = 12'h777;
rom[17675] = 12'h777;
rom[17676] = 12'h777;
rom[17677] = 12'h777;
rom[17678] = 12'h777;
rom[17679] = 12'h777;
rom[17680] = 12'h777;
rom[17681] = 12'h777;
rom[17682] = 12'h666;
rom[17683] = 12'h666;
rom[17684] = 12'h555;
rom[17685] = 12'h444;
rom[17686] = 12'h444;
rom[17687] = 12'h333;
rom[17688] = 12'h333;
rom[17689] = 12'h222;
rom[17690] = 12'h222;
rom[17691] = 12'h222;
rom[17692] = 12'h111;
rom[17693] = 12'h111;
rom[17694] = 12'h111;
rom[17695] = 12'h111;
rom[17696] = 12'h  0;
rom[17697] = 12'h  0;
rom[17698] = 12'h  0;
rom[17699] = 12'h  0;
rom[17700] = 12'h  0;
rom[17701] = 12'h  0;
rom[17702] = 12'h  0;
rom[17703] = 12'h  0;
rom[17704] = 12'h  0;
rom[17705] = 12'h  0;
rom[17706] = 12'h  0;
rom[17707] = 12'h  0;
rom[17708] = 12'h  0;
rom[17709] = 12'h  0;
rom[17710] = 12'h  0;
rom[17711] = 12'h  0;
rom[17712] = 12'h  0;
rom[17713] = 12'h  0;
rom[17714] = 12'h100;
rom[17715] = 12'h100;
rom[17716] = 12'h200;
rom[17717] = 12'h300;
rom[17718] = 12'h500;
rom[17719] = 12'h710;
rom[17720] = 12'h821;
rom[17721] = 12'h921;
rom[17722] = 12'h920;
rom[17723] = 12'h920;
rom[17724] = 12'ha20;
rom[17725] = 12'ha20;
rom[17726] = 12'ha20;
rom[17727] = 12'h920;
rom[17728] = 12'h920;
rom[17729] = 12'h810;
rom[17730] = 12'h710;
rom[17731] = 12'h710;
rom[17732] = 12'h610;
rom[17733] = 12'h610;
rom[17734] = 12'h600;
rom[17735] = 12'h500;
rom[17736] = 12'h400;
rom[17737] = 12'h400;
rom[17738] = 12'h300;
rom[17739] = 12'h200;
rom[17740] = 12'h200;
rom[17741] = 12'h100;
rom[17742] = 12'h100;
rom[17743] = 12'h100;
rom[17744] = 12'h100;
rom[17745] = 12'h  0;
rom[17746] = 12'h  0;
rom[17747] = 12'h  0;
rom[17748] = 12'h  0;
rom[17749] = 12'h  0;
rom[17750] = 12'h  0;
rom[17751] = 12'h  0;
rom[17752] = 12'h  0;
rom[17753] = 12'h  0;
rom[17754] = 12'h  0;
rom[17755] = 12'h  0;
rom[17756] = 12'h  0;
rom[17757] = 12'h  0;
rom[17758] = 12'h  0;
rom[17759] = 12'h  0;
rom[17760] = 12'h  0;
rom[17761] = 12'h100;
rom[17762] = 12'h100;
rom[17763] = 12'h100;
rom[17764] = 12'h100;
rom[17765] = 12'h100;
rom[17766] = 12'h100;
rom[17767] = 12'h100;
rom[17768] = 12'h200;
rom[17769] = 12'h200;
rom[17770] = 12'h200;
rom[17771] = 12'h200;
rom[17772] = 12'h300;
rom[17773] = 12'h300;
rom[17774] = 12'h300;
rom[17775] = 12'h300;
rom[17776] = 12'h300;
rom[17777] = 12'h300;
rom[17778] = 12'h300;
rom[17779] = 12'h300;
rom[17780] = 12'h300;
rom[17781] = 12'h300;
rom[17782] = 12'h200;
rom[17783] = 12'h200;
rom[17784] = 12'h200;
rom[17785] = 12'h200;
rom[17786] = 12'h200;
rom[17787] = 12'h200;
rom[17788] = 12'h200;
rom[17789] = 12'h200;
rom[17790] = 12'h200;
rom[17791] = 12'h200;
rom[17792] = 12'h100;
rom[17793] = 12'h100;
rom[17794] = 12'h101;
rom[17795] = 12'h211;
rom[17796] = 12'h322;
rom[17797] = 12'h444;
rom[17798] = 12'h766;
rom[17799] = 12'h988;
rom[17800] = 12'ha9a;
rom[17801] = 12'hbbb;
rom[17802] = 12'hcbb;
rom[17803] = 12'hcbb;
rom[17804] = 12'hbbb;
rom[17805] = 12'hbbb;
rom[17806] = 12'hbbb;
rom[17807] = 12'hbbb;
rom[17808] = 12'haba;
rom[17809] = 12'haaa;
rom[17810] = 12'h9aa;
rom[17811] = 12'h999;
rom[17812] = 12'h999;
rom[17813] = 12'h899;
rom[17814] = 12'h899;
rom[17815] = 12'h888;
rom[17816] = 12'h888;
rom[17817] = 12'h888;
rom[17818] = 12'h888;
rom[17819] = 12'h888;
rom[17820] = 12'h888;
rom[17821] = 12'h888;
rom[17822] = 12'h888;
rom[17823] = 12'h888;
rom[17824] = 12'h888;
rom[17825] = 12'h888;
rom[17826] = 12'h777;
rom[17827] = 12'h777;
rom[17828] = 12'h777;
rom[17829] = 12'h777;
rom[17830] = 12'h777;
rom[17831] = 12'h777;
rom[17832] = 12'h666;
rom[17833] = 12'h666;
rom[17834] = 12'h666;
rom[17835] = 12'h666;
rom[17836] = 12'h666;
rom[17837] = 12'h666;
rom[17838] = 12'h666;
rom[17839] = 12'h666;
rom[17840] = 12'h666;
rom[17841] = 12'h666;
rom[17842] = 12'h777;
rom[17843] = 12'h777;
rom[17844] = 12'h666;
rom[17845] = 12'h555;
rom[17846] = 12'h555;
rom[17847] = 12'h444;
rom[17848] = 12'h333;
rom[17849] = 12'h333;
rom[17850] = 12'h333;
rom[17851] = 12'h333;
rom[17852] = 12'h333;
rom[17853] = 12'h333;
rom[17854] = 12'h222;
rom[17855] = 12'h222;
rom[17856] = 12'h222;
rom[17857] = 12'h222;
rom[17858] = 12'h111;
rom[17859] = 12'h111;
rom[17860] = 12'h111;
rom[17861] = 12'h111;
rom[17862] = 12'h111;
rom[17863] = 12'h111;
rom[17864] = 12'h111;
rom[17865] = 12'h  0;
rom[17866] = 12'h  0;
rom[17867] = 12'h  0;
rom[17868] = 12'h  0;
rom[17869] = 12'h  0;
rom[17870] = 12'h  0;
rom[17871] = 12'h  0;
rom[17872] = 12'h  0;
rom[17873] = 12'h  0;
rom[17874] = 12'h  0;
rom[17875] = 12'h  0;
rom[17876] = 12'h  0;
rom[17877] = 12'h  0;
rom[17878] = 12'h  0;
rom[17879] = 12'h  0;
rom[17880] = 12'h  0;
rom[17881] = 12'h  0;
rom[17882] = 12'h  0;
rom[17883] = 12'h  0;
rom[17884] = 12'h  0;
rom[17885] = 12'h  0;
rom[17886] = 12'h  0;
rom[17887] = 12'h  0;
rom[17888] = 12'h  0;
rom[17889] = 12'h  0;
rom[17890] = 12'h  0;
rom[17891] = 12'h  0;
rom[17892] = 12'h  0;
rom[17893] = 12'h  0;
rom[17894] = 12'h  0;
rom[17895] = 12'h  0;
rom[17896] = 12'h111;
rom[17897] = 12'h111;
rom[17898] = 12'h111;
rom[17899] = 12'h111;
rom[17900] = 12'h111;
rom[17901] = 12'h111;
rom[17902] = 12'h111;
rom[17903] = 12'h111;
rom[17904] = 12'h111;
rom[17905] = 12'h111;
rom[17906] = 12'h111;
rom[17907] = 12'h222;
rom[17908] = 12'h333;
rom[17909] = 12'h333;
rom[17910] = 12'h333;
rom[17911] = 12'h333;
rom[17912] = 12'h333;
rom[17913] = 12'h333;
rom[17914] = 12'h333;
rom[17915] = 12'h333;
rom[17916] = 12'h333;
rom[17917] = 12'h444;
rom[17918] = 12'h444;
rom[17919] = 12'h333;
rom[17920] = 12'h333;
rom[17921] = 12'h333;
rom[17922] = 12'h333;
rom[17923] = 12'h333;
rom[17924] = 12'h333;
rom[17925] = 12'h444;
rom[17926] = 12'h444;
rom[17927] = 12'h444;
rom[17928] = 12'h333;
rom[17929] = 12'h333;
rom[17930] = 12'h222;
rom[17931] = 12'h222;
rom[17932] = 12'h111;
rom[17933] = 12'h111;
rom[17934] = 12'h111;
rom[17935] = 12'h111;
rom[17936] = 12'h111;
rom[17937] = 12'h111;
rom[17938] = 12'h111;
rom[17939] = 12'h111;
rom[17940] = 12'h111;
rom[17941] = 12'h111;
rom[17942] = 12'h111;
rom[17943] = 12'h222;
rom[17944] = 12'h333;
rom[17945] = 12'h333;
rom[17946] = 12'h444;
rom[17947] = 12'h444;
rom[17948] = 12'h555;
rom[17949] = 12'h555;
rom[17950] = 12'h555;
rom[17951] = 12'h666;
rom[17952] = 12'h555;
rom[17953] = 12'h555;
rom[17954] = 12'h555;
rom[17955] = 12'h555;
rom[17956] = 12'h555;
rom[17957] = 12'h555;
rom[17958] = 12'h555;
rom[17959] = 12'h555;
rom[17960] = 12'h555;
rom[17961] = 12'h555;
rom[17962] = 12'h555;
rom[17963] = 12'h444;
rom[17964] = 12'h444;
rom[17965] = 12'h444;
rom[17966] = 12'h555;
rom[17967] = 12'h555;
rom[17968] = 12'h555;
rom[17969] = 12'h555;
rom[17970] = 12'h555;
rom[17971] = 12'h555;
rom[17972] = 12'h555;
rom[17973] = 12'h555;
rom[17974] = 12'h555;
rom[17975] = 12'h555;
rom[17976] = 12'h555;
rom[17977] = 12'h666;
rom[17978] = 12'h666;
rom[17979] = 12'h666;
rom[17980] = 12'h666;
rom[17981] = 12'h777;
rom[17982] = 12'h777;
rom[17983] = 12'h777;
rom[17984] = 12'h888;
rom[17985] = 12'h888;
rom[17986] = 12'h888;
rom[17987] = 12'h888;
rom[17988] = 12'h888;
rom[17989] = 12'h888;
rom[17990] = 12'h777;
rom[17991] = 12'h777;
rom[17992] = 12'h888;
rom[17993] = 12'h888;
rom[17994] = 12'h888;
rom[17995] = 12'h999;
rom[17996] = 12'haaa;
rom[17997] = 12'haaa;
rom[17998] = 12'haaa;
rom[17999] = 12'haaa;
rom[18000] = 12'h222;
rom[18001] = 12'h222;
rom[18002] = 12'h222;
rom[18003] = 12'h222;
rom[18004] = 12'h222;
rom[18005] = 12'h222;
rom[18006] = 12'h222;
rom[18007] = 12'h222;
rom[18008] = 12'h222;
rom[18009] = 12'h222;
rom[18010] = 12'h222;
rom[18011] = 12'h222;
rom[18012] = 12'h333;
rom[18013] = 12'h333;
rom[18014] = 12'h333;
rom[18015] = 12'h333;
rom[18016] = 12'h333;
rom[18017] = 12'h333;
rom[18018] = 12'h444;
rom[18019] = 12'h444;
rom[18020] = 12'h444;
rom[18021] = 12'h444;
rom[18022] = 12'h444;
rom[18023] = 12'h444;
rom[18024] = 12'h444;
rom[18025] = 12'h555;
rom[18026] = 12'h555;
rom[18027] = 12'h555;
rom[18028] = 12'h555;
rom[18029] = 12'h666;
rom[18030] = 12'h666;
rom[18031] = 12'h666;
rom[18032] = 12'h666;
rom[18033] = 12'h666;
rom[18034] = 12'h666;
rom[18035] = 12'h666;
rom[18036] = 12'h777;
rom[18037] = 12'h777;
rom[18038] = 12'h777;
rom[18039] = 12'h777;
rom[18040] = 12'h666;
rom[18041] = 12'h666;
rom[18042] = 12'h666;
rom[18043] = 12'h666;
rom[18044] = 12'h666;
rom[18045] = 12'h666;
rom[18046] = 12'h555;
rom[18047] = 12'h555;
rom[18048] = 12'h555;
rom[18049] = 12'h555;
rom[18050] = 12'h555;
rom[18051] = 12'h555;
rom[18052] = 12'h555;
rom[18053] = 12'h555;
rom[18054] = 12'h555;
rom[18055] = 12'h555;
rom[18056] = 12'h555;
rom[18057] = 12'h555;
rom[18058] = 12'h555;
rom[18059] = 12'h555;
rom[18060] = 12'h555;
rom[18061] = 12'h555;
rom[18062] = 12'h555;
rom[18063] = 12'h555;
rom[18064] = 12'h555;
rom[18065] = 12'h555;
rom[18066] = 12'h555;
rom[18067] = 12'h666;
rom[18068] = 12'h666;
rom[18069] = 12'h777;
rom[18070] = 12'h777;
rom[18071] = 12'h777;
rom[18072] = 12'h666;
rom[18073] = 12'h777;
rom[18074] = 12'h777;
rom[18075] = 12'h777;
rom[18076] = 12'h777;
rom[18077] = 12'h777;
rom[18078] = 12'h777;
rom[18079] = 12'h777;
rom[18080] = 12'h777;
rom[18081] = 12'h777;
rom[18082] = 12'h777;
rom[18083] = 12'h666;
rom[18084] = 12'h555;
rom[18085] = 12'h555;
rom[18086] = 12'h444;
rom[18087] = 12'h333;
rom[18088] = 12'h333;
rom[18089] = 12'h222;
rom[18090] = 12'h222;
rom[18091] = 12'h222;
rom[18092] = 12'h111;
rom[18093] = 12'h111;
rom[18094] = 12'h111;
rom[18095] = 12'h111;
rom[18096] = 12'h  0;
rom[18097] = 12'h  0;
rom[18098] = 12'h  0;
rom[18099] = 12'h  0;
rom[18100] = 12'h  0;
rom[18101] = 12'h  0;
rom[18102] = 12'h  0;
rom[18103] = 12'h  0;
rom[18104] = 12'h  0;
rom[18105] = 12'h  0;
rom[18106] = 12'h  0;
rom[18107] = 12'h  0;
rom[18108] = 12'h  0;
rom[18109] = 12'h  0;
rom[18110] = 12'h  0;
rom[18111] = 12'h  0;
rom[18112] = 12'h  0;
rom[18113] = 12'h  0;
rom[18114] = 12'h100;
rom[18115] = 12'h200;
rom[18116] = 12'h200;
rom[18117] = 12'h300;
rom[18118] = 12'h500;
rom[18119] = 12'h710;
rom[18120] = 12'h821;
rom[18121] = 12'h921;
rom[18122] = 12'ha31;
rom[18123] = 12'ha30;
rom[18124] = 12'ha30;
rom[18125] = 12'ha20;
rom[18126] = 12'ha30;
rom[18127] = 12'ha20;
rom[18128] = 12'h921;
rom[18129] = 12'h820;
rom[18130] = 12'h710;
rom[18131] = 12'h710;
rom[18132] = 12'h710;
rom[18133] = 12'h610;
rom[18134] = 12'h610;
rom[18135] = 12'h500;
rom[18136] = 12'h400;
rom[18137] = 12'h400;
rom[18138] = 12'h300;
rom[18139] = 12'h200;
rom[18140] = 12'h200;
rom[18141] = 12'h100;
rom[18142] = 12'h100;
rom[18143] = 12'h100;
rom[18144] = 12'h100;
rom[18145] = 12'h100;
rom[18146] = 12'h  0;
rom[18147] = 12'h  0;
rom[18148] = 12'h  0;
rom[18149] = 12'h  0;
rom[18150] = 12'h  0;
rom[18151] = 12'h  0;
rom[18152] = 12'h  0;
rom[18153] = 12'h  0;
rom[18154] = 12'h  0;
rom[18155] = 12'h  0;
rom[18156] = 12'h  0;
rom[18157] = 12'h  0;
rom[18158] = 12'h  0;
rom[18159] = 12'h  0;
rom[18160] = 12'h  0;
rom[18161] = 12'h100;
rom[18162] = 12'h100;
rom[18163] = 12'h100;
rom[18164] = 12'h100;
rom[18165] = 12'h100;
rom[18166] = 12'h100;
rom[18167] = 12'h100;
rom[18168] = 12'h200;
rom[18169] = 12'h200;
rom[18170] = 12'h200;
rom[18171] = 12'h300;
rom[18172] = 12'h300;
rom[18173] = 12'h300;
rom[18174] = 12'h300;
rom[18175] = 12'h300;
rom[18176] = 12'h300;
rom[18177] = 12'h300;
rom[18178] = 12'h300;
rom[18179] = 12'h300;
rom[18180] = 12'h300;
rom[18181] = 12'h300;
rom[18182] = 12'h200;
rom[18183] = 12'h200;
rom[18184] = 12'h200;
rom[18185] = 12'h200;
rom[18186] = 12'h200;
rom[18187] = 12'h200;
rom[18188] = 12'h200;
rom[18189] = 12'h200;
rom[18190] = 12'h200;
rom[18191] = 12'h200;
rom[18192] = 12'h100;
rom[18193] = 12'h100;
rom[18194] = 12'h100;
rom[18195] = 12'h211;
rom[18196] = 12'h322;
rom[18197] = 12'h433;
rom[18198] = 12'h655;
rom[18199] = 12'h877;
rom[18200] = 12'h999;
rom[18201] = 12'haaa;
rom[18202] = 12'hcbb;
rom[18203] = 12'hcbc;
rom[18204] = 12'hcbb;
rom[18205] = 12'hbbb;
rom[18206] = 12'hbbb;
rom[18207] = 12'hbbb;
rom[18208] = 12'habb;
rom[18209] = 12'haaa;
rom[18210] = 12'h9aa;
rom[18211] = 12'h999;
rom[18212] = 12'h999;
rom[18213] = 12'h999;
rom[18214] = 12'h899;
rom[18215] = 12'h888;
rom[18216] = 12'h888;
rom[18217] = 12'h888;
rom[18218] = 12'h888;
rom[18219] = 12'h888;
rom[18220] = 12'h888;
rom[18221] = 12'h888;
rom[18222] = 12'h888;
rom[18223] = 12'h877;
rom[18224] = 12'h888;
rom[18225] = 12'h888;
rom[18226] = 12'h888;
rom[18227] = 12'h888;
rom[18228] = 12'h888;
rom[18229] = 12'h888;
rom[18230] = 12'h777;
rom[18231] = 12'h777;
rom[18232] = 12'h666;
rom[18233] = 12'h666;
rom[18234] = 12'h666;
rom[18235] = 12'h666;
rom[18236] = 12'h777;
rom[18237] = 12'h777;
rom[18238] = 12'h777;
rom[18239] = 12'h666;
rom[18240] = 12'h777;
rom[18241] = 12'h777;
rom[18242] = 12'h777;
rom[18243] = 12'h666;
rom[18244] = 12'h555;
rom[18245] = 12'h444;
rom[18246] = 12'h444;
rom[18247] = 12'h444;
rom[18248] = 12'h333;
rom[18249] = 12'h333;
rom[18250] = 12'h333;
rom[18251] = 12'h333;
rom[18252] = 12'h333;
rom[18253] = 12'h333;
rom[18254] = 12'h222;
rom[18255] = 12'h222;
rom[18256] = 12'h222;
rom[18257] = 12'h222;
rom[18258] = 12'h111;
rom[18259] = 12'h111;
rom[18260] = 12'h111;
rom[18261] = 12'h111;
rom[18262] = 12'h111;
rom[18263] = 12'h111;
rom[18264] = 12'h  0;
rom[18265] = 12'h  0;
rom[18266] = 12'h  0;
rom[18267] = 12'h  0;
rom[18268] = 12'h  0;
rom[18269] = 12'h  0;
rom[18270] = 12'h  0;
rom[18271] = 12'h  0;
rom[18272] = 12'h  0;
rom[18273] = 12'h  0;
rom[18274] = 12'h  0;
rom[18275] = 12'h  0;
rom[18276] = 12'h  0;
rom[18277] = 12'h  0;
rom[18278] = 12'h  0;
rom[18279] = 12'h  0;
rom[18280] = 12'h  0;
rom[18281] = 12'h  0;
rom[18282] = 12'h  0;
rom[18283] = 12'h  0;
rom[18284] = 12'h  0;
rom[18285] = 12'h  0;
rom[18286] = 12'h  0;
rom[18287] = 12'h  0;
rom[18288] = 12'h  0;
rom[18289] = 12'h  0;
rom[18290] = 12'h  0;
rom[18291] = 12'h  0;
rom[18292] = 12'h  0;
rom[18293] = 12'h  0;
rom[18294] = 12'h  0;
rom[18295] = 12'h  0;
rom[18296] = 12'h111;
rom[18297] = 12'h111;
rom[18298] = 12'h111;
rom[18299] = 12'h111;
rom[18300] = 12'h111;
rom[18301] = 12'h111;
rom[18302] = 12'h111;
rom[18303] = 12'h111;
rom[18304] = 12'h111;
rom[18305] = 12'h111;
rom[18306] = 12'h111;
rom[18307] = 12'h222;
rom[18308] = 12'h333;
rom[18309] = 12'h333;
rom[18310] = 12'h333;
rom[18311] = 12'h333;
rom[18312] = 12'h333;
rom[18313] = 12'h333;
rom[18314] = 12'h333;
rom[18315] = 12'h333;
rom[18316] = 12'h333;
rom[18317] = 12'h444;
rom[18318] = 12'h333;
rom[18319] = 12'h333;
rom[18320] = 12'h333;
rom[18321] = 12'h333;
rom[18322] = 12'h333;
rom[18323] = 12'h333;
rom[18324] = 12'h333;
rom[18325] = 12'h444;
rom[18326] = 12'h444;
rom[18327] = 12'h444;
rom[18328] = 12'h333;
rom[18329] = 12'h333;
rom[18330] = 12'h222;
rom[18331] = 12'h222;
rom[18332] = 12'h111;
rom[18333] = 12'h111;
rom[18334] = 12'h111;
rom[18335] = 12'h111;
rom[18336] = 12'h111;
rom[18337] = 12'h111;
rom[18338] = 12'h111;
rom[18339] = 12'h111;
rom[18340] = 12'h222;
rom[18341] = 12'h222;
rom[18342] = 12'h222;
rom[18343] = 12'h333;
rom[18344] = 12'h444;
rom[18345] = 12'h444;
rom[18346] = 12'h444;
rom[18347] = 12'h555;
rom[18348] = 12'h555;
rom[18349] = 12'h555;
rom[18350] = 12'h555;
rom[18351] = 12'h666;
rom[18352] = 12'h666;
rom[18353] = 12'h666;
rom[18354] = 12'h555;
rom[18355] = 12'h555;
rom[18356] = 12'h555;
rom[18357] = 12'h555;
rom[18358] = 12'h555;
rom[18359] = 12'h555;
rom[18360] = 12'h555;
rom[18361] = 12'h555;
rom[18362] = 12'h555;
rom[18363] = 12'h444;
rom[18364] = 12'h444;
rom[18365] = 12'h444;
rom[18366] = 12'h444;
rom[18367] = 12'h444;
rom[18368] = 12'h444;
rom[18369] = 12'h555;
rom[18370] = 12'h555;
rom[18371] = 12'h555;
rom[18372] = 12'h555;
rom[18373] = 12'h555;
rom[18374] = 12'h555;
rom[18375] = 12'h555;
rom[18376] = 12'h666;
rom[18377] = 12'h666;
rom[18378] = 12'h555;
rom[18379] = 12'h666;
rom[18380] = 12'h666;
rom[18381] = 12'h666;
rom[18382] = 12'h666;
rom[18383] = 12'h666;
rom[18384] = 12'h777;
rom[18385] = 12'h888;
rom[18386] = 12'h888;
rom[18387] = 12'h888;
rom[18388] = 12'h888;
rom[18389] = 12'h888;
rom[18390] = 12'h888;
rom[18391] = 12'h888;
rom[18392] = 12'h888;
rom[18393] = 12'h888;
rom[18394] = 12'h888;
rom[18395] = 12'h999;
rom[18396] = 12'haaa;
rom[18397] = 12'haaa;
rom[18398] = 12'haaa;
rom[18399] = 12'haaa;
rom[18400] = 12'h333;
rom[18401] = 12'h333;
rom[18402] = 12'h333;
rom[18403] = 12'h333;
rom[18404] = 12'h333;
rom[18405] = 12'h333;
rom[18406] = 12'h333;
rom[18407] = 12'h333;
rom[18408] = 12'h333;
rom[18409] = 12'h333;
rom[18410] = 12'h333;
rom[18411] = 12'h333;
rom[18412] = 12'h333;
rom[18413] = 12'h333;
rom[18414] = 12'h333;
rom[18415] = 12'h333;
rom[18416] = 12'h444;
rom[18417] = 12'h444;
rom[18418] = 12'h444;
rom[18419] = 12'h444;
rom[18420] = 12'h555;
rom[18421] = 12'h555;
rom[18422] = 12'h555;
rom[18423] = 12'h555;
rom[18424] = 12'h555;
rom[18425] = 12'h555;
rom[18426] = 12'h666;
rom[18427] = 12'h666;
rom[18428] = 12'h666;
rom[18429] = 12'h666;
rom[18430] = 12'h666;
rom[18431] = 12'h666;
rom[18432] = 12'h666;
rom[18433] = 12'h666;
rom[18434] = 12'h777;
rom[18435] = 12'h777;
rom[18436] = 12'h777;
rom[18437] = 12'h777;
rom[18438] = 12'h777;
rom[18439] = 12'h777;
rom[18440] = 12'h777;
rom[18441] = 12'h777;
rom[18442] = 12'h666;
rom[18443] = 12'h666;
rom[18444] = 12'h666;
rom[18445] = 12'h666;
rom[18446] = 12'h555;
rom[18447] = 12'h555;
rom[18448] = 12'h555;
rom[18449] = 12'h555;
rom[18450] = 12'h555;
rom[18451] = 12'h555;
rom[18452] = 12'h555;
rom[18453] = 12'h555;
rom[18454] = 12'h555;
rom[18455] = 12'h555;
rom[18456] = 12'h555;
rom[18457] = 12'h555;
rom[18458] = 12'h555;
rom[18459] = 12'h555;
rom[18460] = 12'h555;
rom[18461] = 12'h555;
rom[18462] = 12'h555;
rom[18463] = 12'h555;
rom[18464] = 12'h555;
rom[18465] = 12'h555;
rom[18466] = 12'h555;
rom[18467] = 12'h555;
rom[18468] = 12'h555;
rom[18469] = 12'h666;
rom[18470] = 12'h777;
rom[18471] = 12'h777;
rom[18472] = 12'h777;
rom[18473] = 12'h777;
rom[18474] = 12'h777;
rom[18475] = 12'h777;
rom[18476] = 12'h777;
rom[18477] = 12'h777;
rom[18478] = 12'h777;
rom[18479] = 12'h777;
rom[18480] = 12'h777;
rom[18481] = 12'h777;
rom[18482] = 12'h777;
rom[18483] = 12'h666;
rom[18484] = 12'h666;
rom[18485] = 12'h555;
rom[18486] = 12'h444;
rom[18487] = 12'h333;
rom[18488] = 12'h333;
rom[18489] = 12'h222;
rom[18490] = 12'h222;
rom[18491] = 12'h222;
rom[18492] = 12'h111;
rom[18493] = 12'h111;
rom[18494] = 12'h111;
rom[18495] = 12'h111;
rom[18496] = 12'h  0;
rom[18497] = 12'h  0;
rom[18498] = 12'h  0;
rom[18499] = 12'h  0;
rom[18500] = 12'h  0;
rom[18501] = 12'h  0;
rom[18502] = 12'h  0;
rom[18503] = 12'h  0;
rom[18504] = 12'h  0;
rom[18505] = 12'h  0;
rom[18506] = 12'h  0;
rom[18507] = 12'h  0;
rom[18508] = 12'h  0;
rom[18509] = 12'h  0;
rom[18510] = 12'h  0;
rom[18511] = 12'h  0;
rom[18512] = 12'h  0;
rom[18513] = 12'h  0;
rom[18514] = 12'h100;
rom[18515] = 12'h200;
rom[18516] = 12'h300;
rom[18517] = 12'h400;
rom[18518] = 12'h500;
rom[18519] = 12'h710;
rom[18520] = 12'h820;
rom[18521] = 12'h921;
rom[18522] = 12'ha31;
rom[18523] = 12'hb31;
rom[18524] = 12'hb30;
rom[18525] = 12'ha20;
rom[18526] = 12'ha30;
rom[18527] = 12'ha30;
rom[18528] = 12'h931;
rom[18529] = 12'h821;
rom[18530] = 12'h810;
rom[18531] = 12'h710;
rom[18532] = 12'h710;
rom[18533] = 12'h610;
rom[18534] = 12'h610;
rom[18535] = 12'h510;
rom[18536] = 12'h510;
rom[18537] = 12'h410;
rom[18538] = 12'h300;
rom[18539] = 12'h200;
rom[18540] = 12'h200;
rom[18541] = 12'h100;
rom[18542] = 12'h100;
rom[18543] = 12'h100;
rom[18544] = 12'h100;
rom[18545] = 12'h100;
rom[18546] = 12'h100;
rom[18547] = 12'h  0;
rom[18548] = 12'h  0;
rom[18549] = 12'h  0;
rom[18550] = 12'h  0;
rom[18551] = 12'h  0;
rom[18552] = 12'h  0;
rom[18553] = 12'h  0;
rom[18554] = 12'h  0;
rom[18555] = 12'h  0;
rom[18556] = 12'h  0;
rom[18557] = 12'h  0;
rom[18558] = 12'h  0;
rom[18559] = 12'h  0;
rom[18560] = 12'h  0;
rom[18561] = 12'h100;
rom[18562] = 12'h100;
rom[18563] = 12'h100;
rom[18564] = 12'h100;
rom[18565] = 12'h100;
rom[18566] = 12'h100;
rom[18567] = 12'h100;
rom[18568] = 12'h200;
rom[18569] = 12'h200;
rom[18570] = 12'h200;
rom[18571] = 12'h300;
rom[18572] = 12'h300;
rom[18573] = 12'h300;
rom[18574] = 12'h300;
rom[18575] = 12'h300;
rom[18576] = 12'h300;
rom[18577] = 12'h300;
rom[18578] = 12'h300;
rom[18579] = 12'h300;
rom[18580] = 12'h300;
rom[18581] = 12'h300;
rom[18582] = 12'h200;
rom[18583] = 12'h200;
rom[18584] = 12'h200;
rom[18585] = 12'h100;
rom[18586] = 12'h100;
rom[18587] = 12'h100;
rom[18588] = 12'h100;
rom[18589] = 12'h100;
rom[18590] = 12'h100;
rom[18591] = 12'h100;
rom[18592] = 12'h100;
rom[18593] = 12'h100;
rom[18594] = 12'h100;
rom[18595] = 12'h211;
rom[18596] = 12'h322;
rom[18597] = 12'h433;
rom[18598] = 12'h545;
rom[18599] = 12'h766;
rom[18600] = 12'h888;
rom[18601] = 12'ha9a;
rom[18602] = 12'hcbb;
rom[18603] = 12'hccc;
rom[18604] = 12'hcbb;
rom[18605] = 12'hbbb;
rom[18606] = 12'hbbb;
rom[18607] = 12'hbbb;
rom[18608] = 12'habb;
rom[18609] = 12'haaa;
rom[18610] = 12'haaa;
rom[18611] = 12'h9aa;
rom[18612] = 12'h999;
rom[18613] = 12'h999;
rom[18614] = 12'h899;
rom[18615] = 12'h888;
rom[18616] = 12'h899;
rom[18617] = 12'h888;
rom[18618] = 12'h888;
rom[18619] = 12'h888;
rom[18620] = 12'h888;
rom[18621] = 12'h888;
rom[18622] = 12'h888;
rom[18623] = 12'h888;
rom[18624] = 12'h777;
rom[18625] = 12'h888;
rom[18626] = 12'h888;
rom[18627] = 12'h888;
rom[18628] = 12'h888;
rom[18629] = 12'h888;
rom[18630] = 12'h777;
rom[18631] = 12'h777;
rom[18632] = 12'h777;
rom[18633] = 12'h777;
rom[18634] = 12'h666;
rom[18635] = 12'h777;
rom[18636] = 12'h777;
rom[18637] = 12'h777;
rom[18638] = 12'h777;
rom[18639] = 12'h777;
rom[18640] = 12'h777;
rom[18641] = 12'h777;
rom[18642] = 12'h666;
rom[18643] = 12'h555;
rom[18644] = 12'h444;
rom[18645] = 12'h444;
rom[18646] = 12'h444;
rom[18647] = 12'h444;
rom[18648] = 12'h333;
rom[18649] = 12'h333;
rom[18650] = 12'h333;
rom[18651] = 12'h333;
rom[18652] = 12'h333;
rom[18653] = 12'h222;
rom[18654] = 12'h222;
rom[18655] = 12'h222;
rom[18656] = 12'h222;
rom[18657] = 12'h222;
rom[18658] = 12'h111;
rom[18659] = 12'h111;
rom[18660] = 12'h111;
rom[18661] = 12'h111;
rom[18662] = 12'h111;
rom[18663] = 12'h111;
rom[18664] = 12'h  0;
rom[18665] = 12'h  0;
rom[18666] = 12'h  0;
rom[18667] = 12'h  0;
rom[18668] = 12'h  0;
rom[18669] = 12'h  0;
rom[18670] = 12'h  0;
rom[18671] = 12'h  0;
rom[18672] = 12'h  0;
rom[18673] = 12'h  0;
rom[18674] = 12'h  0;
rom[18675] = 12'h  0;
rom[18676] = 12'h  0;
rom[18677] = 12'h  0;
rom[18678] = 12'h  0;
rom[18679] = 12'h  0;
rom[18680] = 12'h  0;
rom[18681] = 12'h  0;
rom[18682] = 12'h  0;
rom[18683] = 12'h  0;
rom[18684] = 12'h  0;
rom[18685] = 12'h  0;
rom[18686] = 12'h  0;
rom[18687] = 12'h  0;
rom[18688] = 12'h  0;
rom[18689] = 12'h  0;
rom[18690] = 12'h  0;
rom[18691] = 12'h  0;
rom[18692] = 12'h  0;
rom[18693] = 12'h  0;
rom[18694] = 12'h  0;
rom[18695] = 12'h111;
rom[18696] = 12'h111;
rom[18697] = 12'h111;
rom[18698] = 12'h111;
rom[18699] = 12'h111;
rom[18700] = 12'h111;
rom[18701] = 12'h111;
rom[18702] = 12'h111;
rom[18703] = 12'h111;
rom[18704] = 12'h111;
rom[18705] = 12'h111;
rom[18706] = 12'h222;
rom[18707] = 12'h222;
rom[18708] = 12'h333;
rom[18709] = 12'h333;
rom[18710] = 12'h333;
rom[18711] = 12'h333;
rom[18712] = 12'h333;
rom[18713] = 12'h333;
rom[18714] = 12'h333;
rom[18715] = 12'h333;
rom[18716] = 12'h333;
rom[18717] = 12'h444;
rom[18718] = 12'h333;
rom[18719] = 12'h222;
rom[18720] = 12'h333;
rom[18721] = 12'h333;
rom[18722] = 12'h333;
rom[18723] = 12'h333;
rom[18724] = 12'h333;
rom[18725] = 12'h333;
rom[18726] = 12'h444;
rom[18727] = 12'h444;
rom[18728] = 12'h333;
rom[18729] = 12'h333;
rom[18730] = 12'h222;
rom[18731] = 12'h222;
rom[18732] = 12'h222;
rom[18733] = 12'h111;
rom[18734] = 12'h111;
rom[18735] = 12'h111;
rom[18736] = 12'h111;
rom[18737] = 12'h111;
rom[18738] = 12'h222;
rom[18739] = 12'h222;
rom[18740] = 12'h333;
rom[18741] = 12'h333;
rom[18742] = 12'h333;
rom[18743] = 12'h333;
rom[18744] = 12'h333;
rom[18745] = 12'h444;
rom[18746] = 12'h444;
rom[18747] = 12'h555;
rom[18748] = 12'h555;
rom[18749] = 12'h555;
rom[18750] = 12'h666;
rom[18751] = 12'h666;
rom[18752] = 12'h555;
rom[18753] = 12'h555;
rom[18754] = 12'h555;
rom[18755] = 12'h555;
rom[18756] = 12'h555;
rom[18757] = 12'h555;
rom[18758] = 12'h555;
rom[18759] = 12'h555;
rom[18760] = 12'h555;
rom[18761] = 12'h555;
rom[18762] = 12'h444;
rom[18763] = 12'h444;
rom[18764] = 12'h444;
rom[18765] = 12'h444;
rom[18766] = 12'h444;
rom[18767] = 12'h444;
rom[18768] = 12'h444;
rom[18769] = 12'h444;
rom[18770] = 12'h555;
rom[18771] = 12'h555;
rom[18772] = 12'h555;
rom[18773] = 12'h555;
rom[18774] = 12'h555;
rom[18775] = 12'h555;
rom[18776] = 12'h555;
rom[18777] = 12'h555;
rom[18778] = 12'h555;
rom[18779] = 12'h555;
rom[18780] = 12'h666;
rom[18781] = 12'h666;
rom[18782] = 12'h666;
rom[18783] = 12'h666;
rom[18784] = 12'h666;
rom[18785] = 12'h777;
rom[18786] = 12'h888;
rom[18787] = 12'h888;
rom[18788] = 12'h888;
rom[18789] = 12'h888;
rom[18790] = 12'h888;
rom[18791] = 12'h888;
rom[18792] = 12'h888;
rom[18793] = 12'h888;
rom[18794] = 12'h999;
rom[18795] = 12'h999;
rom[18796] = 12'haaa;
rom[18797] = 12'haaa;
rom[18798] = 12'haaa;
rom[18799] = 12'haaa;
rom[18800] = 12'h333;
rom[18801] = 12'h333;
rom[18802] = 12'h333;
rom[18803] = 12'h333;
rom[18804] = 12'h333;
rom[18805] = 12'h333;
rom[18806] = 12'h333;
rom[18807] = 12'h333;
rom[18808] = 12'h333;
rom[18809] = 12'h333;
rom[18810] = 12'h333;
rom[18811] = 12'h333;
rom[18812] = 12'h333;
rom[18813] = 12'h333;
rom[18814] = 12'h333;
rom[18815] = 12'h444;
rom[18816] = 12'h444;
rom[18817] = 12'h444;
rom[18818] = 12'h444;
rom[18819] = 12'h555;
rom[18820] = 12'h555;
rom[18821] = 12'h555;
rom[18822] = 12'h555;
rom[18823] = 12'h555;
rom[18824] = 12'h666;
rom[18825] = 12'h666;
rom[18826] = 12'h666;
rom[18827] = 12'h666;
rom[18828] = 12'h666;
rom[18829] = 12'h666;
rom[18830] = 12'h666;
rom[18831] = 12'h666;
rom[18832] = 12'h666;
rom[18833] = 12'h777;
rom[18834] = 12'h777;
rom[18835] = 12'h777;
rom[18836] = 12'h777;
rom[18837] = 12'h777;
rom[18838] = 12'h777;
rom[18839] = 12'h777;
rom[18840] = 12'h777;
rom[18841] = 12'h777;
rom[18842] = 12'h777;
rom[18843] = 12'h666;
rom[18844] = 12'h666;
rom[18845] = 12'h666;
rom[18846] = 12'h666;
rom[18847] = 12'h666;
rom[18848] = 12'h666;
rom[18849] = 12'h666;
rom[18850] = 12'h555;
rom[18851] = 12'h555;
rom[18852] = 12'h555;
rom[18853] = 12'h555;
rom[18854] = 12'h555;
rom[18855] = 12'h555;
rom[18856] = 12'h555;
rom[18857] = 12'h555;
rom[18858] = 12'h555;
rom[18859] = 12'h555;
rom[18860] = 12'h555;
rom[18861] = 12'h555;
rom[18862] = 12'h555;
rom[18863] = 12'h555;
rom[18864] = 12'h555;
rom[18865] = 12'h555;
rom[18866] = 12'h555;
rom[18867] = 12'h555;
rom[18868] = 12'h555;
rom[18869] = 12'h555;
rom[18870] = 12'h666;
rom[18871] = 12'h666;
rom[18872] = 12'h777;
rom[18873] = 12'h777;
rom[18874] = 12'h777;
rom[18875] = 12'h777;
rom[18876] = 12'h777;
rom[18877] = 12'h777;
rom[18878] = 12'h777;
rom[18879] = 12'h777;
rom[18880] = 12'h777;
rom[18881] = 12'h777;
rom[18882] = 12'h777;
rom[18883] = 12'h666;
rom[18884] = 12'h666;
rom[18885] = 12'h555;
rom[18886] = 12'h444;
rom[18887] = 12'h444;
rom[18888] = 12'h333;
rom[18889] = 12'h222;
rom[18890] = 12'h222;
rom[18891] = 12'h222;
rom[18892] = 12'h111;
rom[18893] = 12'h111;
rom[18894] = 12'h111;
rom[18895] = 12'h111;
rom[18896] = 12'h  0;
rom[18897] = 12'h  0;
rom[18898] = 12'h  0;
rom[18899] = 12'h  0;
rom[18900] = 12'h  0;
rom[18901] = 12'h  0;
rom[18902] = 12'h  0;
rom[18903] = 12'h  0;
rom[18904] = 12'h  0;
rom[18905] = 12'h  0;
rom[18906] = 12'h  0;
rom[18907] = 12'h  0;
rom[18908] = 12'h  0;
rom[18909] = 12'h  0;
rom[18910] = 12'h  0;
rom[18911] = 12'h  0;
rom[18912] = 12'h  0;
rom[18913] = 12'h  0;
rom[18914] = 12'h100;
rom[18915] = 12'h200;
rom[18916] = 12'h300;
rom[18917] = 12'h400;
rom[18918] = 12'h500;
rom[18919] = 12'h610;
rom[18920] = 12'h810;
rom[18921] = 12'h921;
rom[18922] = 12'hb31;
rom[18923] = 12'hb41;
rom[18924] = 12'hb30;
rom[18925] = 12'ha30;
rom[18926] = 12'hb30;
rom[18927] = 12'ha30;
rom[18928] = 12'ha30;
rom[18929] = 12'h920;
rom[18930] = 12'h820;
rom[18931] = 12'h710;
rom[18932] = 12'h710;
rom[18933] = 12'h610;
rom[18934] = 12'h610;
rom[18935] = 12'h510;
rom[18936] = 12'h510;
rom[18937] = 12'h410;
rom[18938] = 12'h300;
rom[18939] = 12'h200;
rom[18940] = 12'h200;
rom[18941] = 12'h100;
rom[18942] = 12'h100;
rom[18943] = 12'h100;
rom[18944] = 12'h100;
rom[18945] = 12'h100;
rom[18946] = 12'h100;
rom[18947] = 12'h  0;
rom[18948] = 12'h  0;
rom[18949] = 12'h  0;
rom[18950] = 12'h  0;
rom[18951] = 12'h  0;
rom[18952] = 12'h  0;
rom[18953] = 12'h  0;
rom[18954] = 12'h  0;
rom[18955] = 12'h  0;
rom[18956] = 12'h  0;
rom[18957] = 12'h  0;
rom[18958] = 12'h  0;
rom[18959] = 12'h  0;
rom[18960] = 12'h  0;
rom[18961] = 12'h100;
rom[18962] = 12'h100;
rom[18963] = 12'h100;
rom[18964] = 12'h100;
rom[18965] = 12'h100;
rom[18966] = 12'h100;
rom[18967] = 12'h200;
rom[18968] = 12'h200;
rom[18969] = 12'h200;
rom[18970] = 12'h300;
rom[18971] = 12'h300;
rom[18972] = 12'h300;
rom[18973] = 12'h300;
rom[18974] = 12'h400;
rom[18975] = 12'h400;
rom[18976] = 12'h300;
rom[18977] = 12'h300;
rom[18978] = 12'h300;
rom[18979] = 12'h300;
rom[18980] = 12'h300;
rom[18981] = 12'h200;
rom[18982] = 12'h200;
rom[18983] = 12'h200;
rom[18984] = 12'h100;
rom[18985] = 12'h100;
rom[18986] = 12'h100;
rom[18987] = 12'h100;
rom[18988] = 12'h100;
rom[18989] = 12'h100;
rom[18990] = 12'h100;
rom[18991] = 12'h100;
rom[18992] = 12'h100;
rom[18993] = 12'h  0;
rom[18994] = 12'h100;
rom[18995] = 12'h211;
rom[18996] = 12'h322;
rom[18997] = 12'h333;
rom[18998] = 12'h544;
rom[18999] = 12'h655;
rom[19000] = 12'h877;
rom[19001] = 12'ha99;
rom[19002] = 12'hcbb;
rom[19003] = 12'hccc;
rom[19004] = 12'hcbb;
rom[19005] = 12'hbbb;
rom[19006] = 12'hbbb;
rom[19007] = 12'hbbb;
rom[19008] = 12'hbbb;
rom[19009] = 12'haaa;
rom[19010] = 12'haaa;
rom[19011] = 12'haaa;
rom[19012] = 12'h9aa;
rom[19013] = 12'h999;
rom[19014] = 12'h999;
rom[19015] = 12'h888;
rom[19016] = 12'h899;
rom[19017] = 12'h888;
rom[19018] = 12'h888;
rom[19019] = 12'h888;
rom[19020] = 12'h888;
rom[19021] = 12'h888;
rom[19022] = 12'h888;
rom[19023] = 12'h888;
rom[19024] = 12'h888;
rom[19025] = 12'h888;
rom[19026] = 12'h888;
rom[19027] = 12'h888;
rom[19028] = 12'h888;
rom[19029] = 12'h888;
rom[19030] = 12'h777;
rom[19031] = 12'h777;
rom[19032] = 12'h777;
rom[19033] = 12'h777;
rom[19034] = 12'h777;
rom[19035] = 12'h777;
rom[19036] = 12'h777;
rom[19037] = 12'h888;
rom[19038] = 12'h888;
rom[19039] = 12'h888;
rom[19040] = 12'h777;
rom[19041] = 12'h666;
rom[19042] = 12'h555;
rom[19043] = 12'h444;
rom[19044] = 12'h444;
rom[19045] = 12'h444;
rom[19046] = 12'h444;
rom[19047] = 12'h444;
rom[19048] = 12'h333;
rom[19049] = 12'h333;
rom[19050] = 12'h333;
rom[19051] = 12'h333;
rom[19052] = 12'h333;
rom[19053] = 12'h222;
rom[19054] = 12'h222;
rom[19055] = 12'h222;
rom[19056] = 12'h222;
rom[19057] = 12'h111;
rom[19058] = 12'h111;
rom[19059] = 12'h111;
rom[19060] = 12'h111;
rom[19061] = 12'h111;
rom[19062] = 12'h111;
rom[19063] = 12'h111;
rom[19064] = 12'h  0;
rom[19065] = 12'h  0;
rom[19066] = 12'h  0;
rom[19067] = 12'h  0;
rom[19068] = 12'h  0;
rom[19069] = 12'h  0;
rom[19070] = 12'h  0;
rom[19071] = 12'h  0;
rom[19072] = 12'h  0;
rom[19073] = 12'h  0;
rom[19074] = 12'h  0;
rom[19075] = 12'h  0;
rom[19076] = 12'h  0;
rom[19077] = 12'h  0;
rom[19078] = 12'h  0;
rom[19079] = 12'h  0;
rom[19080] = 12'h  0;
rom[19081] = 12'h  0;
rom[19082] = 12'h  0;
rom[19083] = 12'h  0;
rom[19084] = 12'h  0;
rom[19085] = 12'h  0;
rom[19086] = 12'h  0;
rom[19087] = 12'h  0;
rom[19088] = 12'h  0;
rom[19089] = 12'h  0;
rom[19090] = 12'h  0;
rom[19091] = 12'h  0;
rom[19092] = 12'h  0;
rom[19093] = 12'h  0;
rom[19094] = 12'h111;
rom[19095] = 12'h111;
rom[19096] = 12'h111;
rom[19097] = 12'h111;
rom[19098] = 12'h111;
rom[19099] = 12'h111;
rom[19100] = 12'h111;
rom[19101] = 12'h111;
rom[19102] = 12'h111;
rom[19103] = 12'h111;
rom[19104] = 12'h111;
rom[19105] = 12'h111;
rom[19106] = 12'h222;
rom[19107] = 12'h222;
rom[19108] = 12'h333;
rom[19109] = 12'h333;
rom[19110] = 12'h333;
rom[19111] = 12'h333;
rom[19112] = 12'h222;
rom[19113] = 12'h333;
rom[19114] = 12'h333;
rom[19115] = 12'h333;
rom[19116] = 12'h333;
rom[19117] = 12'h333;
rom[19118] = 12'h333;
rom[19119] = 12'h222;
rom[19120] = 12'h333;
rom[19121] = 12'h333;
rom[19122] = 12'h333;
rom[19123] = 12'h333;
rom[19124] = 12'h333;
rom[19125] = 12'h333;
rom[19126] = 12'h444;
rom[19127] = 12'h444;
rom[19128] = 12'h444;
rom[19129] = 12'h333;
rom[19130] = 12'h222;
rom[19131] = 12'h222;
rom[19132] = 12'h222;
rom[19133] = 12'h222;
rom[19134] = 12'h222;
rom[19135] = 12'h222;
rom[19136] = 12'h222;
rom[19137] = 12'h222;
rom[19138] = 12'h333;
rom[19139] = 12'h333;
rom[19140] = 12'h444;
rom[19141] = 12'h444;
rom[19142] = 12'h333;
rom[19143] = 12'h333;
rom[19144] = 12'h333;
rom[19145] = 12'h333;
rom[19146] = 12'h444;
rom[19147] = 12'h444;
rom[19148] = 12'h555;
rom[19149] = 12'h555;
rom[19150] = 12'h666;
rom[19151] = 12'h666;
rom[19152] = 12'h555;
rom[19153] = 12'h555;
rom[19154] = 12'h555;
rom[19155] = 12'h555;
rom[19156] = 12'h555;
rom[19157] = 12'h555;
rom[19158] = 12'h555;
rom[19159] = 12'h555;
rom[19160] = 12'h444;
rom[19161] = 12'h444;
rom[19162] = 12'h444;
rom[19163] = 12'h444;
rom[19164] = 12'h444;
rom[19165] = 12'h444;
rom[19166] = 12'h444;
rom[19167] = 12'h444;
rom[19168] = 12'h444;
rom[19169] = 12'h444;
rom[19170] = 12'h555;
rom[19171] = 12'h555;
rom[19172] = 12'h555;
rom[19173] = 12'h555;
rom[19174] = 12'h555;
rom[19175] = 12'h555;
rom[19176] = 12'h555;
rom[19177] = 12'h666;
rom[19178] = 12'h666;
rom[19179] = 12'h666;
rom[19180] = 12'h666;
rom[19181] = 12'h666;
rom[19182] = 12'h666;
rom[19183] = 12'h666;
rom[19184] = 12'h666;
rom[19185] = 12'h666;
rom[19186] = 12'h777;
rom[19187] = 12'h888;
rom[19188] = 12'h888;
rom[19189] = 12'h888;
rom[19190] = 12'h888;
rom[19191] = 12'h888;
rom[19192] = 12'h888;
rom[19193] = 12'h888;
rom[19194] = 12'h999;
rom[19195] = 12'h999;
rom[19196] = 12'haaa;
rom[19197] = 12'haaa;
rom[19198] = 12'haaa;
rom[19199] = 12'haaa;
rom[19200] = 12'h333;
rom[19201] = 12'h333;
rom[19202] = 12'h333;
rom[19203] = 12'h333;
rom[19204] = 12'h333;
rom[19205] = 12'h333;
rom[19206] = 12'h333;
rom[19207] = 12'h333;
rom[19208] = 12'h333;
rom[19209] = 12'h333;
rom[19210] = 12'h333;
rom[19211] = 12'h444;
rom[19212] = 12'h444;
rom[19213] = 12'h444;
rom[19214] = 12'h444;
rom[19215] = 12'h444;
rom[19216] = 12'h555;
rom[19217] = 12'h555;
rom[19218] = 12'h555;
rom[19219] = 12'h555;
rom[19220] = 12'h555;
rom[19221] = 12'h555;
rom[19222] = 12'h666;
rom[19223] = 12'h666;
rom[19224] = 12'h666;
rom[19225] = 12'h666;
rom[19226] = 12'h777;
rom[19227] = 12'h777;
rom[19228] = 12'h777;
rom[19229] = 12'h777;
rom[19230] = 12'h777;
rom[19231] = 12'h777;
rom[19232] = 12'h777;
rom[19233] = 12'h777;
rom[19234] = 12'h777;
rom[19235] = 12'h777;
rom[19236] = 12'h777;
rom[19237] = 12'h777;
rom[19238] = 12'h777;
rom[19239] = 12'h777;
rom[19240] = 12'h777;
rom[19241] = 12'h777;
rom[19242] = 12'h777;
rom[19243] = 12'h777;
rom[19244] = 12'h777;
rom[19245] = 12'h777;
rom[19246] = 12'h777;
rom[19247] = 12'h777;
rom[19248] = 12'h666;
rom[19249] = 12'h666;
rom[19250] = 12'h555;
rom[19251] = 12'h555;
rom[19252] = 12'h555;
rom[19253] = 12'h555;
rom[19254] = 12'h555;
rom[19255] = 12'h555;
rom[19256] = 12'h555;
rom[19257] = 12'h555;
rom[19258] = 12'h555;
rom[19259] = 12'h555;
rom[19260] = 12'h555;
rom[19261] = 12'h555;
rom[19262] = 12'h555;
rom[19263] = 12'h555;
rom[19264] = 12'h555;
rom[19265] = 12'h555;
rom[19266] = 12'h555;
rom[19267] = 12'h555;
rom[19268] = 12'h666;
rom[19269] = 12'h666;
rom[19270] = 12'h666;
rom[19271] = 12'h666;
rom[19272] = 12'h666;
rom[19273] = 12'h666;
rom[19274] = 12'h666;
rom[19275] = 12'h777;
rom[19276] = 12'h777;
rom[19277] = 12'h888;
rom[19278] = 12'h777;
rom[19279] = 12'h777;
rom[19280] = 12'h777;
rom[19281] = 12'h777;
rom[19282] = 12'h777;
rom[19283] = 12'h777;
rom[19284] = 12'h666;
rom[19285] = 12'h666;
rom[19286] = 12'h555;
rom[19287] = 12'h444;
rom[19288] = 12'h333;
rom[19289] = 12'h222;
rom[19290] = 12'h222;
rom[19291] = 12'h222;
rom[19292] = 12'h111;
rom[19293] = 12'h111;
rom[19294] = 12'h111;
rom[19295] = 12'h  0;
rom[19296] = 12'h  0;
rom[19297] = 12'h  0;
rom[19298] = 12'h  0;
rom[19299] = 12'h  0;
rom[19300] = 12'h  0;
rom[19301] = 12'h  0;
rom[19302] = 12'h  0;
rom[19303] = 12'h  0;
rom[19304] = 12'h  0;
rom[19305] = 12'h  0;
rom[19306] = 12'h  0;
rom[19307] = 12'h  0;
rom[19308] = 12'h  0;
rom[19309] = 12'h  0;
rom[19310] = 12'h  0;
rom[19311] = 12'h  0;
rom[19312] = 12'h  0;
rom[19313] = 12'h  0;
rom[19314] = 12'h100;
rom[19315] = 12'h200;
rom[19316] = 12'h200;
rom[19317] = 12'h400;
rom[19318] = 12'h510;
rom[19319] = 12'h610;
rom[19320] = 12'h820;
rom[19321] = 12'h920;
rom[19322] = 12'hb31;
rom[19323] = 12'hb41;
rom[19324] = 12'hb30;
rom[19325] = 12'hb30;
rom[19326] = 12'hb30;
rom[19327] = 12'hb30;
rom[19328] = 12'h930;
rom[19329] = 12'h930;
rom[19330] = 12'h830;
rom[19331] = 12'h820;
rom[19332] = 12'h720;
rom[19333] = 12'h710;
rom[19334] = 12'h610;
rom[19335] = 12'h510;
rom[19336] = 12'h510;
rom[19337] = 12'h400;
rom[19338] = 12'h300;
rom[19339] = 12'h200;
rom[19340] = 12'h200;
rom[19341] = 12'h100;
rom[19342] = 12'h100;
rom[19343] = 12'h100;
rom[19344] = 12'h100;
rom[19345] = 12'h  0;
rom[19346] = 12'h  0;
rom[19347] = 12'h  0;
rom[19348] = 12'h  0;
rom[19349] = 12'h  0;
rom[19350] = 12'h  0;
rom[19351] = 12'h  0;
rom[19352] = 12'h  0;
rom[19353] = 12'h  0;
rom[19354] = 12'h  0;
rom[19355] = 12'h  0;
rom[19356] = 12'h  0;
rom[19357] = 12'h  0;
rom[19358] = 12'h  0;
rom[19359] = 12'h  0;
rom[19360] = 12'h  0;
rom[19361] = 12'h  0;
rom[19362] = 12'h  0;
rom[19363] = 12'h100;
rom[19364] = 12'h100;
rom[19365] = 12'h200;
rom[19366] = 12'h200;
rom[19367] = 12'h300;
rom[19368] = 12'h300;
rom[19369] = 12'h300;
rom[19370] = 12'h300;
rom[19371] = 12'h400;
rom[19372] = 12'h400;
rom[19373] = 12'h400;
rom[19374] = 12'h400;
rom[19375] = 12'h400;
rom[19376] = 12'h300;
rom[19377] = 12'h300;
rom[19378] = 12'h300;
rom[19379] = 12'h300;
rom[19380] = 12'h300;
rom[19381] = 12'h200;
rom[19382] = 12'h200;
rom[19383] = 12'h200;
rom[19384] = 12'h100;
rom[19385] = 12'h100;
rom[19386] = 12'h100;
rom[19387] = 12'h100;
rom[19388] = 12'h100;
rom[19389] = 12'h100;
rom[19390] = 12'h100;
rom[19391] = 12'h100;
rom[19392] = 12'h100;
rom[19393] = 12'h100;
rom[19394] = 12'h100;
rom[19395] = 12'h212;
rom[19396] = 12'h322;
rom[19397] = 12'h333;
rom[19398] = 12'h444;
rom[19399] = 12'h655;
rom[19400] = 12'h766;
rom[19401] = 12'h988;
rom[19402] = 12'hbab;
rom[19403] = 12'hcbb;
rom[19404] = 12'hbbb;
rom[19405] = 12'hbbb;
rom[19406] = 12'hbbb;
rom[19407] = 12'hbbb;
rom[19408] = 12'haaa;
rom[19409] = 12'haaa;
rom[19410] = 12'haaa;
rom[19411] = 12'haaa;
rom[19412] = 12'h9aa;
rom[19413] = 12'h999;
rom[19414] = 12'h999;
rom[19415] = 12'h999;
rom[19416] = 12'h888;
rom[19417] = 12'h888;
rom[19418] = 12'h888;
rom[19419] = 12'h888;
rom[19420] = 12'h888;
rom[19421] = 12'h888;
rom[19422] = 12'h888;
rom[19423] = 12'h888;
rom[19424] = 12'h888;
rom[19425] = 12'h888;
rom[19426] = 12'h888;
rom[19427] = 12'h888;
rom[19428] = 12'h888;
rom[19429] = 12'h888;
rom[19430] = 12'h888;
rom[19431] = 12'h777;
rom[19432] = 12'h888;
rom[19433] = 12'h888;
rom[19434] = 12'h888;
rom[19435] = 12'h888;
rom[19436] = 12'h888;
rom[19437] = 12'h888;
rom[19438] = 12'h777;
rom[19439] = 12'h666;
rom[19440] = 12'h555;
rom[19441] = 12'h555;
rom[19442] = 12'h555;
rom[19443] = 12'h555;
rom[19444] = 12'h555;
rom[19445] = 12'h444;
rom[19446] = 12'h444;
rom[19447] = 12'h444;
rom[19448] = 12'h444;
rom[19449] = 12'h333;
rom[19450] = 12'h333;
rom[19451] = 12'h222;
rom[19452] = 12'h222;
rom[19453] = 12'h222;
rom[19454] = 12'h222;
rom[19455] = 12'h222;
rom[19456] = 12'h111;
rom[19457] = 12'h111;
rom[19458] = 12'h111;
rom[19459] = 12'h111;
rom[19460] = 12'h111;
rom[19461] = 12'h111;
rom[19462] = 12'h  0;
rom[19463] = 12'h  0;
rom[19464] = 12'h  0;
rom[19465] = 12'h  0;
rom[19466] = 12'h  0;
rom[19467] = 12'h  0;
rom[19468] = 12'h  0;
rom[19469] = 12'h  0;
rom[19470] = 12'h  0;
rom[19471] = 12'h  0;
rom[19472] = 12'h  0;
rom[19473] = 12'h  0;
rom[19474] = 12'h  0;
rom[19475] = 12'h  0;
rom[19476] = 12'h  0;
rom[19477] = 12'h  0;
rom[19478] = 12'h  0;
rom[19479] = 12'h  0;
rom[19480] = 12'h  0;
rom[19481] = 12'h  0;
rom[19482] = 12'h  0;
rom[19483] = 12'h  0;
rom[19484] = 12'h  0;
rom[19485] = 12'h  0;
rom[19486] = 12'h  0;
rom[19487] = 12'h  0;
rom[19488] = 12'h  0;
rom[19489] = 12'h  0;
rom[19490] = 12'h  0;
rom[19491] = 12'h  0;
rom[19492] = 12'h  0;
rom[19493] = 12'h  0;
rom[19494] = 12'h111;
rom[19495] = 12'h111;
rom[19496] = 12'h111;
rom[19497] = 12'h111;
rom[19498] = 12'h111;
rom[19499] = 12'h111;
rom[19500] = 12'h111;
rom[19501] = 12'h111;
rom[19502] = 12'h111;
rom[19503] = 12'h111;
rom[19504] = 12'h111;
rom[19505] = 12'h222;
rom[19506] = 12'h222;
rom[19507] = 12'h333;
rom[19508] = 12'h333;
rom[19509] = 12'h333;
rom[19510] = 12'h333;
rom[19511] = 12'h333;
rom[19512] = 12'h333;
rom[19513] = 12'h333;
rom[19514] = 12'h333;
rom[19515] = 12'h333;
rom[19516] = 12'h333;
rom[19517] = 12'h333;
rom[19518] = 12'h333;
rom[19519] = 12'h222;
rom[19520] = 12'h333;
rom[19521] = 12'h333;
rom[19522] = 12'h333;
rom[19523] = 12'h333;
rom[19524] = 12'h333;
rom[19525] = 12'h444;
rom[19526] = 12'h444;
rom[19527] = 12'h444;
rom[19528] = 12'h333;
rom[19529] = 12'h333;
rom[19530] = 12'h333;
rom[19531] = 12'h222;
rom[19532] = 12'h222;
rom[19533] = 12'h222;
rom[19534] = 12'h222;
rom[19535] = 12'h222;
rom[19536] = 12'h222;
rom[19537] = 12'h333;
rom[19538] = 12'h333;
rom[19539] = 12'h333;
rom[19540] = 12'h333;
rom[19541] = 12'h333;
rom[19542] = 12'h333;
rom[19543] = 12'h333;
rom[19544] = 12'h333;
rom[19545] = 12'h444;
rom[19546] = 12'h555;
rom[19547] = 12'h555;
rom[19548] = 12'h655;
rom[19549] = 12'h555;
rom[19550] = 12'h555;
rom[19551] = 12'h555;
rom[19552] = 12'h555;
rom[19553] = 12'h555;
rom[19554] = 12'h555;
rom[19555] = 12'h555;
rom[19556] = 12'h555;
rom[19557] = 12'h455;
rom[19558] = 12'h455;
rom[19559] = 12'h455;
rom[19560] = 12'h555;
rom[19561] = 12'h455;
rom[19562] = 12'h455;
rom[19563] = 12'h455;
rom[19564] = 12'h455;
rom[19565] = 12'h555;
rom[19566] = 12'h555;
rom[19567] = 12'h555;
rom[19568] = 12'h555;
rom[19569] = 12'h555;
rom[19570] = 12'h555;
rom[19571] = 12'h555;
rom[19572] = 12'h555;
rom[19573] = 12'h555;
rom[19574] = 12'h555;
rom[19575] = 12'h555;
rom[19576] = 12'h555;
rom[19577] = 12'h555;
rom[19578] = 12'h666;
rom[19579] = 12'h666;
rom[19580] = 12'h666;
rom[19581] = 12'h666;
rom[19582] = 12'h666;
rom[19583] = 12'h666;
rom[19584] = 12'h666;
rom[19585] = 12'h666;
rom[19586] = 12'h666;
rom[19587] = 12'h777;
rom[19588] = 12'h777;
rom[19589] = 12'h888;
rom[19590] = 12'h888;
rom[19591] = 12'h888;
rom[19592] = 12'h888;
rom[19593] = 12'h888;
rom[19594] = 12'h999;
rom[19595] = 12'h999;
rom[19596] = 12'haaa;
rom[19597] = 12'haaa;
rom[19598] = 12'haaa;
rom[19599] = 12'haaa;
rom[19600] = 12'h333;
rom[19601] = 12'h333;
rom[19602] = 12'h333;
rom[19603] = 12'h333;
rom[19604] = 12'h444;
rom[19605] = 12'h444;
rom[19606] = 12'h444;
rom[19607] = 12'h444;
rom[19608] = 12'h444;
rom[19609] = 12'h444;
rom[19610] = 12'h444;
rom[19611] = 12'h444;
rom[19612] = 12'h555;
rom[19613] = 12'h555;
rom[19614] = 12'h555;
rom[19615] = 12'h555;
rom[19616] = 12'h555;
rom[19617] = 12'h555;
rom[19618] = 12'h666;
rom[19619] = 12'h666;
rom[19620] = 12'h666;
rom[19621] = 12'h666;
rom[19622] = 12'h666;
rom[19623] = 12'h666;
rom[19624] = 12'h777;
rom[19625] = 12'h777;
rom[19626] = 12'h777;
rom[19627] = 12'h777;
rom[19628] = 12'h777;
rom[19629] = 12'h777;
rom[19630] = 12'h777;
rom[19631] = 12'h777;
rom[19632] = 12'h777;
rom[19633] = 12'h777;
rom[19634] = 12'h777;
rom[19635] = 12'h777;
rom[19636] = 12'h777;
rom[19637] = 12'h777;
rom[19638] = 12'h777;
rom[19639] = 12'h777;
rom[19640] = 12'h777;
rom[19641] = 12'h777;
rom[19642] = 12'h777;
rom[19643] = 12'h777;
rom[19644] = 12'h777;
rom[19645] = 12'h777;
rom[19646] = 12'h777;
rom[19647] = 12'h777;
rom[19648] = 12'h666;
rom[19649] = 12'h666;
rom[19650] = 12'h666;
rom[19651] = 12'h666;
rom[19652] = 12'h666;
rom[19653] = 12'h666;
rom[19654] = 12'h555;
rom[19655] = 12'h555;
rom[19656] = 12'h555;
rom[19657] = 12'h555;
rom[19658] = 12'h555;
rom[19659] = 12'h555;
rom[19660] = 12'h555;
rom[19661] = 12'h555;
rom[19662] = 12'h666;
rom[19663] = 12'h666;
rom[19664] = 12'h555;
rom[19665] = 12'h555;
rom[19666] = 12'h555;
rom[19667] = 12'h555;
rom[19668] = 12'h555;
rom[19669] = 12'h666;
rom[19670] = 12'h666;
rom[19671] = 12'h666;
rom[19672] = 12'h666;
rom[19673] = 12'h666;
rom[19674] = 12'h666;
rom[19675] = 12'h777;
rom[19676] = 12'h777;
rom[19677] = 12'h888;
rom[19678] = 12'h888;
rom[19679] = 12'h777;
rom[19680] = 12'h777;
rom[19681] = 12'h777;
rom[19682] = 12'h777;
rom[19683] = 12'h777;
rom[19684] = 12'h666;
rom[19685] = 12'h666;
rom[19686] = 12'h555;
rom[19687] = 12'h444;
rom[19688] = 12'h333;
rom[19689] = 12'h333;
rom[19690] = 12'h222;
rom[19691] = 12'h222;
rom[19692] = 12'h111;
rom[19693] = 12'h111;
rom[19694] = 12'h111;
rom[19695] = 12'h  0;
rom[19696] = 12'h  0;
rom[19697] = 12'h  0;
rom[19698] = 12'h  0;
rom[19699] = 12'h  0;
rom[19700] = 12'h  0;
rom[19701] = 12'h  0;
rom[19702] = 12'h  0;
rom[19703] = 12'h  0;
rom[19704] = 12'h  0;
rom[19705] = 12'h  0;
rom[19706] = 12'h  0;
rom[19707] = 12'h  0;
rom[19708] = 12'h  0;
rom[19709] = 12'h  0;
rom[19710] = 12'h  0;
rom[19711] = 12'h  0;
rom[19712] = 12'h  0;
rom[19713] = 12'h  0;
rom[19714] = 12'h100;
rom[19715] = 12'h200;
rom[19716] = 12'h200;
rom[19717] = 12'h300;
rom[19718] = 12'h510;
rom[19719] = 12'h610;
rom[19720] = 12'h720;
rom[19721] = 12'h930;
rom[19722] = 12'hb41;
rom[19723] = 12'hb41;
rom[19724] = 12'hb40;
rom[19725] = 12'hb30;
rom[19726] = 12'hb30;
rom[19727] = 12'hb30;
rom[19728] = 12'ha40;
rom[19729] = 12'h930;
rom[19730] = 12'h930;
rom[19731] = 12'h830;
rom[19732] = 12'h820;
rom[19733] = 12'h720;
rom[19734] = 12'h610;
rom[19735] = 12'h610;
rom[19736] = 12'h510;
rom[19737] = 12'h410;
rom[19738] = 12'h400;
rom[19739] = 12'h300;
rom[19740] = 12'h200;
rom[19741] = 12'h200;
rom[19742] = 12'h100;
rom[19743] = 12'h100;
rom[19744] = 12'h  0;
rom[19745] = 12'h  0;
rom[19746] = 12'h  0;
rom[19747] = 12'h  0;
rom[19748] = 12'h  0;
rom[19749] = 12'h  0;
rom[19750] = 12'h  0;
rom[19751] = 12'h  0;
rom[19752] = 12'h  0;
rom[19753] = 12'h  0;
rom[19754] = 12'h  0;
rom[19755] = 12'h  0;
rom[19756] = 12'h  0;
rom[19757] = 12'h  0;
rom[19758] = 12'h  0;
rom[19759] = 12'h  0;
rom[19760] = 12'h  0;
rom[19761] = 12'h  0;
rom[19762] = 12'h  0;
rom[19763] = 12'h100;
rom[19764] = 12'h100;
rom[19765] = 12'h200;
rom[19766] = 12'h200;
rom[19767] = 12'h300;
rom[19768] = 12'h300;
rom[19769] = 12'h300;
rom[19770] = 12'h400;
rom[19771] = 12'h400;
rom[19772] = 12'h400;
rom[19773] = 12'h400;
rom[19774] = 12'h400;
rom[19775] = 12'h400;
rom[19776] = 12'h300;
rom[19777] = 12'h300;
rom[19778] = 12'h300;
rom[19779] = 12'h300;
rom[19780] = 12'h300;
rom[19781] = 12'h200;
rom[19782] = 12'h200;
rom[19783] = 12'h100;
rom[19784] = 12'h100;
rom[19785] = 12'h100;
rom[19786] = 12'h100;
rom[19787] = 12'h100;
rom[19788] = 12'h100;
rom[19789] = 12'h100;
rom[19790] = 12'h100;
rom[19791] = 12'h100;
rom[19792] = 12'h100;
rom[19793] = 12'h100;
rom[19794] = 12'h101;
rom[19795] = 12'h222;
rom[19796] = 12'h323;
rom[19797] = 12'h333;
rom[19798] = 12'h444;
rom[19799] = 12'h555;
rom[19800] = 12'h666;
rom[19801] = 12'h888;
rom[19802] = 12'haaa;
rom[19803] = 12'hbbb;
rom[19804] = 12'hbbb;
rom[19805] = 12'hbbb;
rom[19806] = 12'hbbb;
rom[19807] = 12'hbbb;
rom[19808] = 12'haaa;
rom[19809] = 12'haaa;
rom[19810] = 12'haaa;
rom[19811] = 12'haaa;
rom[19812] = 12'haaa;
rom[19813] = 12'h999;
rom[19814] = 12'h999;
rom[19815] = 12'h999;
rom[19816] = 12'h888;
rom[19817] = 12'h888;
rom[19818] = 12'h888;
rom[19819] = 12'h888;
rom[19820] = 12'h888;
rom[19821] = 12'h888;
rom[19822] = 12'h888;
rom[19823] = 12'h888;
rom[19824] = 12'h888;
rom[19825] = 12'h888;
rom[19826] = 12'h888;
rom[19827] = 12'h888;
rom[19828] = 12'h888;
rom[19829] = 12'h888;
rom[19830] = 12'h888;
rom[19831] = 12'h888;
rom[19832] = 12'h888;
rom[19833] = 12'h888;
rom[19834] = 12'h888;
rom[19835] = 12'h888;
rom[19836] = 12'h888;
rom[19837] = 12'h777;
rom[19838] = 12'h666;
rom[19839] = 12'h666;
rom[19840] = 12'h555;
rom[19841] = 12'h555;
rom[19842] = 12'h555;
rom[19843] = 12'h555;
rom[19844] = 12'h444;
rom[19845] = 12'h444;
rom[19846] = 12'h444;
rom[19847] = 12'h444;
rom[19848] = 12'h333;
rom[19849] = 12'h333;
rom[19850] = 12'h333;
rom[19851] = 12'h222;
rom[19852] = 12'h222;
rom[19853] = 12'h222;
rom[19854] = 12'h222;
rom[19855] = 12'h222;
rom[19856] = 12'h111;
rom[19857] = 12'h111;
rom[19858] = 12'h111;
rom[19859] = 12'h111;
rom[19860] = 12'h111;
rom[19861] = 12'h111;
rom[19862] = 12'h  0;
rom[19863] = 12'h  0;
rom[19864] = 12'h  0;
rom[19865] = 12'h  0;
rom[19866] = 12'h  0;
rom[19867] = 12'h  0;
rom[19868] = 12'h  0;
rom[19869] = 12'h  0;
rom[19870] = 12'h  0;
rom[19871] = 12'h  0;
rom[19872] = 12'h  0;
rom[19873] = 12'h  0;
rom[19874] = 12'h  0;
rom[19875] = 12'h  0;
rom[19876] = 12'h  0;
rom[19877] = 12'h  0;
rom[19878] = 12'h  0;
rom[19879] = 12'h  0;
rom[19880] = 12'h  0;
rom[19881] = 12'h  0;
rom[19882] = 12'h  0;
rom[19883] = 12'h  0;
rom[19884] = 12'h  0;
rom[19885] = 12'h  0;
rom[19886] = 12'h  0;
rom[19887] = 12'h  0;
rom[19888] = 12'h  0;
rom[19889] = 12'h  0;
rom[19890] = 12'h  0;
rom[19891] = 12'h  0;
rom[19892] = 12'h  0;
rom[19893] = 12'h  0;
rom[19894] = 12'h  0;
rom[19895] = 12'h111;
rom[19896] = 12'h111;
rom[19897] = 12'h111;
rom[19898] = 12'h111;
rom[19899] = 12'h111;
rom[19900] = 12'h111;
rom[19901] = 12'h111;
rom[19902] = 12'h111;
rom[19903] = 12'h111;
rom[19904] = 12'h222;
rom[19905] = 12'h222;
rom[19906] = 12'h222;
rom[19907] = 12'h333;
rom[19908] = 12'h333;
rom[19909] = 12'h333;
rom[19910] = 12'h333;
rom[19911] = 12'h333;
rom[19912] = 12'h333;
rom[19913] = 12'h333;
rom[19914] = 12'h333;
rom[19915] = 12'h333;
rom[19916] = 12'h333;
rom[19917] = 12'h333;
rom[19918] = 12'h333;
rom[19919] = 12'h333;
rom[19920] = 12'h333;
rom[19921] = 12'h333;
rom[19922] = 12'h333;
rom[19923] = 12'h333;
rom[19924] = 12'h333;
rom[19925] = 12'h444;
rom[19926] = 12'h444;
rom[19927] = 12'h444;
rom[19928] = 12'h333;
rom[19929] = 12'h333;
rom[19930] = 12'h333;
rom[19931] = 12'h333;
rom[19932] = 12'h222;
rom[19933] = 12'h222;
rom[19934] = 12'h222;
rom[19935] = 12'h222;
rom[19936] = 12'h222;
rom[19937] = 12'h222;
rom[19938] = 12'h232;
rom[19939] = 12'h232;
rom[19940] = 12'h222;
rom[19941] = 12'h222;
rom[19942] = 12'h233;
rom[19943] = 12'h333;
rom[19944] = 12'h444;
rom[19945] = 12'h444;
rom[19946] = 12'h555;
rom[19947] = 12'h655;
rom[19948] = 12'h655;
rom[19949] = 12'h555;
rom[19950] = 12'h555;
rom[19951] = 12'h555;
rom[19952] = 12'h555;
rom[19953] = 12'h555;
rom[19954] = 12'h555;
rom[19955] = 12'h555;
rom[19956] = 12'h555;
rom[19957] = 12'h555;
rom[19958] = 12'h555;
rom[19959] = 12'h555;
rom[19960] = 12'h555;
rom[19961] = 12'h455;
rom[19962] = 12'h455;
rom[19963] = 12'h455;
rom[19964] = 12'h555;
rom[19965] = 12'h555;
rom[19966] = 12'h555;
rom[19967] = 12'h555;
rom[19968] = 12'h555;
rom[19969] = 12'h555;
rom[19970] = 12'h555;
rom[19971] = 12'h555;
rom[19972] = 12'h555;
rom[19973] = 12'h555;
rom[19974] = 12'h555;
rom[19975] = 12'h555;
rom[19976] = 12'h555;
rom[19977] = 12'h555;
rom[19978] = 12'h666;
rom[19979] = 12'h666;
rom[19980] = 12'h666;
rom[19981] = 12'h666;
rom[19982] = 12'h666;
rom[19983] = 12'h666;
rom[19984] = 12'h666;
rom[19985] = 12'h666;
rom[19986] = 12'h666;
rom[19987] = 12'h777;
rom[19988] = 12'h777;
rom[19989] = 12'h777;
rom[19990] = 12'h888;
rom[19991] = 12'h888;
rom[19992] = 12'h888;
rom[19993] = 12'h888;
rom[19994] = 12'h999;
rom[19995] = 12'h999;
rom[19996] = 12'haaa;
rom[19997] = 12'haaa;
rom[19998] = 12'haaa;
rom[19999] = 12'haaa;
rom[20000] = 12'h444;
rom[20001] = 12'h444;
rom[20002] = 12'h444;
rom[20003] = 12'h444;
rom[20004] = 12'h444;
rom[20005] = 12'h555;
rom[20006] = 12'h555;
rom[20007] = 12'h555;
rom[20008] = 12'h555;
rom[20009] = 12'h555;
rom[20010] = 12'h555;
rom[20011] = 12'h555;
rom[20012] = 12'h666;
rom[20013] = 12'h666;
rom[20014] = 12'h666;
rom[20015] = 12'h666;
rom[20016] = 12'h666;
rom[20017] = 12'h666;
rom[20018] = 12'h666;
rom[20019] = 12'h777;
rom[20020] = 12'h777;
rom[20021] = 12'h777;
rom[20022] = 12'h777;
rom[20023] = 12'h777;
rom[20024] = 12'h777;
rom[20025] = 12'h777;
rom[20026] = 12'h777;
rom[20027] = 12'h777;
rom[20028] = 12'h777;
rom[20029] = 12'h777;
rom[20030] = 12'h777;
rom[20031] = 12'h777;
rom[20032] = 12'h777;
rom[20033] = 12'h777;
rom[20034] = 12'h777;
rom[20035] = 12'h666;
rom[20036] = 12'h666;
rom[20037] = 12'h666;
rom[20038] = 12'h666;
rom[20039] = 12'h666;
rom[20040] = 12'h666;
rom[20041] = 12'h666;
rom[20042] = 12'h777;
rom[20043] = 12'h777;
rom[20044] = 12'h777;
rom[20045] = 12'h777;
rom[20046] = 12'h777;
rom[20047] = 12'h777;
rom[20048] = 12'h666;
rom[20049] = 12'h777;
rom[20050] = 12'h777;
rom[20051] = 12'h777;
rom[20052] = 12'h666;
rom[20053] = 12'h666;
rom[20054] = 12'h666;
rom[20055] = 12'h666;
rom[20056] = 12'h666;
rom[20057] = 12'h666;
rom[20058] = 12'h666;
rom[20059] = 12'h555;
rom[20060] = 12'h555;
rom[20061] = 12'h666;
rom[20062] = 12'h666;
rom[20063] = 12'h666;
rom[20064] = 12'h555;
rom[20065] = 12'h555;
rom[20066] = 12'h555;
rom[20067] = 12'h555;
rom[20068] = 12'h555;
rom[20069] = 12'h555;
rom[20070] = 12'h555;
rom[20071] = 12'h555;
rom[20072] = 12'h666;
rom[20073] = 12'h666;
rom[20074] = 12'h666;
rom[20075] = 12'h666;
rom[20076] = 12'h777;
rom[20077] = 12'h777;
rom[20078] = 12'h777;
rom[20079] = 12'h888;
rom[20080] = 12'h777;
rom[20081] = 12'h777;
rom[20082] = 12'h777;
rom[20083] = 12'h777;
rom[20084] = 12'h666;
rom[20085] = 12'h666;
rom[20086] = 12'h555;
rom[20087] = 12'h555;
rom[20088] = 12'h444;
rom[20089] = 12'h333;
rom[20090] = 12'h222;
rom[20091] = 12'h222;
rom[20092] = 12'h111;
rom[20093] = 12'h111;
rom[20094] = 12'h111;
rom[20095] = 12'h  0;
rom[20096] = 12'h  0;
rom[20097] = 12'h  0;
rom[20098] = 12'h  0;
rom[20099] = 12'h  0;
rom[20100] = 12'h  0;
rom[20101] = 12'h  0;
rom[20102] = 12'h  0;
rom[20103] = 12'h  0;
rom[20104] = 12'h  0;
rom[20105] = 12'h  0;
rom[20106] = 12'h  0;
rom[20107] = 12'h  0;
rom[20108] = 12'h  0;
rom[20109] = 12'h  0;
rom[20110] = 12'h  0;
rom[20111] = 12'h  0;
rom[20112] = 12'h  0;
rom[20113] = 12'h100;
rom[20114] = 12'h100;
rom[20115] = 12'h200;
rom[20116] = 12'h200;
rom[20117] = 12'h300;
rom[20118] = 12'h510;
rom[20119] = 12'h610;
rom[20120] = 12'h710;
rom[20121] = 12'h920;
rom[20122] = 12'hb41;
rom[20123] = 12'hc41;
rom[20124] = 12'hc41;
rom[20125] = 12'hc40;
rom[20126] = 12'hc40;
rom[20127] = 12'hb40;
rom[20128] = 12'hb40;
rom[20129] = 12'ha40;
rom[20130] = 12'ha30;
rom[20131] = 12'h930;
rom[20132] = 12'h820;
rom[20133] = 12'h820;
rom[20134] = 12'h710;
rom[20135] = 12'h610;
rom[20136] = 12'h610;
rom[20137] = 12'h510;
rom[20138] = 12'h400;
rom[20139] = 12'h300;
rom[20140] = 12'h200;
rom[20141] = 12'h200;
rom[20142] = 12'h100;
rom[20143] = 12'h100;
rom[20144] = 12'h  0;
rom[20145] = 12'h  0;
rom[20146] = 12'h  0;
rom[20147] = 12'h  0;
rom[20148] = 12'h  0;
rom[20149] = 12'h  0;
rom[20150] = 12'h  0;
rom[20151] = 12'h  0;
rom[20152] = 12'h  0;
rom[20153] = 12'h  0;
rom[20154] = 12'h  0;
rom[20155] = 12'h  0;
rom[20156] = 12'h  0;
rom[20157] = 12'h  0;
rom[20158] = 12'h  0;
rom[20159] = 12'h  0;
rom[20160] = 12'h  0;
rom[20161] = 12'h  0;
rom[20162] = 12'h100;
rom[20163] = 12'h100;
rom[20164] = 12'h200;
rom[20165] = 12'h200;
rom[20166] = 12'h300;
rom[20167] = 12'h300;
rom[20168] = 12'h300;
rom[20169] = 12'h400;
rom[20170] = 12'h400;
rom[20171] = 12'h400;
rom[20172] = 12'h400;
rom[20173] = 12'h400;
rom[20174] = 12'h400;
rom[20175] = 12'h400;
rom[20176] = 12'h300;
rom[20177] = 12'h300;
rom[20178] = 12'h300;
rom[20179] = 12'h300;
rom[20180] = 12'h300;
rom[20181] = 12'h200;
rom[20182] = 12'h200;
rom[20183] = 12'h100;
rom[20184] = 12'h100;
rom[20185] = 12'h100;
rom[20186] = 12'h100;
rom[20187] = 12'h100;
rom[20188] = 12'h100;
rom[20189] = 12'h100;
rom[20190] = 12'h100;
rom[20191] = 12'h100;
rom[20192] = 12'h100;
rom[20193] = 12'h100;
rom[20194] = 12'h111;
rom[20195] = 12'h322;
rom[20196] = 12'h333;
rom[20197] = 12'h333;
rom[20198] = 12'h444;
rom[20199] = 12'h545;
rom[20200] = 12'h555;
rom[20201] = 12'h777;
rom[20202] = 12'h999;
rom[20203] = 12'hbaa;
rom[20204] = 12'hbbb;
rom[20205] = 12'hbbb;
rom[20206] = 12'hbbb;
rom[20207] = 12'hbbb;
rom[20208] = 12'haaa;
rom[20209] = 12'haaa;
rom[20210] = 12'haaa;
rom[20211] = 12'haaa;
rom[20212] = 12'haaa;
rom[20213] = 12'haaa;
rom[20214] = 12'h999;
rom[20215] = 12'h999;
rom[20216] = 12'h999;
rom[20217] = 12'h888;
rom[20218] = 12'h888;
rom[20219] = 12'h888;
rom[20220] = 12'h888;
rom[20221] = 12'h888;
rom[20222] = 12'h888;
rom[20223] = 12'h888;
rom[20224] = 12'h999;
rom[20225] = 12'h999;
rom[20226] = 12'h888;
rom[20227] = 12'h888;
rom[20228] = 12'h888;
rom[20229] = 12'h888;
rom[20230] = 12'h888;
rom[20231] = 12'h888;
rom[20232] = 12'h888;
rom[20233] = 12'h888;
rom[20234] = 12'h888;
rom[20235] = 12'h777;
rom[20236] = 12'h777;
rom[20237] = 12'h666;
rom[20238] = 12'h666;
rom[20239] = 12'h555;
rom[20240] = 12'h666;
rom[20241] = 12'h555;
rom[20242] = 12'h555;
rom[20243] = 12'h444;
rom[20244] = 12'h444;
rom[20245] = 12'h444;
rom[20246] = 12'h333;
rom[20247] = 12'h333;
rom[20248] = 12'h333;
rom[20249] = 12'h333;
rom[20250] = 12'h333;
rom[20251] = 12'h222;
rom[20252] = 12'h222;
rom[20253] = 12'h222;
rom[20254] = 12'h222;
rom[20255] = 12'h222;
rom[20256] = 12'h111;
rom[20257] = 12'h111;
rom[20258] = 12'h111;
rom[20259] = 12'h111;
rom[20260] = 12'h111;
rom[20261] = 12'h  0;
rom[20262] = 12'h  0;
rom[20263] = 12'h  0;
rom[20264] = 12'h  0;
rom[20265] = 12'h  0;
rom[20266] = 12'h  0;
rom[20267] = 12'h  0;
rom[20268] = 12'h  0;
rom[20269] = 12'h  0;
rom[20270] = 12'h  0;
rom[20271] = 12'h  0;
rom[20272] = 12'h  0;
rom[20273] = 12'h  0;
rom[20274] = 12'h  0;
rom[20275] = 12'h  0;
rom[20276] = 12'h  0;
rom[20277] = 12'h  0;
rom[20278] = 12'h  0;
rom[20279] = 12'h  0;
rom[20280] = 12'h  0;
rom[20281] = 12'h  0;
rom[20282] = 12'h  0;
rom[20283] = 12'h  0;
rom[20284] = 12'h  0;
rom[20285] = 12'h  0;
rom[20286] = 12'h  0;
rom[20287] = 12'h  0;
rom[20288] = 12'h  0;
rom[20289] = 12'h  0;
rom[20290] = 12'h  0;
rom[20291] = 12'h  0;
rom[20292] = 12'h  0;
rom[20293] = 12'h  0;
rom[20294] = 12'h  0;
rom[20295] = 12'h111;
rom[20296] = 12'h111;
rom[20297] = 12'h111;
rom[20298] = 12'h111;
rom[20299] = 12'h111;
rom[20300] = 12'h111;
rom[20301] = 12'h111;
rom[20302] = 12'h111;
rom[20303] = 12'h111;
rom[20304] = 12'h222;
rom[20305] = 12'h222;
rom[20306] = 12'h333;
rom[20307] = 12'h333;
rom[20308] = 12'h333;
rom[20309] = 12'h222;
rom[20310] = 12'h333;
rom[20311] = 12'h333;
rom[20312] = 12'h333;
rom[20313] = 12'h333;
rom[20314] = 12'h333;
rom[20315] = 12'h333;
rom[20316] = 12'h333;
rom[20317] = 12'h333;
rom[20318] = 12'h222;
rom[20319] = 12'h333;
rom[20320] = 12'h333;
rom[20321] = 12'h333;
rom[20322] = 12'h333;
rom[20323] = 12'h333;
rom[20324] = 12'h444;
rom[20325] = 12'h444;
rom[20326] = 12'h444;
rom[20327] = 12'h444;
rom[20328] = 12'h333;
rom[20329] = 12'h333;
rom[20330] = 12'h333;
rom[20331] = 12'h333;
rom[20332] = 12'h333;
rom[20333] = 12'h333;
rom[20334] = 12'h222;
rom[20335] = 12'h222;
rom[20336] = 12'h222;
rom[20337] = 12'h222;
rom[20338] = 12'h222;
rom[20339] = 12'h222;
rom[20340] = 12'h222;
rom[20341] = 12'h222;
rom[20342] = 12'h333;
rom[20343] = 12'h333;
rom[20344] = 12'h555;
rom[20345] = 12'h555;
rom[20346] = 12'h655;
rom[20347] = 12'h666;
rom[20348] = 12'h665;
rom[20349] = 12'h555;
rom[20350] = 12'h555;
rom[20351] = 12'h555;
rom[20352] = 12'h444;
rom[20353] = 12'h555;
rom[20354] = 12'h555;
rom[20355] = 12'h555;
rom[20356] = 12'h555;
rom[20357] = 12'h555;
rom[20358] = 12'h555;
rom[20359] = 12'h555;
rom[20360] = 12'h555;
rom[20361] = 12'h555;
rom[20362] = 12'h555;
rom[20363] = 12'h555;
rom[20364] = 12'h555;
rom[20365] = 12'h555;
rom[20366] = 12'h555;
rom[20367] = 12'h555;
rom[20368] = 12'h555;
rom[20369] = 12'h555;
rom[20370] = 12'h555;
rom[20371] = 12'h555;
rom[20372] = 12'h555;
rom[20373] = 12'h555;
rom[20374] = 12'h555;
rom[20375] = 12'h555;
rom[20376] = 12'h555;
rom[20377] = 12'h555;
rom[20378] = 12'h555;
rom[20379] = 12'h666;
rom[20380] = 12'h666;
rom[20381] = 12'h666;
rom[20382] = 12'h666;
rom[20383] = 12'h666;
rom[20384] = 12'h666;
rom[20385] = 12'h666;
rom[20386] = 12'h666;
rom[20387] = 12'h777;
rom[20388] = 12'h777;
rom[20389] = 12'h777;
rom[20390] = 12'h888;
rom[20391] = 12'h888;
rom[20392] = 12'h888;
rom[20393] = 12'h888;
rom[20394] = 12'h999;
rom[20395] = 12'h999;
rom[20396] = 12'haaa;
rom[20397] = 12'haaa;
rom[20398] = 12'haaa;
rom[20399] = 12'haaa;
rom[20400] = 12'h555;
rom[20401] = 12'h555;
rom[20402] = 12'h555;
rom[20403] = 12'h555;
rom[20404] = 12'h555;
rom[20405] = 12'h555;
rom[20406] = 12'h555;
rom[20407] = 12'h555;
rom[20408] = 12'h666;
rom[20409] = 12'h666;
rom[20410] = 12'h666;
rom[20411] = 12'h666;
rom[20412] = 12'h666;
rom[20413] = 12'h666;
rom[20414] = 12'h777;
rom[20415] = 12'h777;
rom[20416] = 12'h777;
rom[20417] = 12'h777;
rom[20418] = 12'h777;
rom[20419] = 12'h777;
rom[20420] = 12'h777;
rom[20421] = 12'h777;
rom[20422] = 12'h777;
rom[20423] = 12'h888;
rom[20424] = 12'h777;
rom[20425] = 12'h777;
rom[20426] = 12'h777;
rom[20427] = 12'h777;
rom[20428] = 12'h777;
rom[20429] = 12'h777;
rom[20430] = 12'h666;
rom[20431] = 12'h666;
rom[20432] = 12'h777;
rom[20433] = 12'h777;
rom[20434] = 12'h666;
rom[20435] = 12'h666;
rom[20436] = 12'h666;
rom[20437] = 12'h666;
rom[20438] = 12'h666;
rom[20439] = 12'h666;
rom[20440] = 12'h666;
rom[20441] = 12'h666;
rom[20442] = 12'h666;
rom[20443] = 12'h777;
rom[20444] = 12'h777;
rom[20445] = 12'h777;
rom[20446] = 12'h777;
rom[20447] = 12'h777;
rom[20448] = 12'h777;
rom[20449] = 12'h777;
rom[20450] = 12'h777;
rom[20451] = 12'h777;
rom[20452] = 12'h777;
rom[20453] = 12'h666;
rom[20454] = 12'h666;
rom[20455] = 12'h666;
rom[20456] = 12'h666;
rom[20457] = 12'h666;
rom[20458] = 12'h666;
rom[20459] = 12'h555;
rom[20460] = 12'h555;
rom[20461] = 12'h555;
rom[20462] = 12'h555;
rom[20463] = 12'h555;
rom[20464] = 12'h555;
rom[20465] = 12'h555;
rom[20466] = 12'h555;
rom[20467] = 12'h555;
rom[20468] = 12'h555;
rom[20469] = 12'h555;
rom[20470] = 12'h555;
rom[20471] = 12'h555;
rom[20472] = 12'h666;
rom[20473] = 12'h666;
rom[20474] = 12'h666;
rom[20475] = 12'h666;
rom[20476] = 12'h666;
rom[20477] = 12'h666;
rom[20478] = 12'h777;
rom[20479] = 12'h777;
rom[20480] = 12'h777;
rom[20481] = 12'h777;
rom[20482] = 12'h777;
rom[20483] = 12'h777;
rom[20484] = 12'h777;
rom[20485] = 12'h666;
rom[20486] = 12'h555;
rom[20487] = 12'h555;
rom[20488] = 12'h444;
rom[20489] = 12'h333;
rom[20490] = 12'h333;
rom[20491] = 12'h222;
rom[20492] = 12'h111;
rom[20493] = 12'h111;
rom[20494] = 12'h111;
rom[20495] = 12'h  0;
rom[20496] = 12'h  0;
rom[20497] = 12'h  0;
rom[20498] = 12'h  0;
rom[20499] = 12'h  0;
rom[20500] = 12'h  0;
rom[20501] = 12'h  0;
rom[20502] = 12'h  0;
rom[20503] = 12'h  0;
rom[20504] = 12'h  0;
rom[20505] = 12'h  0;
rom[20506] = 12'h  0;
rom[20507] = 12'h  0;
rom[20508] = 12'h  0;
rom[20509] = 12'h  0;
rom[20510] = 12'h  0;
rom[20511] = 12'h  0;
rom[20512] = 12'h  0;
rom[20513] = 12'h100;
rom[20514] = 12'h100;
rom[20515] = 12'h200;
rom[20516] = 12'h200;
rom[20517] = 12'h300;
rom[20518] = 12'h510;
rom[20519] = 12'h610;
rom[20520] = 12'h710;
rom[20521] = 12'h920;
rom[20522] = 12'hb41;
rom[20523] = 12'hc51;
rom[20524] = 12'hd51;
rom[20525] = 12'hd51;
rom[20526] = 12'hc40;
rom[20527] = 12'hc40;
rom[20528] = 12'hb40;
rom[20529] = 12'hb40;
rom[20530] = 12'hb40;
rom[20531] = 12'ha30;
rom[20532] = 12'h930;
rom[20533] = 12'h820;
rom[20534] = 12'h820;
rom[20535] = 12'h720;
rom[20536] = 12'h610;
rom[20537] = 12'h510;
rom[20538] = 12'h400;
rom[20539] = 12'h300;
rom[20540] = 12'h200;
rom[20541] = 12'h200;
rom[20542] = 12'h100;
rom[20543] = 12'h100;
rom[20544] = 12'h  0;
rom[20545] = 12'h  0;
rom[20546] = 12'h  0;
rom[20547] = 12'h  0;
rom[20548] = 12'h  0;
rom[20549] = 12'h  0;
rom[20550] = 12'h  0;
rom[20551] = 12'h  0;
rom[20552] = 12'h  0;
rom[20553] = 12'h  0;
rom[20554] = 12'h  0;
rom[20555] = 12'h  0;
rom[20556] = 12'h  0;
rom[20557] = 12'h  0;
rom[20558] = 12'h  0;
rom[20559] = 12'h  0;
rom[20560] = 12'h  0;
rom[20561] = 12'h  0;
rom[20562] = 12'h100;
rom[20563] = 12'h100;
rom[20564] = 12'h200;
rom[20565] = 12'h200;
rom[20566] = 12'h300;
rom[20567] = 12'h300;
rom[20568] = 12'h400;
rom[20569] = 12'h400;
rom[20570] = 12'h400;
rom[20571] = 12'h400;
rom[20572] = 12'h400;
rom[20573] = 12'h400;
rom[20574] = 12'h400;
rom[20575] = 12'h400;
rom[20576] = 12'h300;
rom[20577] = 12'h300;
rom[20578] = 12'h300;
rom[20579] = 12'h300;
rom[20580] = 12'h200;
rom[20581] = 12'h200;
rom[20582] = 12'h200;
rom[20583] = 12'h100;
rom[20584] = 12'h100;
rom[20585] = 12'h100;
rom[20586] = 12'h100;
rom[20587] = 12'h100;
rom[20588] = 12'h100;
rom[20589] = 12'h  0;
rom[20590] = 12'h100;
rom[20591] = 12'h100;
rom[20592] = 12'h100;
rom[20593] = 12'h100;
rom[20594] = 12'h111;
rom[20595] = 12'h222;
rom[20596] = 12'h333;
rom[20597] = 12'h433;
rom[20598] = 12'h444;
rom[20599] = 12'h555;
rom[20600] = 12'h555;
rom[20601] = 12'h766;
rom[20602] = 12'h988;
rom[20603] = 12'haaa;
rom[20604] = 12'hbbb;
rom[20605] = 12'hbbb;
rom[20606] = 12'hbbb;
rom[20607] = 12'hbbb;
rom[20608] = 12'haaa;
rom[20609] = 12'haaa;
rom[20610] = 12'haaa;
rom[20611] = 12'haaa;
rom[20612] = 12'haaa;
rom[20613] = 12'haaa;
rom[20614] = 12'haaa;
rom[20615] = 12'h999;
rom[20616] = 12'h999;
rom[20617] = 12'h999;
rom[20618] = 12'h888;
rom[20619] = 12'h888;
rom[20620] = 12'h888;
rom[20621] = 12'h888;
rom[20622] = 12'h888;
rom[20623] = 12'h888;
rom[20624] = 12'h999;
rom[20625] = 12'h999;
rom[20626] = 12'h888;
rom[20627] = 12'h888;
rom[20628] = 12'h888;
rom[20629] = 12'h888;
rom[20630] = 12'h888;
rom[20631] = 12'h888;
rom[20632] = 12'h888;
rom[20633] = 12'h888;
rom[20634] = 12'h777;
rom[20635] = 12'h777;
rom[20636] = 12'h777;
rom[20637] = 12'h666;
rom[20638] = 12'h666;
rom[20639] = 12'h555;
rom[20640] = 12'h666;
rom[20641] = 12'h555;
rom[20642] = 12'h555;
rom[20643] = 12'h444;
rom[20644] = 12'h444;
rom[20645] = 12'h333;
rom[20646] = 12'h333;
rom[20647] = 12'h333;
rom[20648] = 12'h333;
rom[20649] = 12'h333;
rom[20650] = 12'h333;
rom[20651] = 12'h333;
rom[20652] = 12'h333;
rom[20653] = 12'h222;
rom[20654] = 12'h222;
rom[20655] = 12'h111;
rom[20656] = 12'h111;
rom[20657] = 12'h111;
rom[20658] = 12'h111;
rom[20659] = 12'h111;
rom[20660] = 12'h  0;
rom[20661] = 12'h  0;
rom[20662] = 12'h  0;
rom[20663] = 12'h  0;
rom[20664] = 12'h111;
rom[20665] = 12'h111;
rom[20666] = 12'h111;
rom[20667] = 12'h  0;
rom[20668] = 12'h  0;
rom[20669] = 12'h  0;
rom[20670] = 12'h  0;
rom[20671] = 12'h  0;
rom[20672] = 12'h  0;
rom[20673] = 12'h  0;
rom[20674] = 12'h  0;
rom[20675] = 12'h  0;
rom[20676] = 12'h  0;
rom[20677] = 12'h  0;
rom[20678] = 12'h  0;
rom[20679] = 12'h  0;
rom[20680] = 12'h  0;
rom[20681] = 12'h  0;
rom[20682] = 12'h  0;
rom[20683] = 12'h  0;
rom[20684] = 12'h  0;
rom[20685] = 12'h  0;
rom[20686] = 12'h  0;
rom[20687] = 12'h  0;
rom[20688] = 12'h  0;
rom[20689] = 12'h  0;
rom[20690] = 12'h  0;
rom[20691] = 12'h  0;
rom[20692] = 12'h  0;
rom[20693] = 12'h  0;
rom[20694] = 12'h111;
rom[20695] = 12'h111;
rom[20696] = 12'h111;
rom[20697] = 12'h111;
rom[20698] = 12'h111;
rom[20699] = 12'h111;
rom[20700] = 12'h111;
rom[20701] = 12'h111;
rom[20702] = 12'h111;
rom[20703] = 12'h111;
rom[20704] = 12'h222;
rom[20705] = 12'h222;
rom[20706] = 12'h333;
rom[20707] = 12'h333;
rom[20708] = 12'h222;
rom[20709] = 12'h222;
rom[20710] = 12'h333;
rom[20711] = 12'h333;
rom[20712] = 12'h333;
rom[20713] = 12'h333;
rom[20714] = 12'h333;
rom[20715] = 12'h333;
rom[20716] = 12'h333;
rom[20717] = 12'h333;
rom[20718] = 12'h222;
rom[20719] = 12'h333;
rom[20720] = 12'h333;
rom[20721] = 12'h333;
rom[20722] = 12'h333;
rom[20723] = 12'h333;
rom[20724] = 12'h333;
rom[20725] = 12'h444;
rom[20726] = 12'h444;
rom[20727] = 12'h444;
rom[20728] = 12'h333;
rom[20729] = 12'h333;
rom[20730] = 12'h333;
rom[20731] = 12'h333;
rom[20732] = 12'h333;
rom[20733] = 12'h333;
rom[20734] = 12'h333;
rom[20735] = 12'h233;
rom[20736] = 12'h233;
rom[20737] = 12'h232;
rom[20738] = 12'h222;
rom[20739] = 12'h222;
rom[20740] = 12'h233;
rom[20741] = 12'h333;
rom[20742] = 12'h444;
rom[20743] = 12'h444;
rom[20744] = 12'h555;
rom[20745] = 12'h555;
rom[20746] = 12'h666;
rom[20747] = 12'h666;
rom[20748] = 12'h666;
rom[20749] = 12'h555;
rom[20750] = 12'h555;
rom[20751] = 12'h555;
rom[20752] = 12'h555;
rom[20753] = 12'h555;
rom[20754] = 12'h555;
rom[20755] = 12'h555;
rom[20756] = 12'h555;
rom[20757] = 12'h555;
rom[20758] = 12'h555;
rom[20759] = 12'h555;
rom[20760] = 12'h555;
rom[20761] = 12'h555;
rom[20762] = 12'h555;
rom[20763] = 12'h555;
rom[20764] = 12'h555;
rom[20765] = 12'h555;
rom[20766] = 12'h555;
rom[20767] = 12'h555;
rom[20768] = 12'h555;
rom[20769] = 12'h555;
rom[20770] = 12'h555;
rom[20771] = 12'h555;
rom[20772] = 12'h555;
rom[20773] = 12'h555;
rom[20774] = 12'h555;
rom[20775] = 12'h555;
rom[20776] = 12'h555;
rom[20777] = 12'h555;
rom[20778] = 12'h555;
rom[20779] = 12'h666;
rom[20780] = 12'h666;
rom[20781] = 12'h666;
rom[20782] = 12'h666;
rom[20783] = 12'h666;
rom[20784] = 12'h666;
rom[20785] = 12'h666;
rom[20786] = 12'h777;
rom[20787] = 12'h777;
rom[20788] = 12'h777;
rom[20789] = 12'h777;
rom[20790] = 12'h888;
rom[20791] = 12'h888;
rom[20792] = 12'h888;
rom[20793] = 12'h888;
rom[20794] = 12'h999;
rom[20795] = 12'h999;
rom[20796] = 12'haaa;
rom[20797] = 12'haaa;
rom[20798] = 12'haaa;
rom[20799] = 12'haaa;
rom[20800] = 12'h555;
rom[20801] = 12'h555;
rom[20802] = 12'h555;
rom[20803] = 12'h555;
rom[20804] = 12'h555;
rom[20805] = 12'h555;
rom[20806] = 12'h555;
rom[20807] = 12'h555;
rom[20808] = 12'h666;
rom[20809] = 12'h666;
rom[20810] = 12'h666;
rom[20811] = 12'h666;
rom[20812] = 12'h777;
rom[20813] = 12'h777;
rom[20814] = 12'h777;
rom[20815] = 12'h777;
rom[20816] = 12'h777;
rom[20817] = 12'h777;
rom[20818] = 12'h777;
rom[20819] = 12'h777;
rom[20820] = 12'h777;
rom[20821] = 12'h777;
rom[20822] = 12'h777;
rom[20823] = 12'h777;
rom[20824] = 12'h777;
rom[20825] = 12'h777;
rom[20826] = 12'h777;
rom[20827] = 12'h777;
rom[20828] = 12'h777;
rom[20829] = 12'h666;
rom[20830] = 12'h666;
rom[20831] = 12'h666;
rom[20832] = 12'h777;
rom[20833] = 12'h777;
rom[20834] = 12'h777;
rom[20835] = 12'h777;
rom[20836] = 12'h666;
rom[20837] = 12'h666;
rom[20838] = 12'h666;
rom[20839] = 12'h666;
rom[20840] = 12'h666;
rom[20841] = 12'h666;
rom[20842] = 12'h666;
rom[20843] = 12'h777;
rom[20844] = 12'h777;
rom[20845] = 12'h777;
rom[20846] = 12'h777;
rom[20847] = 12'h777;
rom[20848] = 12'h777;
rom[20849] = 12'h666;
rom[20850] = 12'h666;
rom[20851] = 12'h666;
rom[20852] = 12'h666;
rom[20853] = 12'h666;
rom[20854] = 12'h666;
rom[20855] = 12'h666;
rom[20856] = 12'h666;
rom[20857] = 12'h666;
rom[20858] = 12'h666;
rom[20859] = 12'h666;
rom[20860] = 12'h555;
rom[20861] = 12'h555;
rom[20862] = 12'h555;
rom[20863] = 12'h555;
rom[20864] = 12'h555;
rom[20865] = 12'h555;
rom[20866] = 12'h555;
rom[20867] = 12'h555;
rom[20868] = 12'h555;
rom[20869] = 12'h555;
rom[20870] = 12'h555;
rom[20871] = 12'h555;
rom[20872] = 12'h666;
rom[20873] = 12'h666;
rom[20874] = 12'h666;
rom[20875] = 12'h666;
rom[20876] = 12'h666;
rom[20877] = 12'h666;
rom[20878] = 12'h666;
rom[20879] = 12'h777;
rom[20880] = 12'h777;
rom[20881] = 12'h777;
rom[20882] = 12'h777;
rom[20883] = 12'h777;
rom[20884] = 12'h777;
rom[20885] = 12'h666;
rom[20886] = 12'h555;
rom[20887] = 12'h555;
rom[20888] = 12'h444;
rom[20889] = 12'h444;
rom[20890] = 12'h333;
rom[20891] = 12'h222;
rom[20892] = 12'h111;
rom[20893] = 12'h111;
rom[20894] = 12'h111;
rom[20895] = 12'h111;
rom[20896] = 12'h  0;
rom[20897] = 12'h  0;
rom[20898] = 12'h  0;
rom[20899] = 12'h  0;
rom[20900] = 12'h  0;
rom[20901] = 12'h  0;
rom[20902] = 12'h  0;
rom[20903] = 12'h  0;
rom[20904] = 12'h  0;
rom[20905] = 12'h  0;
rom[20906] = 12'h  0;
rom[20907] = 12'h  0;
rom[20908] = 12'h  0;
rom[20909] = 12'h  0;
rom[20910] = 12'h  0;
rom[20911] = 12'h  0;
rom[20912] = 12'h  0;
rom[20913] = 12'h100;
rom[20914] = 12'h100;
rom[20915] = 12'h200;
rom[20916] = 12'h200;
rom[20917] = 12'h300;
rom[20918] = 12'h510;
rom[20919] = 12'h610;
rom[20920] = 12'h710;
rom[20921] = 12'h820;
rom[20922] = 12'ha30;
rom[20923] = 12'hc51;
rom[20924] = 12'hd51;
rom[20925] = 12'hd51;
rom[20926] = 12'hd51;
rom[20927] = 12'hd50;
rom[20928] = 12'hc40;
rom[20929] = 12'hc40;
rom[20930] = 12'hb40;
rom[20931] = 12'hb30;
rom[20932] = 12'ha30;
rom[20933] = 12'h930;
rom[20934] = 12'h920;
rom[20935] = 12'h820;
rom[20936] = 12'h710;
rom[20937] = 12'h510;
rom[20938] = 12'h400;
rom[20939] = 12'h300;
rom[20940] = 12'h200;
rom[20941] = 12'h200;
rom[20942] = 12'h100;
rom[20943] = 12'h100;
rom[20944] = 12'h  0;
rom[20945] = 12'h  0;
rom[20946] = 12'h  0;
rom[20947] = 12'h  0;
rom[20948] = 12'h  0;
rom[20949] = 12'h  0;
rom[20950] = 12'h  0;
rom[20951] = 12'h  0;
rom[20952] = 12'h  0;
rom[20953] = 12'h  0;
rom[20954] = 12'h  0;
rom[20955] = 12'h  0;
rom[20956] = 12'h  0;
rom[20957] = 12'h  0;
rom[20958] = 12'h  0;
rom[20959] = 12'h  0;
rom[20960] = 12'h  0;
rom[20961] = 12'h  0;
rom[20962] = 12'h100;
rom[20963] = 12'h100;
rom[20964] = 12'h200;
rom[20965] = 12'h200;
rom[20966] = 12'h300;
rom[20967] = 12'h300;
rom[20968] = 12'h400;
rom[20969] = 12'h400;
rom[20970] = 12'h400;
rom[20971] = 12'h400;
rom[20972] = 12'h400;
rom[20973] = 12'h400;
rom[20974] = 12'h400;
rom[20975] = 12'h400;
rom[20976] = 12'h300;
rom[20977] = 12'h300;
rom[20978] = 12'h300;
rom[20979] = 12'h300;
rom[20980] = 12'h200;
rom[20981] = 12'h200;
rom[20982] = 12'h100;
rom[20983] = 12'h100;
rom[20984] = 12'h100;
rom[20985] = 12'h100;
rom[20986] = 12'h100;
rom[20987] = 12'h100;
rom[20988] = 12'h  0;
rom[20989] = 12'h  0;
rom[20990] = 12'h  0;
rom[20991] = 12'h  0;
rom[20992] = 12'h100;
rom[20993] = 12'h100;
rom[20994] = 12'h111;
rom[20995] = 12'h222;
rom[20996] = 12'h333;
rom[20997] = 12'h444;
rom[20998] = 12'h544;
rom[20999] = 12'h555;
rom[21000] = 12'h555;
rom[21001] = 12'h666;
rom[21002] = 12'h888;
rom[21003] = 12'haaa;
rom[21004] = 12'hbbb;
rom[21005] = 12'hbbb;
rom[21006] = 12'hbbb;
rom[21007] = 12'hbbb;
rom[21008] = 12'hbbb;
rom[21009] = 12'haaa;
rom[21010] = 12'haaa;
rom[21011] = 12'haaa;
rom[21012] = 12'haaa;
rom[21013] = 12'haaa;
rom[21014] = 12'haaa;
rom[21015] = 12'h999;
rom[21016] = 12'h999;
rom[21017] = 12'h999;
rom[21018] = 12'h999;
rom[21019] = 12'h888;
rom[21020] = 12'h999;
rom[21021] = 12'h999;
rom[21022] = 12'h999;
rom[21023] = 12'h999;
rom[21024] = 12'h999;
rom[21025] = 12'h999;
rom[21026] = 12'h888;
rom[21027] = 12'h888;
rom[21028] = 12'h888;
rom[21029] = 12'h888;
rom[21030] = 12'h888;
rom[21031] = 12'h888;
rom[21032] = 12'h777;
rom[21033] = 12'h777;
rom[21034] = 12'h777;
rom[21035] = 12'h777;
rom[21036] = 12'h666;
rom[21037] = 12'h666;
rom[21038] = 12'h666;
rom[21039] = 12'h666;
rom[21040] = 12'h555;
rom[21041] = 12'h555;
rom[21042] = 12'h444;
rom[21043] = 12'h444;
rom[21044] = 12'h444;
rom[21045] = 12'h333;
rom[21046] = 12'h333;
rom[21047] = 12'h333;
rom[21048] = 12'h333;
rom[21049] = 12'h333;
rom[21050] = 12'h333;
rom[21051] = 12'h333;
rom[21052] = 12'h333;
rom[21053] = 12'h222;
rom[21054] = 12'h111;
rom[21055] = 12'h111;
rom[21056] = 12'h111;
rom[21057] = 12'h111;
rom[21058] = 12'h111;
rom[21059] = 12'h  0;
rom[21060] = 12'h  0;
rom[21061] = 12'h  0;
rom[21062] = 12'h  0;
rom[21063] = 12'h111;
rom[21064] = 12'h111;
rom[21065] = 12'h111;
rom[21066] = 12'h111;
rom[21067] = 12'h  0;
rom[21068] = 12'h  0;
rom[21069] = 12'h  0;
rom[21070] = 12'h  0;
rom[21071] = 12'h  0;
rom[21072] = 12'h  0;
rom[21073] = 12'h  0;
rom[21074] = 12'h  0;
rom[21075] = 12'h  0;
rom[21076] = 12'h  0;
rom[21077] = 12'h  0;
rom[21078] = 12'h  0;
rom[21079] = 12'h  0;
rom[21080] = 12'h  0;
rom[21081] = 12'h  0;
rom[21082] = 12'h  0;
rom[21083] = 12'h  0;
rom[21084] = 12'h  0;
rom[21085] = 12'h  0;
rom[21086] = 12'h  0;
rom[21087] = 12'h  0;
rom[21088] = 12'h  0;
rom[21089] = 12'h  0;
rom[21090] = 12'h  0;
rom[21091] = 12'h  0;
rom[21092] = 12'h  0;
rom[21093] = 12'h  0;
rom[21094] = 12'h111;
rom[21095] = 12'h111;
rom[21096] = 12'h111;
rom[21097] = 12'h111;
rom[21098] = 12'h111;
rom[21099] = 12'h111;
rom[21100] = 12'h111;
rom[21101] = 12'h111;
rom[21102] = 12'h111;
rom[21103] = 12'h222;
rom[21104] = 12'h222;
rom[21105] = 12'h333;
rom[21106] = 12'h333;
rom[21107] = 12'h333;
rom[21108] = 12'h222;
rom[21109] = 12'h333;
rom[21110] = 12'h333;
rom[21111] = 12'h333;
rom[21112] = 12'h333;
rom[21113] = 12'h333;
rom[21114] = 12'h333;
rom[21115] = 12'h333;
rom[21116] = 12'h333;
rom[21117] = 12'h333;
rom[21118] = 12'h333;
rom[21119] = 12'h333;
rom[21120] = 12'h333;
rom[21121] = 12'h333;
rom[21122] = 12'h333;
rom[21123] = 12'h333;
rom[21124] = 12'h333;
rom[21125] = 12'h444;
rom[21126] = 12'h444;
rom[21127] = 12'h333;
rom[21128] = 12'h333;
rom[21129] = 12'h333;
rom[21130] = 12'h333;
rom[21131] = 12'h333;
rom[21132] = 12'h333;
rom[21133] = 12'h333;
rom[21134] = 12'h333;
rom[21135] = 12'h333;
rom[21136] = 12'h333;
rom[21137] = 12'h233;
rom[21138] = 12'h232;
rom[21139] = 12'h333;
rom[21140] = 12'h333;
rom[21141] = 12'h444;
rom[21142] = 12'h444;
rom[21143] = 12'h555;
rom[21144] = 12'h555;
rom[21145] = 12'h666;
rom[21146] = 12'h666;
rom[21147] = 12'h666;
rom[21148] = 12'h666;
rom[21149] = 12'h555;
rom[21150] = 12'h555;
rom[21151] = 12'h554;
rom[21152] = 12'h544;
rom[21153] = 12'h555;
rom[21154] = 12'h555;
rom[21155] = 12'h555;
rom[21156] = 12'h555;
rom[21157] = 12'h555;
rom[21158] = 12'h555;
rom[21159] = 12'h555;
rom[21160] = 12'h555;
rom[21161] = 12'h555;
rom[21162] = 12'h555;
rom[21163] = 12'h555;
rom[21164] = 12'h666;
rom[21165] = 12'h666;
rom[21166] = 12'h666;
rom[21167] = 12'h666;
rom[21168] = 12'h666;
rom[21169] = 12'h666;
rom[21170] = 12'h666;
rom[21171] = 12'h666;
rom[21172] = 12'h666;
rom[21173] = 12'h666;
rom[21174] = 12'h666;
rom[21175] = 12'h666;
rom[21176] = 12'h666;
rom[21177] = 12'h666;
rom[21178] = 12'h666;
rom[21179] = 12'h666;
rom[21180] = 12'h666;
rom[21181] = 12'h666;
rom[21182] = 12'h666;
rom[21183] = 12'h777;
rom[21184] = 12'h777;
rom[21185] = 12'h777;
rom[21186] = 12'h777;
rom[21187] = 12'h777;
rom[21188] = 12'h777;
rom[21189] = 12'h777;
rom[21190] = 12'h777;
rom[21191] = 12'h888;
rom[21192] = 12'h888;
rom[21193] = 12'h888;
rom[21194] = 12'h999;
rom[21195] = 12'h999;
rom[21196] = 12'haaa;
rom[21197] = 12'haaa;
rom[21198] = 12'haaa;
rom[21199] = 12'haaa;
rom[21200] = 12'h555;
rom[21201] = 12'h555;
rom[21202] = 12'h555;
rom[21203] = 12'h555;
rom[21204] = 12'h555;
rom[21205] = 12'h666;
rom[21206] = 12'h666;
rom[21207] = 12'h666;
rom[21208] = 12'h666;
rom[21209] = 12'h666;
rom[21210] = 12'h777;
rom[21211] = 12'h777;
rom[21212] = 12'h777;
rom[21213] = 12'h777;
rom[21214] = 12'h777;
rom[21215] = 12'h777;
rom[21216] = 12'h777;
rom[21217] = 12'h777;
rom[21218] = 12'h777;
rom[21219] = 12'h777;
rom[21220] = 12'h666;
rom[21221] = 12'h666;
rom[21222] = 12'h666;
rom[21223] = 12'h666;
rom[21224] = 12'h666;
rom[21225] = 12'h666;
rom[21226] = 12'h666;
rom[21227] = 12'h666;
rom[21228] = 12'h666;
rom[21229] = 12'h666;
rom[21230] = 12'h666;
rom[21231] = 12'h666;
rom[21232] = 12'h777;
rom[21233] = 12'h777;
rom[21234] = 12'h777;
rom[21235] = 12'h777;
rom[21236] = 12'h777;
rom[21237] = 12'h777;
rom[21238] = 12'h777;
rom[21239] = 12'h777;
rom[21240] = 12'h666;
rom[21241] = 12'h777;
rom[21242] = 12'h777;
rom[21243] = 12'h777;
rom[21244] = 12'h777;
rom[21245] = 12'h777;
rom[21246] = 12'h777;
rom[21247] = 12'h777;
rom[21248] = 12'h777;
rom[21249] = 12'h666;
rom[21250] = 12'h666;
rom[21251] = 12'h666;
rom[21252] = 12'h666;
rom[21253] = 12'h666;
rom[21254] = 12'h666;
rom[21255] = 12'h666;
rom[21256] = 12'h666;
rom[21257] = 12'h666;
rom[21258] = 12'h666;
rom[21259] = 12'h666;
rom[21260] = 12'h666;
rom[21261] = 12'h555;
rom[21262] = 12'h555;
rom[21263] = 12'h555;
rom[21264] = 12'h555;
rom[21265] = 12'h555;
rom[21266] = 12'h555;
rom[21267] = 12'h555;
rom[21268] = 12'h555;
rom[21269] = 12'h666;
rom[21270] = 12'h666;
rom[21271] = 12'h666;
rom[21272] = 12'h666;
rom[21273] = 12'h666;
rom[21274] = 12'h666;
rom[21275] = 12'h555;
rom[21276] = 12'h555;
rom[21277] = 12'h555;
rom[21278] = 12'h666;
rom[21279] = 12'h666;
rom[21280] = 12'h777;
rom[21281] = 12'h777;
rom[21282] = 12'h777;
rom[21283] = 12'h777;
rom[21284] = 12'h777;
rom[21285] = 12'h777;
rom[21286] = 12'h666;
rom[21287] = 12'h555;
rom[21288] = 12'h444;
rom[21289] = 12'h444;
rom[21290] = 12'h333;
rom[21291] = 12'h222;
rom[21292] = 12'h222;
rom[21293] = 12'h111;
rom[21294] = 12'h111;
rom[21295] = 12'h111;
rom[21296] = 12'h  0;
rom[21297] = 12'h  0;
rom[21298] = 12'h  0;
rom[21299] = 12'h  0;
rom[21300] = 12'h  0;
rom[21301] = 12'h  0;
rom[21302] = 12'h  0;
rom[21303] = 12'h  0;
rom[21304] = 12'h  0;
rom[21305] = 12'h  0;
rom[21306] = 12'h  0;
rom[21307] = 12'h  0;
rom[21308] = 12'h  0;
rom[21309] = 12'h  0;
rom[21310] = 12'h  0;
rom[21311] = 12'h  0;
rom[21312] = 12'h100;
rom[21313] = 12'h100;
rom[21314] = 12'h100;
rom[21315] = 12'h200;
rom[21316] = 12'h200;
rom[21317] = 12'h300;
rom[21318] = 12'h410;
rom[21319] = 12'h510;
rom[21320] = 12'h710;
rom[21321] = 12'h820;
rom[21322] = 12'ha30;
rom[21323] = 12'hb41;
rom[21324] = 12'hc51;
rom[21325] = 12'hd61;
rom[21326] = 12'hd51;
rom[21327] = 12'hd51;
rom[21328] = 12'hd50;
rom[21329] = 12'hd40;
rom[21330] = 12'hc40;
rom[21331] = 12'hc40;
rom[21332] = 12'hb30;
rom[21333] = 12'ha30;
rom[21334] = 12'h920;
rom[21335] = 12'h920;
rom[21336] = 12'h710;
rom[21337] = 12'h610;
rom[21338] = 12'h500;
rom[21339] = 12'h300;
rom[21340] = 12'h300;
rom[21341] = 12'h200;
rom[21342] = 12'h100;
rom[21343] = 12'h100;
rom[21344] = 12'h  0;
rom[21345] = 12'h  0;
rom[21346] = 12'h  0;
rom[21347] = 12'h  0;
rom[21348] = 12'h  0;
rom[21349] = 12'h  0;
rom[21350] = 12'h  0;
rom[21351] = 12'h  0;
rom[21352] = 12'h  0;
rom[21353] = 12'h  0;
rom[21354] = 12'h  0;
rom[21355] = 12'h  0;
rom[21356] = 12'h  0;
rom[21357] = 12'h  0;
rom[21358] = 12'h  0;
rom[21359] = 12'h  0;
rom[21360] = 12'h  0;
rom[21361] = 12'h100;
rom[21362] = 12'h100;
rom[21363] = 12'h200;
rom[21364] = 12'h200;
rom[21365] = 12'h300;
rom[21366] = 12'h300;
rom[21367] = 12'h400;
rom[21368] = 12'h400;
rom[21369] = 12'h400;
rom[21370] = 12'h400;
rom[21371] = 12'h400;
rom[21372] = 12'h400;
rom[21373] = 12'h400;
rom[21374] = 12'h400;
rom[21375] = 12'h400;
rom[21376] = 12'h300;
rom[21377] = 12'h300;
rom[21378] = 12'h300;
rom[21379] = 12'h200;
rom[21380] = 12'h200;
rom[21381] = 12'h200;
rom[21382] = 12'h100;
rom[21383] = 12'h100;
rom[21384] = 12'h100;
rom[21385] = 12'h100;
rom[21386] = 12'h100;
rom[21387] = 12'h  0;
rom[21388] = 12'h  0;
rom[21389] = 12'h  0;
rom[21390] = 12'h  0;
rom[21391] = 12'h  0;
rom[21392] = 12'h  0;
rom[21393] = 12'h100;
rom[21394] = 12'h111;
rom[21395] = 12'h222;
rom[21396] = 12'h333;
rom[21397] = 12'h444;
rom[21398] = 12'h544;
rom[21399] = 12'h555;
rom[21400] = 12'h555;
rom[21401] = 12'h555;
rom[21402] = 12'h777;
rom[21403] = 12'h999;
rom[21404] = 12'hbbb;
rom[21405] = 12'hbbb;
rom[21406] = 12'hbbb;
rom[21407] = 12'hbaa;
rom[21408] = 12'hbbb;
rom[21409] = 12'haaa;
rom[21410] = 12'haaa;
rom[21411] = 12'h999;
rom[21412] = 12'haaa;
rom[21413] = 12'haaa;
rom[21414] = 12'haaa;
rom[21415] = 12'haaa;
rom[21416] = 12'h999;
rom[21417] = 12'h999;
rom[21418] = 12'h999;
rom[21419] = 12'h999;
rom[21420] = 12'h999;
rom[21421] = 12'h999;
rom[21422] = 12'h999;
rom[21423] = 12'h999;
rom[21424] = 12'h999;
rom[21425] = 12'h999;
rom[21426] = 12'h888;
rom[21427] = 12'h888;
rom[21428] = 12'h888;
rom[21429] = 12'h888;
rom[21430] = 12'h888;
rom[21431] = 12'h888;
rom[21432] = 12'h777;
rom[21433] = 12'h777;
rom[21434] = 12'h777;
rom[21435] = 12'h666;
rom[21436] = 12'h666;
rom[21437] = 12'h666;
rom[21438] = 12'h666;
rom[21439] = 12'h666;
rom[21440] = 12'h555;
rom[21441] = 12'h555;
rom[21442] = 12'h444;
rom[21443] = 12'h444;
rom[21444] = 12'h444;
rom[21445] = 12'h444;
rom[21446] = 12'h444;
rom[21447] = 12'h444;
rom[21448] = 12'h333;
rom[21449] = 12'h333;
rom[21450] = 12'h222;
rom[21451] = 12'h222;
rom[21452] = 12'h222;
rom[21453] = 12'h222;
rom[21454] = 12'h111;
rom[21455] = 12'h111;
rom[21456] = 12'h111;
rom[21457] = 12'h111;
rom[21458] = 12'h  0;
rom[21459] = 12'h  0;
rom[21460] = 12'h  0;
rom[21461] = 12'h  0;
rom[21462] = 12'h111;
rom[21463] = 12'h111;
rom[21464] = 12'h111;
rom[21465] = 12'h111;
rom[21466] = 12'h111;
rom[21467] = 12'h  0;
rom[21468] = 12'h  0;
rom[21469] = 12'h  0;
rom[21470] = 12'h  0;
rom[21471] = 12'h  0;
rom[21472] = 12'h  0;
rom[21473] = 12'h  0;
rom[21474] = 12'h  0;
rom[21475] = 12'h  0;
rom[21476] = 12'h  0;
rom[21477] = 12'h  0;
rom[21478] = 12'h  0;
rom[21479] = 12'h  0;
rom[21480] = 12'h  0;
rom[21481] = 12'h  0;
rom[21482] = 12'h  0;
rom[21483] = 12'h  0;
rom[21484] = 12'h  0;
rom[21485] = 12'h  0;
rom[21486] = 12'h  0;
rom[21487] = 12'h  0;
rom[21488] = 12'h  0;
rom[21489] = 12'h  0;
rom[21490] = 12'h  0;
rom[21491] = 12'h  0;
rom[21492] = 12'h  0;
rom[21493] = 12'h  0;
rom[21494] = 12'h111;
rom[21495] = 12'h111;
rom[21496] = 12'h111;
rom[21497] = 12'h  0;
rom[21498] = 12'h111;
rom[21499] = 12'h111;
rom[21500] = 12'h111;
rom[21501] = 12'h111;
rom[21502] = 12'h222;
rom[21503] = 12'h222;
rom[21504] = 12'h222;
rom[21505] = 12'h333;
rom[21506] = 12'h333;
rom[21507] = 12'h333;
rom[21508] = 12'h222;
rom[21509] = 12'h333;
rom[21510] = 12'h333;
rom[21511] = 12'h333;
rom[21512] = 12'h333;
rom[21513] = 12'h333;
rom[21514] = 12'h333;
rom[21515] = 12'h333;
rom[21516] = 12'h333;
rom[21517] = 12'h333;
rom[21518] = 12'h333;
rom[21519] = 12'h333;
rom[21520] = 12'h333;
rom[21521] = 12'h333;
rom[21522] = 12'h333;
rom[21523] = 12'h333;
rom[21524] = 12'h333;
rom[21525] = 12'h444;
rom[21526] = 12'h444;
rom[21527] = 12'h333;
rom[21528] = 12'h333;
rom[21529] = 12'h333;
rom[21530] = 12'h333;
rom[21531] = 12'h333;
rom[21532] = 12'h333;
rom[21533] = 12'h333;
rom[21534] = 12'h333;
rom[21535] = 12'h333;
rom[21536] = 12'h333;
rom[21537] = 12'h233;
rom[21538] = 12'h333;
rom[21539] = 12'h333;
rom[21540] = 12'h344;
rom[21541] = 12'h444;
rom[21542] = 12'h555;
rom[21543] = 12'h555;
rom[21544] = 12'h666;
rom[21545] = 12'h666;
rom[21546] = 12'h666;
rom[21547] = 12'h666;
rom[21548] = 12'h665;
rom[21549] = 12'h555;
rom[21550] = 12'h555;
rom[21551] = 12'h544;
rom[21552] = 12'h555;
rom[21553] = 12'h555;
rom[21554] = 12'h555;
rom[21555] = 12'h555;
rom[21556] = 12'h555;
rom[21557] = 12'h666;
rom[21558] = 12'h666;
rom[21559] = 12'h666;
rom[21560] = 12'h666;
rom[21561] = 12'h666;
rom[21562] = 12'h666;
rom[21563] = 12'h666;
rom[21564] = 12'h666;
rom[21565] = 12'h666;
rom[21566] = 12'h666;
rom[21567] = 12'h666;
rom[21568] = 12'h666;
rom[21569] = 12'h666;
rom[21570] = 12'h666;
rom[21571] = 12'h666;
rom[21572] = 12'h666;
rom[21573] = 12'h666;
rom[21574] = 12'h666;
rom[21575] = 12'h666;
rom[21576] = 12'h777;
rom[21577] = 12'h777;
rom[21578] = 12'h666;
rom[21579] = 12'h666;
rom[21580] = 12'h666;
rom[21581] = 12'h666;
rom[21582] = 12'h666;
rom[21583] = 12'h666;
rom[21584] = 12'h777;
rom[21585] = 12'h777;
rom[21586] = 12'h777;
rom[21587] = 12'h777;
rom[21588] = 12'h777;
rom[21589] = 12'h777;
rom[21590] = 12'h888;
rom[21591] = 12'h888;
rom[21592] = 12'h888;
rom[21593] = 12'h888;
rom[21594] = 12'h999;
rom[21595] = 12'h999;
rom[21596] = 12'haaa;
rom[21597] = 12'haaa;
rom[21598] = 12'haaa;
rom[21599] = 12'haaa;
rom[21600] = 12'h555;
rom[21601] = 12'h555;
rom[21602] = 12'h555;
rom[21603] = 12'h666;
rom[21604] = 12'h666;
rom[21605] = 12'h666;
rom[21606] = 12'h666;
rom[21607] = 12'h777;
rom[21608] = 12'h777;
rom[21609] = 12'h777;
rom[21610] = 12'h777;
rom[21611] = 12'h777;
rom[21612] = 12'h777;
rom[21613] = 12'h777;
rom[21614] = 12'h666;
rom[21615] = 12'h666;
rom[21616] = 12'h666;
rom[21617] = 12'h666;
rom[21618] = 12'h666;
rom[21619] = 12'h666;
rom[21620] = 12'h666;
rom[21621] = 12'h666;
rom[21622] = 12'h666;
rom[21623] = 12'h666;
rom[21624] = 12'h666;
rom[21625] = 12'h666;
rom[21626] = 12'h666;
rom[21627] = 12'h666;
rom[21628] = 12'h666;
rom[21629] = 12'h666;
rom[21630] = 12'h666;
rom[21631] = 12'h666;
rom[21632] = 12'h666;
rom[21633] = 12'h666;
rom[21634] = 12'h777;
rom[21635] = 12'h777;
rom[21636] = 12'h777;
rom[21637] = 12'h777;
rom[21638] = 12'h777;
rom[21639] = 12'h777;
rom[21640] = 12'h777;
rom[21641] = 12'h777;
rom[21642] = 12'h777;
rom[21643] = 12'h777;
rom[21644] = 12'h777;
rom[21645] = 12'h777;
rom[21646] = 12'h777;
rom[21647] = 12'h777;
rom[21648] = 12'h777;
rom[21649] = 12'h777;
rom[21650] = 12'h666;
rom[21651] = 12'h666;
rom[21652] = 12'h666;
rom[21653] = 12'h666;
rom[21654] = 12'h666;
rom[21655] = 12'h666;
rom[21656] = 12'h666;
rom[21657] = 12'h666;
rom[21658] = 12'h666;
rom[21659] = 12'h666;
rom[21660] = 12'h666;
rom[21661] = 12'h666;
rom[21662] = 12'h666;
rom[21663] = 12'h555;
rom[21664] = 12'h555;
rom[21665] = 12'h555;
rom[21666] = 12'h555;
rom[21667] = 12'h555;
rom[21668] = 12'h666;
rom[21669] = 12'h666;
rom[21670] = 12'h666;
rom[21671] = 12'h666;
rom[21672] = 12'h666;
rom[21673] = 12'h666;
rom[21674] = 12'h666;
rom[21675] = 12'h555;
rom[21676] = 12'h555;
rom[21677] = 12'h555;
rom[21678] = 12'h555;
rom[21679] = 12'h666;
rom[21680] = 12'h666;
rom[21681] = 12'h666;
rom[21682] = 12'h666;
rom[21683] = 12'h777;
rom[21684] = 12'h777;
rom[21685] = 12'h777;
rom[21686] = 12'h666;
rom[21687] = 12'h666;
rom[21688] = 12'h444;
rom[21689] = 12'h444;
rom[21690] = 12'h444;
rom[21691] = 12'h333;
rom[21692] = 12'h222;
rom[21693] = 12'h111;
rom[21694] = 12'h111;
rom[21695] = 12'h111;
rom[21696] = 12'h  0;
rom[21697] = 12'h  0;
rom[21698] = 12'h  0;
rom[21699] = 12'h  0;
rom[21700] = 12'h  0;
rom[21701] = 12'h  0;
rom[21702] = 12'h  0;
rom[21703] = 12'h  0;
rom[21704] = 12'h  0;
rom[21705] = 12'h  0;
rom[21706] = 12'h  0;
rom[21707] = 12'h  0;
rom[21708] = 12'h  0;
rom[21709] = 12'h  0;
rom[21710] = 12'h  0;
rom[21711] = 12'h  0;
rom[21712] = 12'h100;
rom[21713] = 12'h100;
rom[21714] = 12'h100;
rom[21715] = 12'h200;
rom[21716] = 12'h200;
rom[21717] = 12'h300;
rom[21718] = 12'h410;
rom[21719] = 12'h510;
rom[21720] = 12'h620;
rom[21721] = 12'h720;
rom[21722] = 12'h930;
rom[21723] = 12'hb40;
rom[21724] = 12'hc51;
rom[21725] = 12'hd61;
rom[21726] = 12'hd61;
rom[21727] = 12'he61;
rom[21728] = 12'he50;
rom[21729] = 12'he50;
rom[21730] = 12'hd50;
rom[21731] = 12'hd40;
rom[21732] = 12'hc40;
rom[21733] = 12'hb30;
rom[21734] = 12'ha30;
rom[21735] = 12'h920;
rom[21736] = 12'h820;
rom[21737] = 12'h710;
rom[21738] = 12'h510;
rom[21739] = 12'h400;
rom[21740] = 12'h300;
rom[21741] = 12'h200;
rom[21742] = 12'h200;
rom[21743] = 12'h100;
rom[21744] = 12'h  0;
rom[21745] = 12'h  0;
rom[21746] = 12'h  0;
rom[21747] = 12'h  0;
rom[21748] = 12'h  0;
rom[21749] = 12'h  0;
rom[21750] = 12'h  0;
rom[21751] = 12'h  0;
rom[21752] = 12'h  0;
rom[21753] = 12'h  0;
rom[21754] = 12'h  0;
rom[21755] = 12'h  0;
rom[21756] = 12'h  0;
rom[21757] = 12'h  0;
rom[21758] = 12'h  0;
rom[21759] = 12'h  0;
rom[21760] = 12'h100;
rom[21761] = 12'h100;
rom[21762] = 12'h200;
rom[21763] = 12'h200;
rom[21764] = 12'h300;
rom[21765] = 12'h300;
rom[21766] = 12'h400;
rom[21767] = 12'h400;
rom[21768] = 12'h400;
rom[21769] = 12'h500;
rom[21770] = 12'h500;
rom[21771] = 12'h500;
rom[21772] = 12'h500;
rom[21773] = 12'h500;
rom[21774] = 12'h400;
rom[21775] = 12'h400;
rom[21776] = 12'h300;
rom[21777] = 12'h300;
rom[21778] = 12'h300;
rom[21779] = 12'h200;
rom[21780] = 12'h200;
rom[21781] = 12'h200;
rom[21782] = 12'h100;
rom[21783] = 12'h100;
rom[21784] = 12'h100;
rom[21785] = 12'h100;
rom[21786] = 12'h100;
rom[21787] = 12'h  0;
rom[21788] = 12'h  0;
rom[21789] = 12'h  0;
rom[21790] = 12'h  0;
rom[21791] = 12'h  0;
rom[21792] = 12'h  0;
rom[21793] = 12'h100;
rom[21794] = 12'h211;
rom[21795] = 12'h322;
rom[21796] = 12'h433;
rom[21797] = 12'h444;
rom[21798] = 12'h444;
rom[21799] = 12'h444;
rom[21800] = 12'h544;
rom[21801] = 12'h545;
rom[21802] = 12'h666;
rom[21803] = 12'h988;
rom[21804] = 12'hbaa;
rom[21805] = 12'hbbb;
rom[21806] = 12'hbbb;
rom[21807] = 12'haaa;
rom[21808] = 12'haaa;
rom[21809] = 12'haaa;
rom[21810] = 12'haaa;
rom[21811] = 12'h999;
rom[21812] = 12'h999;
rom[21813] = 12'h999;
rom[21814] = 12'h999;
rom[21815] = 12'haaa;
rom[21816] = 12'h999;
rom[21817] = 12'h999;
rom[21818] = 12'h999;
rom[21819] = 12'h999;
rom[21820] = 12'h999;
rom[21821] = 12'h999;
rom[21822] = 12'h999;
rom[21823] = 12'h999;
rom[21824] = 12'h999;
rom[21825] = 12'h888;
rom[21826] = 12'h888;
rom[21827] = 12'h888;
rom[21828] = 12'h888;
rom[21829] = 12'h888;
rom[21830] = 12'h888;
rom[21831] = 12'h777;
rom[21832] = 12'h777;
rom[21833] = 12'h777;
rom[21834] = 12'h666;
rom[21835] = 12'h666;
rom[21836] = 12'h666;
rom[21837] = 12'h666;
rom[21838] = 12'h555;
rom[21839] = 12'h555;
rom[21840] = 12'h555;
rom[21841] = 12'h555;
rom[21842] = 12'h555;
rom[21843] = 12'h555;
rom[21844] = 12'h555;
rom[21845] = 12'h444;
rom[21846] = 12'h444;
rom[21847] = 12'h444;
rom[21848] = 12'h333;
rom[21849] = 12'h222;
rom[21850] = 12'h222;
rom[21851] = 12'h222;
rom[21852] = 12'h111;
rom[21853] = 12'h111;
rom[21854] = 12'h111;
rom[21855] = 12'h111;
rom[21856] = 12'h111;
rom[21857] = 12'h111;
rom[21858] = 12'h  0;
rom[21859] = 12'h  0;
rom[21860] = 12'h  0;
rom[21861] = 12'h111;
rom[21862] = 12'h111;
rom[21863] = 12'h111;
rom[21864] = 12'h111;
rom[21865] = 12'h111;
rom[21866] = 12'h  0;
rom[21867] = 12'h  0;
rom[21868] = 12'h  0;
rom[21869] = 12'h  0;
rom[21870] = 12'h  0;
rom[21871] = 12'h  0;
rom[21872] = 12'h  0;
rom[21873] = 12'h  0;
rom[21874] = 12'h  0;
rom[21875] = 12'h  0;
rom[21876] = 12'h  0;
rom[21877] = 12'h  0;
rom[21878] = 12'h  0;
rom[21879] = 12'h  0;
rom[21880] = 12'h  0;
rom[21881] = 12'h  0;
rom[21882] = 12'h  0;
rom[21883] = 12'h  0;
rom[21884] = 12'h  0;
rom[21885] = 12'h  0;
rom[21886] = 12'h  0;
rom[21887] = 12'h  0;
rom[21888] = 12'h  0;
rom[21889] = 12'h  0;
rom[21890] = 12'h  0;
rom[21891] = 12'h  0;
rom[21892] = 12'h  0;
rom[21893] = 12'h  0;
rom[21894] = 12'h111;
rom[21895] = 12'h111;
rom[21896] = 12'h111;
rom[21897] = 12'h  0;
rom[21898] = 12'h111;
rom[21899] = 12'h111;
rom[21900] = 12'h111;
rom[21901] = 12'h111;
rom[21902] = 12'h222;
rom[21903] = 12'h222;
rom[21904] = 12'h222;
rom[21905] = 12'h333;
rom[21906] = 12'h333;
rom[21907] = 12'h333;
rom[21908] = 12'h333;
rom[21909] = 12'h333;
rom[21910] = 12'h333;
rom[21911] = 12'h333;
rom[21912] = 12'h333;
rom[21913] = 12'h333;
rom[21914] = 12'h333;
rom[21915] = 12'h333;
rom[21916] = 12'h333;
rom[21917] = 12'h333;
rom[21918] = 12'h333;
rom[21919] = 12'h333;
rom[21920] = 12'h333;
rom[21921] = 12'h333;
rom[21922] = 12'h333;
rom[21923] = 12'h333;
rom[21924] = 12'h444;
rom[21925] = 12'h444;
rom[21926] = 12'h444;
rom[21927] = 12'h444;
rom[21928] = 12'h333;
rom[21929] = 12'h333;
rom[21930] = 12'h333;
rom[21931] = 12'h333;
rom[21932] = 12'h333;
rom[21933] = 12'h333;
rom[21934] = 12'h333;
rom[21935] = 12'h333;
rom[21936] = 12'h333;
rom[21937] = 12'h333;
rom[21938] = 12'h333;
rom[21939] = 12'h444;
rom[21940] = 12'h555;
rom[21941] = 12'h555;
rom[21942] = 12'h666;
rom[21943] = 12'h666;
rom[21944] = 12'h666;
rom[21945] = 12'h666;
rom[21946] = 12'h666;
rom[21947] = 12'h666;
rom[21948] = 12'h655;
rom[21949] = 12'h655;
rom[21950] = 12'h655;
rom[21951] = 12'h655;
rom[21952] = 12'h655;
rom[21953] = 12'h665;
rom[21954] = 12'h666;
rom[21955] = 12'h666;
rom[21956] = 12'h666;
rom[21957] = 12'h666;
rom[21958] = 12'h666;
rom[21959] = 12'h666;
rom[21960] = 12'h666;
rom[21961] = 12'h666;
rom[21962] = 12'h666;
rom[21963] = 12'h666;
rom[21964] = 12'h666;
rom[21965] = 12'h666;
rom[21966] = 12'h666;
rom[21967] = 12'h666;
rom[21968] = 12'h666;
rom[21969] = 12'h666;
rom[21970] = 12'h666;
rom[21971] = 12'h666;
rom[21972] = 12'h666;
rom[21973] = 12'h666;
rom[21974] = 12'h666;
rom[21975] = 12'h666;
rom[21976] = 12'h777;
rom[21977] = 12'h777;
rom[21978] = 12'h777;
rom[21979] = 12'h777;
rom[21980] = 12'h777;
rom[21981] = 12'h777;
rom[21982] = 12'h777;
rom[21983] = 12'h777;
rom[21984] = 12'h777;
rom[21985] = 12'h777;
rom[21986] = 12'h777;
rom[21987] = 12'h777;
rom[21988] = 12'h777;
rom[21989] = 12'h777;
rom[21990] = 12'h888;
rom[21991] = 12'h888;
rom[21992] = 12'h888;
rom[21993] = 12'h888;
rom[21994] = 12'h999;
rom[21995] = 12'h999;
rom[21996] = 12'haaa;
rom[21997] = 12'haaa;
rom[21998] = 12'haaa;
rom[21999] = 12'haaa;
rom[22000] = 12'h666;
rom[22001] = 12'h666;
rom[22002] = 12'h666;
rom[22003] = 12'h666;
rom[22004] = 12'h777;
rom[22005] = 12'h777;
rom[22006] = 12'h777;
rom[22007] = 12'h777;
rom[22008] = 12'h777;
rom[22009] = 12'h777;
rom[22010] = 12'h777;
rom[22011] = 12'h777;
rom[22012] = 12'h777;
rom[22013] = 12'h666;
rom[22014] = 12'h666;
rom[22015] = 12'h666;
rom[22016] = 12'h666;
rom[22017] = 12'h666;
rom[22018] = 12'h666;
rom[22019] = 12'h666;
rom[22020] = 12'h666;
rom[22021] = 12'h666;
rom[22022] = 12'h666;
rom[22023] = 12'h666;
rom[22024] = 12'h666;
rom[22025] = 12'h666;
rom[22026] = 12'h666;
rom[22027] = 12'h666;
rom[22028] = 12'h666;
rom[22029] = 12'h666;
rom[22030] = 12'h666;
rom[22031] = 12'h666;
rom[22032] = 12'h666;
rom[22033] = 12'h666;
rom[22034] = 12'h666;
rom[22035] = 12'h777;
rom[22036] = 12'h777;
rom[22037] = 12'h777;
rom[22038] = 12'h777;
rom[22039] = 12'h777;
rom[22040] = 12'h777;
rom[22041] = 12'h777;
rom[22042] = 12'h777;
rom[22043] = 12'h777;
rom[22044] = 12'h777;
rom[22045] = 12'h777;
rom[22046] = 12'h777;
rom[22047] = 12'h777;
rom[22048] = 12'h777;
rom[22049] = 12'h777;
rom[22050] = 12'h777;
rom[22051] = 12'h777;
rom[22052] = 12'h666;
rom[22053] = 12'h666;
rom[22054] = 12'h666;
rom[22055] = 12'h666;
rom[22056] = 12'h555;
rom[22057] = 12'h666;
rom[22058] = 12'h666;
rom[22059] = 12'h666;
rom[22060] = 12'h666;
rom[22061] = 12'h666;
rom[22062] = 12'h666;
rom[22063] = 12'h666;
rom[22064] = 12'h555;
rom[22065] = 12'h555;
rom[22066] = 12'h555;
rom[22067] = 12'h555;
rom[22068] = 12'h666;
rom[22069] = 12'h666;
rom[22070] = 12'h666;
rom[22071] = 12'h666;
rom[22072] = 12'h666;
rom[22073] = 12'h666;
rom[22074] = 12'h666;
rom[22075] = 12'h555;
rom[22076] = 12'h555;
rom[22077] = 12'h555;
rom[22078] = 12'h555;
rom[22079] = 12'h555;
rom[22080] = 12'h666;
rom[22081] = 12'h666;
rom[22082] = 12'h666;
rom[22083] = 12'h777;
rom[22084] = 12'h777;
rom[22085] = 12'h777;
rom[22086] = 12'h777;
rom[22087] = 12'h666;
rom[22088] = 12'h555;
rom[22089] = 12'h444;
rom[22090] = 12'h444;
rom[22091] = 12'h333;
rom[22092] = 12'h222;
rom[22093] = 12'h222;
rom[22094] = 12'h111;
rom[22095] = 12'h111;
rom[22096] = 12'h  0;
rom[22097] = 12'h  0;
rom[22098] = 12'h  0;
rom[22099] = 12'h  0;
rom[22100] = 12'h  0;
rom[22101] = 12'h  0;
rom[22102] = 12'h  0;
rom[22103] = 12'h  0;
rom[22104] = 12'h  0;
rom[22105] = 12'h  0;
rom[22106] = 12'h  0;
rom[22107] = 12'h  0;
rom[22108] = 12'h  0;
rom[22109] = 12'h  0;
rom[22110] = 12'h  0;
rom[22111] = 12'h  0;
rom[22112] = 12'h100;
rom[22113] = 12'h100;
rom[22114] = 12'h100;
rom[22115] = 12'h200;
rom[22116] = 12'h200;
rom[22117] = 12'h300;
rom[22118] = 12'h410;
rom[22119] = 12'h510;
rom[22120] = 12'h610;
rom[22121] = 12'h720;
rom[22122] = 12'h830;
rom[22123] = 12'ha40;
rom[22124] = 12'hc51;
rom[22125] = 12'hd61;
rom[22126] = 12'hd61;
rom[22127] = 12'he61;
rom[22128] = 12'he60;
rom[22129] = 12'hf60;
rom[22130] = 12'he50;
rom[22131] = 12'hd50;
rom[22132] = 12'hc40;
rom[22133] = 12'hc30;
rom[22134] = 12'hb30;
rom[22135] = 12'ha30;
rom[22136] = 12'h820;
rom[22137] = 12'h710;
rom[22138] = 12'h610;
rom[22139] = 12'h400;
rom[22140] = 12'h300;
rom[22141] = 12'h300;
rom[22142] = 12'h200;
rom[22143] = 12'h100;
rom[22144] = 12'h100;
rom[22145] = 12'h  0;
rom[22146] = 12'h  0;
rom[22147] = 12'h  0;
rom[22148] = 12'h  0;
rom[22149] = 12'h  0;
rom[22150] = 12'h  0;
rom[22151] = 12'h  0;
rom[22152] = 12'h  0;
rom[22153] = 12'h  0;
rom[22154] = 12'h  0;
rom[22155] = 12'h  0;
rom[22156] = 12'h  0;
rom[22157] = 12'h  0;
rom[22158] = 12'h  0;
rom[22159] = 12'h100;
rom[22160] = 12'h100;
rom[22161] = 12'h200;
rom[22162] = 12'h200;
rom[22163] = 12'h300;
rom[22164] = 12'h300;
rom[22165] = 12'h400;
rom[22166] = 12'h400;
rom[22167] = 12'h400;
rom[22168] = 12'h500;
rom[22169] = 12'h500;
rom[22170] = 12'h500;
rom[22171] = 12'h500;
rom[22172] = 12'h500;
rom[22173] = 12'h500;
rom[22174] = 12'h500;
rom[22175] = 12'h400;
rom[22176] = 12'h300;
rom[22177] = 12'h300;
rom[22178] = 12'h300;
rom[22179] = 12'h200;
rom[22180] = 12'h200;
rom[22181] = 12'h200;
rom[22182] = 12'h100;
rom[22183] = 12'h100;
rom[22184] = 12'h100;
rom[22185] = 12'h100;
rom[22186] = 12'h100;
rom[22187] = 12'h  0;
rom[22188] = 12'h  0;
rom[22189] = 12'h  0;
rom[22190] = 12'h  0;
rom[22191] = 12'h  0;
rom[22192] = 12'h  0;
rom[22193] = 12'h111;
rom[22194] = 12'h222;
rom[22195] = 12'h333;
rom[22196] = 12'h444;
rom[22197] = 12'h444;
rom[22198] = 12'h444;
rom[22199] = 12'h433;
rom[22200] = 12'h444;
rom[22201] = 12'h444;
rom[22202] = 12'h655;
rom[22203] = 12'h888;
rom[22204] = 12'haaa;
rom[22205] = 12'hbbb;
rom[22206] = 12'hbaa;
rom[22207] = 12'haaa;
rom[22208] = 12'haaa;
rom[22209] = 12'haaa;
rom[22210] = 12'haaa;
rom[22211] = 12'h999;
rom[22212] = 12'h999;
rom[22213] = 12'h999;
rom[22214] = 12'h999;
rom[22215] = 12'haaa;
rom[22216] = 12'haaa;
rom[22217] = 12'h999;
rom[22218] = 12'h999;
rom[22219] = 12'h999;
rom[22220] = 12'h999;
rom[22221] = 12'h999;
rom[22222] = 12'h999;
rom[22223] = 12'h999;
rom[22224] = 12'h888;
rom[22225] = 12'h888;
rom[22226] = 12'h888;
rom[22227] = 12'h888;
rom[22228] = 12'h888;
rom[22229] = 12'h888;
rom[22230] = 12'h777;
rom[22231] = 12'h777;
rom[22232] = 12'h777;
rom[22233] = 12'h666;
rom[22234] = 12'h666;
rom[22235] = 12'h666;
rom[22236] = 12'h666;
rom[22237] = 12'h666;
rom[22238] = 12'h555;
rom[22239] = 12'h555;
rom[22240] = 12'h555;
rom[22241] = 12'h555;
rom[22242] = 12'h555;
rom[22243] = 12'h555;
rom[22244] = 12'h555;
rom[22245] = 12'h444;
rom[22246] = 12'h333;
rom[22247] = 12'h333;
rom[22248] = 12'h222;
rom[22249] = 12'h222;
rom[22250] = 12'h222;
rom[22251] = 12'h111;
rom[22252] = 12'h111;
rom[22253] = 12'h111;
rom[22254] = 12'h111;
rom[22255] = 12'h111;
rom[22256] = 12'h111;
rom[22257] = 12'h  0;
rom[22258] = 12'h  0;
rom[22259] = 12'h  0;
rom[22260] = 12'h  0;
rom[22261] = 12'h111;
rom[22262] = 12'h111;
rom[22263] = 12'h111;
rom[22264] = 12'h111;
rom[22265] = 12'h  0;
rom[22266] = 12'h  0;
rom[22267] = 12'h  0;
rom[22268] = 12'h  0;
rom[22269] = 12'h  0;
rom[22270] = 12'h  0;
rom[22271] = 12'h  0;
rom[22272] = 12'h  0;
rom[22273] = 12'h  0;
rom[22274] = 12'h  0;
rom[22275] = 12'h  0;
rom[22276] = 12'h  0;
rom[22277] = 12'h  0;
rom[22278] = 12'h  0;
rom[22279] = 12'h  0;
rom[22280] = 12'h  0;
rom[22281] = 12'h  0;
rom[22282] = 12'h  0;
rom[22283] = 12'h  0;
rom[22284] = 12'h  0;
rom[22285] = 12'h  0;
rom[22286] = 12'h  0;
rom[22287] = 12'h  0;
rom[22288] = 12'h  0;
rom[22289] = 12'h  0;
rom[22290] = 12'h  0;
rom[22291] = 12'h  0;
rom[22292] = 12'h  0;
rom[22293] = 12'h  0;
rom[22294] = 12'h111;
rom[22295] = 12'h222;
rom[22296] = 12'h111;
rom[22297] = 12'h  0;
rom[22298] = 12'h111;
rom[22299] = 12'h111;
rom[22300] = 12'h111;
rom[22301] = 12'h111;
rom[22302] = 12'h222;
rom[22303] = 12'h222;
rom[22304] = 12'h222;
rom[22305] = 12'h333;
rom[22306] = 12'h333;
rom[22307] = 12'h333;
rom[22308] = 12'h333;
rom[22309] = 12'h333;
rom[22310] = 12'h333;
rom[22311] = 12'h333;
rom[22312] = 12'h333;
rom[22313] = 12'h333;
rom[22314] = 12'h333;
rom[22315] = 12'h333;
rom[22316] = 12'h333;
rom[22317] = 12'h333;
rom[22318] = 12'h333;
rom[22319] = 12'h333;
rom[22320] = 12'h333;
rom[22321] = 12'h333;
rom[22322] = 12'h333;
rom[22323] = 12'h444;
rom[22324] = 12'h444;
rom[22325] = 12'h444;
rom[22326] = 12'h444;
rom[22327] = 12'h444;
rom[22328] = 12'h333;
rom[22329] = 12'h333;
rom[22330] = 12'h333;
rom[22331] = 12'h333;
rom[22332] = 12'h333;
rom[22333] = 12'h333;
rom[22334] = 12'h333;
rom[22335] = 12'h333;
rom[22336] = 12'h444;
rom[22337] = 12'h444;
rom[22338] = 12'h444;
rom[22339] = 12'h555;
rom[22340] = 12'h665;
rom[22341] = 12'h666;
rom[22342] = 12'h776;
rom[22343] = 12'h777;
rom[22344] = 12'h666;
rom[22345] = 12'h666;
rom[22346] = 12'h666;
rom[22347] = 12'h666;
rom[22348] = 12'h665;
rom[22349] = 12'h666;
rom[22350] = 12'h766;
rom[22351] = 12'h777;
rom[22352] = 12'h776;
rom[22353] = 12'h766;
rom[22354] = 12'h766;
rom[22355] = 12'h666;
rom[22356] = 12'h666;
rom[22357] = 12'h666;
rom[22358] = 12'h666;
rom[22359] = 12'h666;
rom[22360] = 12'h666;
rom[22361] = 12'h666;
rom[22362] = 12'h666;
rom[22363] = 12'h666;
rom[22364] = 12'h666;
rom[22365] = 12'h666;
rom[22366] = 12'h666;
rom[22367] = 12'h666;
rom[22368] = 12'h666;
rom[22369] = 12'h666;
rom[22370] = 12'h666;
rom[22371] = 12'h666;
rom[22372] = 12'h666;
rom[22373] = 12'h666;
rom[22374] = 12'h666;
rom[22375] = 12'h666;
rom[22376] = 12'h666;
rom[22377] = 12'h666;
rom[22378] = 12'h777;
rom[22379] = 12'h777;
rom[22380] = 12'h777;
rom[22381] = 12'h777;
rom[22382] = 12'h777;
rom[22383] = 12'h777;
rom[22384] = 12'h777;
rom[22385] = 12'h777;
rom[22386] = 12'h777;
rom[22387] = 12'h777;
rom[22388] = 12'h777;
rom[22389] = 12'h888;
rom[22390] = 12'h888;
rom[22391] = 12'h888;
rom[22392] = 12'h888;
rom[22393] = 12'h888;
rom[22394] = 12'h999;
rom[22395] = 12'h999;
rom[22396] = 12'haaa;
rom[22397] = 12'haaa;
rom[22398] = 12'haaa;
rom[22399] = 12'haaa;
rom[22400] = 12'h777;
rom[22401] = 12'h777;
rom[22402] = 12'h777;
rom[22403] = 12'h777;
rom[22404] = 12'h777;
rom[22405] = 12'h777;
rom[22406] = 12'h777;
rom[22407] = 12'h777;
rom[22408] = 12'h777;
rom[22409] = 12'h777;
rom[22410] = 12'h777;
rom[22411] = 12'h666;
rom[22412] = 12'h666;
rom[22413] = 12'h666;
rom[22414] = 12'h666;
rom[22415] = 12'h666;
rom[22416] = 12'h666;
rom[22417] = 12'h666;
rom[22418] = 12'h666;
rom[22419] = 12'h666;
rom[22420] = 12'h555;
rom[22421] = 12'h555;
rom[22422] = 12'h555;
rom[22423] = 12'h555;
rom[22424] = 12'h555;
rom[22425] = 12'h555;
rom[22426] = 12'h555;
rom[22427] = 12'h555;
rom[22428] = 12'h666;
rom[22429] = 12'h666;
rom[22430] = 12'h666;
rom[22431] = 12'h666;
rom[22432] = 12'h666;
rom[22433] = 12'h666;
rom[22434] = 12'h666;
rom[22435] = 12'h666;
rom[22436] = 12'h777;
rom[22437] = 12'h777;
rom[22438] = 12'h777;
rom[22439] = 12'h777;
rom[22440] = 12'h777;
rom[22441] = 12'h777;
rom[22442] = 12'h777;
rom[22443] = 12'h777;
rom[22444] = 12'h777;
rom[22445] = 12'h777;
rom[22446] = 12'h777;
rom[22447] = 12'h777;
rom[22448] = 12'h777;
rom[22449] = 12'h777;
rom[22450] = 12'h777;
rom[22451] = 12'h666;
rom[22452] = 12'h666;
rom[22453] = 12'h666;
rom[22454] = 12'h666;
rom[22455] = 12'h666;
rom[22456] = 12'h555;
rom[22457] = 12'h555;
rom[22458] = 12'h555;
rom[22459] = 12'h666;
rom[22460] = 12'h666;
rom[22461] = 12'h666;
rom[22462] = 12'h666;
rom[22463] = 12'h666;
rom[22464] = 12'h666;
rom[22465] = 12'h666;
rom[22466] = 12'h666;
rom[22467] = 12'h666;
rom[22468] = 12'h666;
rom[22469] = 12'h666;
rom[22470] = 12'h666;
rom[22471] = 12'h666;
rom[22472] = 12'h555;
rom[22473] = 12'h555;
rom[22474] = 12'h555;
rom[22475] = 12'h555;
rom[22476] = 12'h555;
rom[22477] = 12'h555;
rom[22478] = 12'h555;
rom[22479] = 12'h555;
rom[22480] = 12'h666;
rom[22481] = 12'h666;
rom[22482] = 12'h666;
rom[22483] = 12'h666;
rom[22484] = 12'h666;
rom[22485] = 12'h666;
rom[22486] = 12'h666;
rom[22487] = 12'h777;
rom[22488] = 12'h555;
rom[22489] = 12'h555;
rom[22490] = 12'h444;
rom[22491] = 12'h333;
rom[22492] = 12'h333;
rom[22493] = 12'h222;
rom[22494] = 12'h222;
rom[22495] = 12'h111;
rom[22496] = 12'h  0;
rom[22497] = 12'h  0;
rom[22498] = 12'h  0;
rom[22499] = 12'h  0;
rom[22500] = 12'h  0;
rom[22501] = 12'h  0;
rom[22502] = 12'h  0;
rom[22503] = 12'h  0;
rom[22504] = 12'h  0;
rom[22505] = 12'h  0;
rom[22506] = 12'h  0;
rom[22507] = 12'h  0;
rom[22508] = 12'h  0;
rom[22509] = 12'h  0;
rom[22510] = 12'h  0;
rom[22511] = 12'h  0;
rom[22512] = 12'h100;
rom[22513] = 12'h100;
rom[22514] = 12'h200;
rom[22515] = 12'h200;
rom[22516] = 12'h200;
rom[22517] = 12'h300;
rom[22518] = 12'h410;
rom[22519] = 12'h410;
rom[22520] = 12'h620;
rom[22521] = 12'h720;
rom[22522] = 12'h830;
rom[22523] = 12'h940;
rom[22524] = 12'hb50;
rom[22525] = 12'hc61;
rom[22526] = 12'hd61;
rom[22527] = 12'he71;
rom[22528] = 12'hf71;
rom[22529] = 12'hf61;
rom[22530] = 12'hf60;
rom[22531] = 12'he50;
rom[22532] = 12'he50;
rom[22533] = 12'hd40;
rom[22534] = 12'hc40;
rom[22535] = 12'hb30;
rom[22536] = 12'ha30;
rom[22537] = 12'h820;
rom[22538] = 12'h710;
rom[22539] = 12'h510;
rom[22540] = 12'h400;
rom[22541] = 12'h300;
rom[22542] = 12'h300;
rom[22543] = 12'h200;
rom[22544] = 12'h100;
rom[22545] = 12'h100;
rom[22546] = 12'h  0;
rom[22547] = 12'h  0;
rom[22548] = 12'h  0;
rom[22549] = 12'h  0;
rom[22550] = 12'h  0;
rom[22551] = 12'h  0;
rom[22552] = 12'h  0;
rom[22553] = 12'h  0;
rom[22554] = 12'h  0;
rom[22555] = 12'h  0;
rom[22556] = 12'h100;
rom[22557] = 12'h100;
rom[22558] = 12'h100;
rom[22559] = 12'h200;
rom[22560] = 12'h200;
rom[22561] = 12'h300;
rom[22562] = 12'h300;
rom[22563] = 12'h300;
rom[22564] = 12'h400;
rom[22565] = 12'h400;
rom[22566] = 12'h500;
rom[22567] = 12'h500;
rom[22568] = 12'h500;
rom[22569] = 12'h500;
rom[22570] = 12'h600;
rom[22571] = 12'h600;
rom[22572] = 12'h500;
rom[22573] = 12'h500;
rom[22574] = 12'h500;
rom[22575] = 12'h400;
rom[22576] = 12'h300;
rom[22577] = 12'h300;
rom[22578] = 12'h300;
rom[22579] = 12'h200;
rom[22580] = 12'h200;
rom[22581] = 12'h200;
rom[22582] = 12'h100;
rom[22583] = 12'h100;
rom[22584] = 12'h100;
rom[22585] = 12'h100;
rom[22586] = 12'h100;
rom[22587] = 12'h100;
rom[22588] = 12'h  0;
rom[22589] = 12'h  0;
rom[22590] = 12'h  0;
rom[22591] = 12'h  0;
rom[22592] = 12'h  0;
rom[22593] = 12'h111;
rom[22594] = 12'h322;
rom[22595] = 12'h433;
rom[22596] = 12'h444;
rom[22597] = 12'h444;
rom[22598] = 12'h444;
rom[22599] = 12'h433;
rom[22600] = 12'h444;
rom[22601] = 12'h444;
rom[22602] = 12'h555;
rom[22603] = 12'h777;
rom[22604] = 12'h999;
rom[22605] = 12'hbaa;
rom[22606] = 12'haaa;
rom[22607] = 12'haaa;
rom[22608] = 12'haaa;
rom[22609] = 12'haaa;
rom[22610] = 12'haaa;
rom[22611] = 12'h999;
rom[22612] = 12'h999;
rom[22613] = 12'h999;
rom[22614] = 12'h999;
rom[22615] = 12'h999;
rom[22616] = 12'h999;
rom[22617] = 12'h999;
rom[22618] = 12'h999;
rom[22619] = 12'h999;
rom[22620] = 12'h999;
rom[22621] = 12'h999;
rom[22622] = 12'h999;
rom[22623] = 12'h888;
rom[22624] = 12'h888;
rom[22625] = 12'h888;
rom[22626] = 12'h888;
rom[22627] = 12'h888;
rom[22628] = 12'h888;
rom[22629] = 12'h777;
rom[22630] = 12'h777;
rom[22631] = 12'h777;
rom[22632] = 12'h666;
rom[22633] = 12'h666;
rom[22634] = 12'h666;
rom[22635] = 12'h666;
rom[22636] = 12'h666;
rom[22637] = 12'h666;
rom[22638] = 12'h666;
rom[22639] = 12'h666;
rom[22640] = 12'h666;
rom[22641] = 12'h555;
rom[22642] = 12'h555;
rom[22643] = 12'h444;
rom[22644] = 12'h444;
rom[22645] = 12'h444;
rom[22646] = 12'h333;
rom[22647] = 12'h333;
rom[22648] = 12'h222;
rom[22649] = 12'h222;
rom[22650] = 12'h111;
rom[22651] = 12'h111;
rom[22652] = 12'h111;
rom[22653] = 12'h111;
rom[22654] = 12'h111;
rom[22655] = 12'h  0;
rom[22656] = 12'h  0;
rom[22657] = 12'h  0;
rom[22658] = 12'h111;
rom[22659] = 12'h111;
rom[22660] = 12'h111;
rom[22661] = 12'h111;
rom[22662] = 12'h111;
rom[22663] = 12'h111;
rom[22664] = 12'h  0;
rom[22665] = 12'h  0;
rom[22666] = 12'h  0;
rom[22667] = 12'h  0;
rom[22668] = 12'h  0;
rom[22669] = 12'h  0;
rom[22670] = 12'h  0;
rom[22671] = 12'h  0;
rom[22672] = 12'h  0;
rom[22673] = 12'h  0;
rom[22674] = 12'h  0;
rom[22675] = 12'h  0;
rom[22676] = 12'h  0;
rom[22677] = 12'h  0;
rom[22678] = 12'h  0;
rom[22679] = 12'h  0;
rom[22680] = 12'h  0;
rom[22681] = 12'h  0;
rom[22682] = 12'h  0;
rom[22683] = 12'h  0;
rom[22684] = 12'h  0;
rom[22685] = 12'h  0;
rom[22686] = 12'h  0;
rom[22687] = 12'h  0;
rom[22688] = 12'h  0;
rom[22689] = 12'h  0;
rom[22690] = 12'h  0;
rom[22691] = 12'h  0;
rom[22692] = 12'h  0;
rom[22693] = 12'h111;
rom[22694] = 12'h111;
rom[22695] = 12'h111;
rom[22696] = 12'h111;
rom[22697] = 12'h111;
rom[22698] = 12'h111;
rom[22699] = 12'h111;
rom[22700] = 12'h111;
rom[22701] = 12'h111;
rom[22702] = 12'h222;
rom[22703] = 12'h333;
rom[22704] = 12'h222;
rom[22705] = 12'h222;
rom[22706] = 12'h333;
rom[22707] = 12'h333;
rom[22708] = 12'h333;
rom[22709] = 12'h333;
rom[22710] = 12'h333;
rom[22711] = 12'h333;
rom[22712] = 12'h333;
rom[22713] = 12'h333;
rom[22714] = 12'h333;
rom[22715] = 12'h333;
rom[22716] = 12'h333;
rom[22717] = 12'h333;
rom[22718] = 12'h333;
rom[22719] = 12'h333;
rom[22720] = 12'h333;
rom[22721] = 12'h333;
rom[22722] = 12'h333;
rom[22723] = 12'h444;
rom[22724] = 12'h444;
rom[22725] = 12'h444;
rom[22726] = 12'h444;
rom[22727] = 12'h444;
rom[22728] = 12'h333;
rom[22729] = 12'h333;
rom[22730] = 12'h333;
rom[22731] = 12'h333;
rom[22732] = 12'h333;
rom[22733] = 12'h333;
rom[22734] = 12'h444;
rom[22735] = 12'h444;
rom[22736] = 12'h444;
rom[22737] = 12'h555;
rom[22738] = 12'h665;
rom[22739] = 12'h666;
rom[22740] = 12'h777;
rom[22741] = 12'h777;
rom[22742] = 12'h776;
rom[22743] = 12'h766;
rom[22744] = 12'h766;
rom[22745] = 12'h666;
rom[22746] = 12'h666;
rom[22747] = 12'h766;
rom[22748] = 12'h777;
rom[22749] = 12'h777;
rom[22750] = 12'h877;
rom[22751] = 12'h877;
rom[22752] = 12'h777;
rom[22753] = 12'h777;
rom[22754] = 12'h777;
rom[22755] = 12'h776;
rom[22756] = 12'h766;
rom[22757] = 12'h666;
rom[22758] = 12'h666;
rom[22759] = 12'h666;
rom[22760] = 12'h666;
rom[22761] = 12'h666;
rom[22762] = 12'h666;
rom[22763] = 12'h666;
rom[22764] = 12'h666;
rom[22765] = 12'h666;
rom[22766] = 12'h666;
rom[22767] = 12'h666;
rom[22768] = 12'h666;
rom[22769] = 12'h666;
rom[22770] = 12'h666;
rom[22771] = 12'h666;
rom[22772] = 12'h666;
rom[22773] = 12'h666;
rom[22774] = 12'h666;
rom[22775] = 12'h666;
rom[22776] = 12'h666;
rom[22777] = 12'h666;
rom[22778] = 12'h666;
rom[22779] = 12'h666;
rom[22780] = 12'h777;
rom[22781] = 12'h777;
rom[22782] = 12'h777;
rom[22783] = 12'h777;
rom[22784] = 12'h777;
rom[22785] = 12'h777;
rom[22786] = 12'h777;
rom[22787] = 12'h777;
rom[22788] = 12'h888;
rom[22789] = 12'h888;
rom[22790] = 12'h888;
rom[22791] = 12'h888;
rom[22792] = 12'h888;
rom[22793] = 12'h888;
rom[22794] = 12'h999;
rom[22795] = 12'h999;
rom[22796] = 12'haaa;
rom[22797] = 12'haaa;
rom[22798] = 12'haaa;
rom[22799] = 12'haaa;
rom[22800] = 12'h777;
rom[22801] = 12'h777;
rom[22802] = 12'h777;
rom[22803] = 12'h777;
rom[22804] = 12'h777;
rom[22805] = 12'h777;
rom[22806] = 12'h777;
rom[22807] = 12'h777;
rom[22808] = 12'h666;
rom[22809] = 12'h666;
rom[22810] = 12'h666;
rom[22811] = 12'h666;
rom[22812] = 12'h666;
rom[22813] = 12'h666;
rom[22814] = 12'h666;
rom[22815] = 12'h666;
rom[22816] = 12'h666;
rom[22817] = 12'h666;
rom[22818] = 12'h666;
rom[22819] = 12'h666;
rom[22820] = 12'h666;
rom[22821] = 12'h666;
rom[22822] = 12'h666;
rom[22823] = 12'h666;
rom[22824] = 12'h555;
rom[22825] = 12'h666;
rom[22826] = 12'h666;
rom[22827] = 12'h666;
rom[22828] = 12'h666;
rom[22829] = 12'h666;
rom[22830] = 12'h666;
rom[22831] = 12'h666;
rom[22832] = 12'h666;
rom[22833] = 12'h666;
rom[22834] = 12'h666;
rom[22835] = 12'h666;
rom[22836] = 12'h777;
rom[22837] = 12'h777;
rom[22838] = 12'h777;
rom[22839] = 12'h777;
rom[22840] = 12'h777;
rom[22841] = 12'h777;
rom[22842] = 12'h777;
rom[22843] = 12'h777;
rom[22844] = 12'h777;
rom[22845] = 12'h777;
rom[22846] = 12'h777;
rom[22847] = 12'h777;
rom[22848] = 12'h777;
rom[22849] = 12'h777;
rom[22850] = 12'h777;
rom[22851] = 12'h777;
rom[22852] = 12'h666;
rom[22853] = 12'h666;
rom[22854] = 12'h666;
rom[22855] = 12'h666;
rom[22856] = 12'h555;
rom[22857] = 12'h555;
rom[22858] = 12'h555;
rom[22859] = 12'h666;
rom[22860] = 12'h666;
rom[22861] = 12'h666;
rom[22862] = 12'h666;
rom[22863] = 12'h666;
rom[22864] = 12'h666;
rom[22865] = 12'h666;
rom[22866] = 12'h666;
rom[22867] = 12'h666;
rom[22868] = 12'h666;
rom[22869] = 12'h666;
rom[22870] = 12'h666;
rom[22871] = 12'h666;
rom[22872] = 12'h555;
rom[22873] = 12'h555;
rom[22874] = 12'h555;
rom[22875] = 12'h555;
rom[22876] = 12'h555;
rom[22877] = 12'h555;
rom[22878] = 12'h555;
rom[22879] = 12'h555;
rom[22880] = 12'h555;
rom[22881] = 12'h555;
rom[22882] = 12'h555;
rom[22883] = 12'h555;
rom[22884] = 12'h555;
rom[22885] = 12'h666;
rom[22886] = 12'h666;
rom[22887] = 12'h666;
rom[22888] = 12'h666;
rom[22889] = 12'h555;
rom[22890] = 12'h444;
rom[22891] = 12'h444;
rom[22892] = 12'h333;
rom[22893] = 12'h222;
rom[22894] = 12'h222;
rom[22895] = 12'h111;
rom[22896] = 12'h100;
rom[22897] = 12'h  0;
rom[22898] = 12'h  0;
rom[22899] = 12'h  0;
rom[22900] = 12'h  0;
rom[22901] = 12'h  0;
rom[22902] = 12'h  0;
rom[22903] = 12'h  0;
rom[22904] = 12'h  0;
rom[22905] = 12'h  0;
rom[22906] = 12'h  0;
rom[22907] = 12'h  0;
rom[22908] = 12'h  0;
rom[22909] = 12'h  0;
rom[22910] = 12'h  0;
rom[22911] = 12'h  0;
rom[22912] = 12'h100;
rom[22913] = 12'h100;
rom[22914] = 12'h100;
rom[22915] = 12'h200;
rom[22916] = 12'h200;
rom[22917] = 12'h200;
rom[22918] = 12'h300;
rom[22919] = 12'h410;
rom[22920] = 12'h510;
rom[22921] = 12'h620;
rom[22922] = 12'h720;
rom[22923] = 12'h930;
rom[22924] = 12'ha40;
rom[22925] = 12'hc51;
rom[22926] = 12'hd61;
rom[22927] = 12'he61;
rom[22928] = 12'hf71;
rom[22929] = 12'hf71;
rom[22930] = 12'hf60;
rom[22931] = 12'hf60;
rom[22932] = 12'hf60;
rom[22933] = 12'he60;
rom[22934] = 12'hd50;
rom[22935] = 12'hc40;
rom[22936] = 12'hb30;
rom[22937] = 12'h930;
rom[22938] = 12'h820;
rom[22939] = 12'h610;
rom[22940] = 12'h500;
rom[22941] = 12'h400;
rom[22942] = 12'h400;
rom[22943] = 12'h300;
rom[22944] = 12'h200;
rom[22945] = 12'h200;
rom[22946] = 12'h100;
rom[22947] = 12'h100;
rom[22948] = 12'h100;
rom[22949] = 12'h  0;
rom[22950] = 12'h  0;
rom[22951] = 12'h  0;
rom[22952] = 12'h  0;
rom[22953] = 12'h  0;
rom[22954] = 12'h100;
rom[22955] = 12'h100;
rom[22956] = 12'h200;
rom[22957] = 12'h200;
rom[22958] = 12'h200;
rom[22959] = 12'h300;
rom[22960] = 12'h300;
rom[22961] = 12'h400;
rom[22962] = 12'h400;
rom[22963] = 12'h400;
rom[22964] = 12'h500;
rom[22965] = 12'h500;
rom[22966] = 12'h500;
rom[22967] = 12'h600;
rom[22968] = 12'h600;
rom[22969] = 12'h600;
rom[22970] = 12'h600;
rom[22971] = 12'h600;
rom[22972] = 12'h600;
rom[22973] = 12'h500;
rom[22974] = 12'h500;
rom[22975] = 12'h400;
rom[22976] = 12'h400;
rom[22977] = 12'h300;
rom[22978] = 12'h300;
rom[22979] = 12'h200;
rom[22980] = 12'h200;
rom[22981] = 12'h200;
rom[22982] = 12'h200;
rom[22983] = 12'h100;
rom[22984] = 12'h100;
rom[22985] = 12'h100;
rom[22986] = 12'h100;
rom[22987] = 12'h100;
rom[22988] = 12'h  0;
rom[22989] = 12'h  0;
rom[22990] = 12'h  0;
rom[22991] = 12'h  0;
rom[22992] = 12'h111;
rom[22993] = 12'h111;
rom[22994] = 12'h333;
rom[22995] = 12'h333;
rom[22996] = 12'h333;
rom[22997] = 12'h333;
rom[22998] = 12'h333;
rom[22999] = 12'h433;
rom[23000] = 12'h444;
rom[23001] = 12'h444;
rom[23002] = 12'h555;
rom[23003] = 12'h777;
rom[23004] = 12'h999;
rom[23005] = 12'haaa;
rom[23006] = 12'haaa;
rom[23007] = 12'haaa;
rom[23008] = 12'haaa;
rom[23009] = 12'haaa;
rom[23010] = 12'haaa;
rom[23011] = 12'h999;
rom[23012] = 12'h999;
rom[23013] = 12'h999;
rom[23014] = 12'h999;
rom[23015] = 12'h999;
rom[23016] = 12'h999;
rom[23017] = 12'h999;
rom[23018] = 12'h999;
rom[23019] = 12'h999;
rom[23020] = 12'h999;
rom[23021] = 12'h999;
rom[23022] = 12'h999;
rom[23023] = 12'h888;
rom[23024] = 12'h888;
rom[23025] = 12'h888;
rom[23026] = 12'h888;
rom[23027] = 12'h888;
rom[23028] = 12'h888;
rom[23029] = 12'h888;
rom[23030] = 12'h777;
rom[23031] = 12'h777;
rom[23032] = 12'h777;
rom[23033] = 12'h777;
rom[23034] = 12'h666;
rom[23035] = 12'h666;
rom[23036] = 12'h666;
rom[23037] = 12'h666;
rom[23038] = 12'h666;
rom[23039] = 12'h666;
rom[23040] = 12'h555;
rom[23041] = 12'h555;
rom[23042] = 12'h444;
rom[23043] = 12'h444;
rom[23044] = 12'h333;
rom[23045] = 12'h333;
rom[23046] = 12'h333;
rom[23047] = 12'h222;
rom[23048] = 12'h222;
rom[23049] = 12'h222;
rom[23050] = 12'h111;
rom[23051] = 12'h111;
rom[23052] = 12'h111;
rom[23053] = 12'h111;
rom[23054] = 12'h111;
rom[23055] = 12'h  0;
rom[23056] = 12'h111;
rom[23057] = 12'h111;
rom[23058] = 12'h111;
rom[23059] = 12'h111;
rom[23060] = 12'h111;
rom[23061] = 12'h111;
rom[23062] = 12'h111;
rom[23063] = 12'h111;
rom[23064] = 12'h  0;
rom[23065] = 12'h  0;
rom[23066] = 12'h  0;
rom[23067] = 12'h  0;
rom[23068] = 12'h  0;
rom[23069] = 12'h  0;
rom[23070] = 12'h  0;
rom[23071] = 12'h  0;
rom[23072] = 12'h  0;
rom[23073] = 12'h  0;
rom[23074] = 12'h  0;
rom[23075] = 12'h  0;
rom[23076] = 12'h  0;
rom[23077] = 12'h  0;
rom[23078] = 12'h  0;
rom[23079] = 12'h  0;
rom[23080] = 12'h  0;
rom[23081] = 12'h  0;
rom[23082] = 12'h  0;
rom[23083] = 12'h  0;
rom[23084] = 12'h  0;
rom[23085] = 12'h  0;
rom[23086] = 12'h  0;
rom[23087] = 12'h  0;
rom[23088] = 12'h  0;
rom[23089] = 12'h  0;
rom[23090] = 12'h  0;
rom[23091] = 12'h  0;
rom[23092] = 12'h  0;
rom[23093] = 12'h111;
rom[23094] = 12'h111;
rom[23095] = 12'h111;
rom[23096] = 12'h111;
rom[23097] = 12'h111;
rom[23098] = 12'h111;
rom[23099] = 12'h111;
rom[23100] = 12'h111;
rom[23101] = 12'h111;
rom[23102] = 12'h222;
rom[23103] = 12'h333;
rom[23104] = 12'h222;
rom[23105] = 12'h222;
rom[23106] = 12'h333;
rom[23107] = 12'h333;
rom[23108] = 12'h333;
rom[23109] = 12'h333;
rom[23110] = 12'h333;
rom[23111] = 12'h333;
rom[23112] = 12'h333;
rom[23113] = 12'h333;
rom[23114] = 12'h333;
rom[23115] = 12'h333;
rom[23116] = 12'h333;
rom[23117] = 12'h333;
rom[23118] = 12'h333;
rom[23119] = 12'h444;
rom[23120] = 12'h333;
rom[23121] = 12'h333;
rom[23122] = 12'h333;
rom[23123] = 12'h444;
rom[23124] = 12'h444;
rom[23125] = 12'h444;
rom[23126] = 12'h444;
rom[23127] = 12'h444;
rom[23128] = 12'h444;
rom[23129] = 12'h444;
rom[23130] = 12'h444;
rom[23131] = 12'h333;
rom[23132] = 12'h333;
rom[23133] = 12'h333;
rom[23134] = 12'h444;
rom[23135] = 12'h555;
rom[23136] = 12'h555;
rom[23137] = 12'h666;
rom[23138] = 12'h666;
rom[23139] = 12'h777;
rom[23140] = 12'h777;
rom[23141] = 12'h777;
rom[23142] = 12'h777;
rom[23143] = 12'h777;
rom[23144] = 12'h777;
rom[23145] = 12'h777;
rom[23146] = 12'h777;
rom[23147] = 12'h777;
rom[23148] = 12'h877;
rom[23149] = 12'h877;
rom[23150] = 12'h777;
rom[23151] = 12'h777;
rom[23152] = 12'h777;
rom[23153] = 12'h776;
rom[23154] = 12'h776;
rom[23155] = 12'h766;
rom[23156] = 12'h666;
rom[23157] = 12'h666;
rom[23158] = 12'h666;
rom[23159] = 12'h666;
rom[23160] = 12'h666;
rom[23161] = 12'h666;
rom[23162] = 12'h666;
rom[23163] = 12'h666;
rom[23164] = 12'h766;
rom[23165] = 12'h766;
rom[23166] = 12'h766;
rom[23167] = 12'h666;
rom[23168] = 12'h666;
rom[23169] = 12'h666;
rom[23170] = 12'h666;
rom[23171] = 12'h666;
rom[23172] = 12'h666;
rom[23173] = 12'h666;
rom[23174] = 12'h666;
rom[23175] = 12'h666;
rom[23176] = 12'h666;
rom[23177] = 12'h666;
rom[23178] = 12'h666;
rom[23179] = 12'h666;
rom[23180] = 12'h666;
rom[23181] = 12'h666;
rom[23182] = 12'h666;
rom[23183] = 12'h666;
rom[23184] = 12'h777;
rom[23185] = 12'h777;
rom[23186] = 12'h777;
rom[23187] = 12'h777;
rom[23188] = 12'h777;
rom[23189] = 12'h888;
rom[23190] = 12'h888;
rom[23191] = 12'h888;
rom[23192] = 12'h888;
rom[23193] = 12'h888;
rom[23194] = 12'h999;
rom[23195] = 12'h999;
rom[23196] = 12'haaa;
rom[23197] = 12'haaa;
rom[23198] = 12'haaa;
rom[23199] = 12'haaa;
rom[23200] = 12'h777;
rom[23201] = 12'h777;
rom[23202] = 12'h777;
rom[23203] = 12'h777;
rom[23204] = 12'h777;
rom[23205] = 12'h777;
rom[23206] = 12'h777;
rom[23207] = 12'h777;
rom[23208] = 12'h666;
rom[23209] = 12'h666;
rom[23210] = 12'h666;
rom[23211] = 12'h666;
rom[23212] = 12'h666;
rom[23213] = 12'h666;
rom[23214] = 12'h666;
rom[23215] = 12'h666;
rom[23216] = 12'h666;
rom[23217] = 12'h666;
rom[23218] = 12'h666;
rom[23219] = 12'h666;
rom[23220] = 12'h666;
rom[23221] = 12'h666;
rom[23222] = 12'h666;
rom[23223] = 12'h666;
rom[23224] = 12'h666;
rom[23225] = 12'h666;
rom[23226] = 12'h666;
rom[23227] = 12'h666;
rom[23228] = 12'h666;
rom[23229] = 12'h666;
rom[23230] = 12'h666;
rom[23231] = 12'h666;
rom[23232] = 12'h666;
rom[23233] = 12'h666;
rom[23234] = 12'h666;
rom[23235] = 12'h666;
rom[23236] = 12'h777;
rom[23237] = 12'h777;
rom[23238] = 12'h777;
rom[23239] = 12'h777;
rom[23240] = 12'h777;
rom[23241] = 12'h777;
rom[23242] = 12'h777;
rom[23243] = 12'h777;
rom[23244] = 12'h777;
rom[23245] = 12'h777;
rom[23246] = 12'h777;
rom[23247] = 12'h777;
rom[23248] = 12'h777;
rom[23249] = 12'h777;
rom[23250] = 12'h777;
rom[23251] = 12'h777;
rom[23252] = 12'h777;
rom[23253] = 12'h666;
rom[23254] = 12'h666;
rom[23255] = 12'h666;
rom[23256] = 12'h666;
rom[23257] = 12'h666;
rom[23258] = 12'h666;
rom[23259] = 12'h666;
rom[23260] = 12'h666;
rom[23261] = 12'h666;
rom[23262] = 12'h666;
rom[23263] = 12'h666;
rom[23264] = 12'h666;
rom[23265] = 12'h666;
rom[23266] = 12'h666;
rom[23267] = 12'h666;
rom[23268] = 12'h666;
rom[23269] = 12'h666;
rom[23270] = 12'h666;
rom[23271] = 12'h666;
rom[23272] = 12'h555;
rom[23273] = 12'h555;
rom[23274] = 12'h666;
rom[23275] = 12'h666;
rom[23276] = 12'h555;
rom[23277] = 12'h555;
rom[23278] = 12'h555;
rom[23279] = 12'h555;
rom[23280] = 12'h555;
rom[23281] = 12'h555;
rom[23282] = 12'h555;
rom[23283] = 12'h555;
rom[23284] = 12'h555;
rom[23285] = 12'h555;
rom[23286] = 12'h555;
rom[23287] = 12'h555;
rom[23288] = 12'h666;
rom[23289] = 12'h555;
rom[23290] = 12'h555;
rom[23291] = 12'h444;
rom[23292] = 12'h444;
rom[23293] = 12'h333;
rom[23294] = 12'h222;
rom[23295] = 12'h111;
rom[23296] = 12'h111;
rom[23297] = 12'h100;
rom[23298] = 12'h  0;
rom[23299] = 12'h  0;
rom[23300] = 12'h  0;
rom[23301] = 12'h  0;
rom[23302] = 12'h  0;
rom[23303] = 12'h  0;
rom[23304] = 12'h  0;
rom[23305] = 12'h  0;
rom[23306] = 12'h  0;
rom[23307] = 12'h  0;
rom[23308] = 12'h  0;
rom[23309] = 12'h  0;
rom[23310] = 12'h  0;
rom[23311] = 12'h  0;
rom[23312] = 12'h100;
rom[23313] = 12'h100;
rom[23314] = 12'h100;
rom[23315] = 12'h100;
rom[23316] = 12'h200;
rom[23317] = 12'h200;
rom[23318] = 12'h300;
rom[23319] = 12'h310;
rom[23320] = 12'h410;
rom[23321] = 12'h510;
rom[23322] = 12'h620;
rom[23323] = 12'h830;
rom[23324] = 12'h940;
rom[23325] = 12'hb50;
rom[23326] = 12'hc51;
rom[23327] = 12'hd61;
rom[23328] = 12'hf71;
rom[23329] = 12'hf71;
rom[23330] = 12'hf71;
rom[23331] = 12'hf71;
rom[23332] = 12'hf71;
rom[23333] = 12'hf71;
rom[23334] = 12'he61;
rom[23335] = 12'hd61;
rom[23336] = 12'hc50;
rom[23337] = 12'ha40;
rom[23338] = 12'h930;
rom[23339] = 12'h720;
rom[23340] = 12'h610;
rom[23341] = 12'h510;
rom[23342] = 12'h510;
rom[23343] = 12'h400;
rom[23344] = 12'h300;
rom[23345] = 12'h200;
rom[23346] = 12'h200;
rom[23347] = 12'h200;
rom[23348] = 12'h100;
rom[23349] = 12'h100;
rom[23350] = 12'h100;
rom[23351] = 12'h100;
rom[23352] = 12'h100;
rom[23353] = 12'h100;
rom[23354] = 12'h200;
rom[23355] = 12'h200;
rom[23356] = 12'h300;
rom[23357] = 12'h300;
rom[23358] = 12'h300;
rom[23359] = 12'h400;
rom[23360] = 12'h400;
rom[23361] = 12'h500;
rom[23362] = 12'h500;
rom[23363] = 12'h500;
rom[23364] = 12'h600;
rom[23365] = 12'h600;
rom[23366] = 12'h610;
rom[23367] = 12'h610;
rom[23368] = 12'h610;
rom[23369] = 12'h610;
rom[23370] = 12'h600;
rom[23371] = 12'h600;
rom[23372] = 12'h600;
rom[23373] = 12'h500;
rom[23374] = 12'h500;
rom[23375] = 12'h400;
rom[23376] = 12'h300;
rom[23377] = 12'h300;
rom[23378] = 12'h300;
rom[23379] = 12'h200;
rom[23380] = 12'h200;
rom[23381] = 12'h200;
rom[23382] = 12'h200;
rom[23383] = 12'h100;
rom[23384] = 12'h100;
rom[23385] = 12'h100;
rom[23386] = 12'h100;
rom[23387] = 12'h  0;
rom[23388] = 12'h  0;
rom[23389] = 12'h  0;
rom[23390] = 12'h  0;
rom[23391] = 12'h  0;
rom[23392] = 12'h111;
rom[23393] = 12'h222;
rom[23394] = 12'h333;
rom[23395] = 12'h333;
rom[23396] = 12'h333;
rom[23397] = 12'h333;
rom[23398] = 12'h333;
rom[23399] = 12'h333;
rom[23400] = 12'h433;
rom[23401] = 12'h433;
rom[23402] = 12'h444;
rom[23403] = 12'h666;
rom[23404] = 12'h888;
rom[23405] = 12'ha9a;
rom[23406] = 12'haaa;
rom[23407] = 12'haaa;
rom[23408] = 12'haaa;
rom[23409] = 12'haaa;
rom[23410] = 12'haaa;
rom[23411] = 12'h999;
rom[23412] = 12'h999;
rom[23413] = 12'h999;
rom[23414] = 12'h999;
rom[23415] = 12'h999;
rom[23416] = 12'h999;
rom[23417] = 12'h999;
rom[23418] = 12'h999;
rom[23419] = 12'h999;
rom[23420] = 12'h999;
rom[23421] = 12'h999;
rom[23422] = 12'h888;
rom[23423] = 12'h888;
rom[23424] = 12'h888;
rom[23425] = 12'h888;
rom[23426] = 12'h888;
rom[23427] = 12'h888;
rom[23428] = 12'h888;
rom[23429] = 12'h888;
rom[23430] = 12'h777;
rom[23431] = 12'h777;
rom[23432] = 12'h777;
rom[23433] = 12'h777;
rom[23434] = 12'h777;
rom[23435] = 12'h777;
rom[23436] = 12'h666;
rom[23437] = 12'h666;
rom[23438] = 12'h666;
rom[23439] = 12'h555;
rom[23440] = 12'h555;
rom[23441] = 12'h444;
rom[23442] = 12'h444;
rom[23443] = 12'h333;
rom[23444] = 12'h333;
rom[23445] = 12'h333;
rom[23446] = 12'h222;
rom[23447] = 12'h222;
rom[23448] = 12'h222;
rom[23449] = 12'h111;
rom[23450] = 12'h111;
rom[23451] = 12'h111;
rom[23452] = 12'h111;
rom[23453] = 12'h111;
rom[23454] = 12'h111;
rom[23455] = 12'h111;
rom[23456] = 12'h111;
rom[23457] = 12'h111;
rom[23458] = 12'h111;
rom[23459] = 12'h111;
rom[23460] = 12'h111;
rom[23461] = 12'h111;
rom[23462] = 12'h111;
rom[23463] = 12'h  0;
rom[23464] = 12'h  0;
rom[23465] = 12'h  0;
rom[23466] = 12'h  0;
rom[23467] = 12'h  0;
rom[23468] = 12'h  0;
rom[23469] = 12'h  0;
rom[23470] = 12'h  0;
rom[23471] = 12'h  0;
rom[23472] = 12'h  0;
rom[23473] = 12'h  0;
rom[23474] = 12'h  0;
rom[23475] = 12'h  0;
rom[23476] = 12'h  0;
rom[23477] = 12'h  0;
rom[23478] = 12'h  0;
rom[23479] = 12'h  0;
rom[23480] = 12'h  0;
rom[23481] = 12'h  0;
rom[23482] = 12'h  0;
rom[23483] = 12'h  0;
rom[23484] = 12'h  0;
rom[23485] = 12'h  0;
rom[23486] = 12'h  0;
rom[23487] = 12'h  0;
rom[23488] = 12'h  0;
rom[23489] = 12'h  0;
rom[23490] = 12'h  0;
rom[23491] = 12'h  0;
rom[23492] = 12'h  0;
rom[23493] = 12'h111;
rom[23494] = 12'h111;
rom[23495] = 12'h111;
rom[23496] = 12'h111;
rom[23497] = 12'h111;
rom[23498] = 12'h111;
rom[23499] = 12'h111;
rom[23500] = 12'h222;
rom[23501] = 12'h222;
rom[23502] = 12'h222;
rom[23503] = 12'h333;
rom[23504] = 12'h222;
rom[23505] = 12'h222;
rom[23506] = 12'h333;
rom[23507] = 12'h333;
rom[23508] = 12'h444;
rom[23509] = 12'h444;
rom[23510] = 12'h333;
rom[23511] = 12'h333;
rom[23512] = 12'h333;
rom[23513] = 12'h333;
rom[23514] = 12'h333;
rom[23515] = 12'h333;
rom[23516] = 12'h333;
rom[23517] = 12'h333;
rom[23518] = 12'h333;
rom[23519] = 12'h444;
rom[23520] = 12'h333;
rom[23521] = 12'h444;
rom[23522] = 12'h444;
rom[23523] = 12'h444;
rom[23524] = 12'h444;
rom[23525] = 12'h444;
rom[23526] = 12'h444;
rom[23527] = 12'h444;
rom[23528] = 12'h444;
rom[23529] = 12'h444;
rom[23530] = 12'h444;
rom[23531] = 12'h444;
rom[23532] = 12'h444;
rom[23533] = 12'h444;
rom[23534] = 12'h555;
rom[23535] = 12'h666;
rom[23536] = 12'h666;
rom[23537] = 12'h777;
rom[23538] = 12'h777;
rom[23539] = 12'h888;
rom[23540] = 12'h888;
rom[23541] = 12'h888;
rom[23542] = 12'h888;
rom[23543] = 12'h888;
rom[23544] = 12'h888;
rom[23545] = 12'h888;
rom[23546] = 12'h888;
rom[23547] = 12'h888;
rom[23548] = 12'h877;
rom[23549] = 12'h777;
rom[23550] = 12'h766;
rom[23551] = 12'h666;
rom[23552] = 12'h666;
rom[23553] = 12'h666;
rom[23554] = 12'h666;
rom[23555] = 12'h666;
rom[23556] = 12'h666;
rom[23557] = 12'h666;
rom[23558] = 12'h666;
rom[23559] = 12'h666;
rom[23560] = 12'h666;
rom[23561] = 12'h666;
rom[23562] = 12'h666;
rom[23563] = 12'h766;
rom[23564] = 12'h766;
rom[23565] = 12'h776;
rom[23566] = 12'h776;
rom[23567] = 12'h776;
rom[23568] = 12'h777;
rom[23569] = 12'h777;
rom[23570] = 12'h777;
rom[23571] = 12'h777;
rom[23572] = 12'h777;
rom[23573] = 12'h777;
rom[23574] = 12'h777;
rom[23575] = 12'h666;
rom[23576] = 12'h666;
rom[23577] = 12'h666;
rom[23578] = 12'h666;
rom[23579] = 12'h666;
rom[23580] = 12'h666;
rom[23581] = 12'h666;
rom[23582] = 12'h666;
rom[23583] = 12'h666;
rom[23584] = 12'h777;
rom[23585] = 12'h777;
rom[23586] = 12'h777;
rom[23587] = 12'h777;
rom[23588] = 12'h777;
rom[23589] = 12'h888;
rom[23590] = 12'h888;
rom[23591] = 12'h888;
rom[23592] = 12'h888;
rom[23593] = 12'h888;
rom[23594] = 12'h999;
rom[23595] = 12'h999;
rom[23596] = 12'haaa;
rom[23597] = 12'haaa;
rom[23598] = 12'haaa;
rom[23599] = 12'haaa;
rom[23600] = 12'h777;
rom[23601] = 12'h777;
rom[23602] = 12'h777;
rom[23603] = 12'h777;
rom[23604] = 12'h777;
rom[23605] = 12'h777;
rom[23606] = 12'h777;
rom[23607] = 12'h666;
rom[23608] = 12'h666;
rom[23609] = 12'h666;
rom[23610] = 12'h666;
rom[23611] = 12'h666;
rom[23612] = 12'h666;
rom[23613] = 12'h666;
rom[23614] = 12'h666;
rom[23615] = 12'h666;
rom[23616] = 12'h666;
rom[23617] = 12'h666;
rom[23618] = 12'h666;
rom[23619] = 12'h666;
rom[23620] = 12'h666;
rom[23621] = 12'h666;
rom[23622] = 12'h666;
rom[23623] = 12'h666;
rom[23624] = 12'h666;
rom[23625] = 12'h666;
rom[23626] = 12'h666;
rom[23627] = 12'h666;
rom[23628] = 12'h666;
rom[23629] = 12'h666;
rom[23630] = 12'h666;
rom[23631] = 12'h666;
rom[23632] = 12'h666;
rom[23633] = 12'h666;
rom[23634] = 12'h666;
rom[23635] = 12'h666;
rom[23636] = 12'h666;
rom[23637] = 12'h777;
rom[23638] = 12'h777;
rom[23639] = 12'h777;
rom[23640] = 12'h777;
rom[23641] = 12'h777;
rom[23642] = 12'h777;
rom[23643] = 12'h777;
rom[23644] = 12'h777;
rom[23645] = 12'h777;
rom[23646] = 12'h777;
rom[23647] = 12'h777;
rom[23648] = 12'h777;
rom[23649] = 12'h777;
rom[23650] = 12'h777;
rom[23651] = 12'h777;
rom[23652] = 12'h777;
rom[23653] = 12'h666;
rom[23654] = 12'h666;
rom[23655] = 12'h666;
rom[23656] = 12'h666;
rom[23657] = 12'h666;
rom[23658] = 12'h666;
rom[23659] = 12'h666;
rom[23660] = 12'h666;
rom[23661] = 12'h666;
rom[23662] = 12'h666;
rom[23663] = 12'h666;
rom[23664] = 12'h666;
rom[23665] = 12'h666;
rom[23666] = 12'h666;
rom[23667] = 12'h666;
rom[23668] = 12'h666;
rom[23669] = 12'h666;
rom[23670] = 12'h666;
rom[23671] = 12'h666;
rom[23672] = 12'h555;
rom[23673] = 12'h555;
rom[23674] = 12'h666;
rom[23675] = 12'h666;
rom[23676] = 12'h555;
rom[23677] = 12'h555;
rom[23678] = 12'h555;
rom[23679] = 12'h444;
rom[23680] = 12'h444;
rom[23681] = 12'h444;
rom[23682] = 12'h555;
rom[23683] = 12'h555;
rom[23684] = 12'h555;
rom[23685] = 12'h555;
rom[23686] = 12'h555;
rom[23687] = 12'h555;
rom[23688] = 12'h555;
rom[23689] = 12'h555;
rom[23690] = 12'h555;
rom[23691] = 12'h444;
rom[23692] = 12'h444;
rom[23693] = 12'h333;
rom[23694] = 12'h333;
rom[23695] = 12'h222;
rom[23696] = 12'h111;
rom[23697] = 12'h111;
rom[23698] = 12'h100;
rom[23699] = 12'h  0;
rom[23700] = 12'h  0;
rom[23701] = 12'h  0;
rom[23702] = 12'h  0;
rom[23703] = 12'h  0;
rom[23704] = 12'h  0;
rom[23705] = 12'h  0;
rom[23706] = 12'h  0;
rom[23707] = 12'h  0;
rom[23708] = 12'h  0;
rom[23709] = 12'h  0;
rom[23710] = 12'h  0;
rom[23711] = 12'h  0;
rom[23712] = 12'h100;
rom[23713] = 12'h100;
rom[23714] = 12'h100;
rom[23715] = 12'h100;
rom[23716] = 12'h100;
rom[23717] = 12'h200;
rom[23718] = 12'h200;
rom[23719] = 12'h300;
rom[23720] = 12'h410;
rom[23721] = 12'h510;
rom[23722] = 12'h620;
rom[23723] = 12'h720;
rom[23724] = 12'h930;
rom[23725] = 12'ha40;
rom[23726] = 12'hc51;
rom[23727] = 12'hd61;
rom[23728] = 12'he71;
rom[23729] = 12'hf71;
rom[23730] = 12'hf71;
rom[23731] = 12'hf81;
rom[23732] = 12'hf81;
rom[23733] = 12'hf81;
rom[23734] = 12'hf71;
rom[23735] = 12'hf71;
rom[23736] = 12'hd60;
rom[23737] = 12'hc50;
rom[23738] = 12'hb40;
rom[23739] = 12'h930;
rom[23740] = 12'h820;
rom[23741] = 12'h720;
rom[23742] = 12'h610;
rom[23743] = 12'h500;
rom[23744] = 12'h400;
rom[23745] = 12'h300;
rom[23746] = 12'h300;
rom[23747] = 12'h200;
rom[23748] = 12'h200;
rom[23749] = 12'h200;
rom[23750] = 12'h200;
rom[23751] = 12'h200;
rom[23752] = 12'h200;
rom[23753] = 12'h200;
rom[23754] = 12'h200;
rom[23755] = 12'h300;
rom[23756] = 12'h300;
rom[23757] = 12'h400;
rom[23758] = 12'h400;
rom[23759] = 12'h500;
rom[23760] = 12'h500;
rom[23761] = 12'h600;
rom[23762] = 12'h600;
rom[23763] = 12'h600;
rom[23764] = 12'h600;
rom[23765] = 12'h710;
rom[23766] = 12'h710;
rom[23767] = 12'h710;
rom[23768] = 12'h710;
rom[23769] = 12'h710;
rom[23770] = 12'h710;
rom[23771] = 12'h600;
rom[23772] = 12'h600;
rom[23773] = 12'h500;
rom[23774] = 12'h500;
rom[23775] = 12'h400;
rom[23776] = 12'h400;
rom[23777] = 12'h300;
rom[23778] = 12'h300;
rom[23779] = 12'h300;
rom[23780] = 12'h200;
rom[23781] = 12'h200;
rom[23782] = 12'h200;
rom[23783] = 12'h100;
rom[23784] = 12'h100;
rom[23785] = 12'h100;
rom[23786] = 12'h100;
rom[23787] = 12'h  0;
rom[23788] = 12'h  0;
rom[23789] = 12'h  0;
rom[23790] = 12'h100;
rom[23791] = 12'h100;
rom[23792] = 12'h222;
rom[23793] = 12'h333;
rom[23794] = 12'h333;
rom[23795] = 12'h333;
rom[23796] = 12'h333;
rom[23797] = 12'h233;
rom[23798] = 12'h333;
rom[23799] = 12'h333;
rom[23800] = 12'h333;
rom[23801] = 12'h333;
rom[23802] = 12'h444;
rom[23803] = 12'h555;
rom[23804] = 12'h877;
rom[23805] = 12'h999;
rom[23806] = 12'haaa;
rom[23807] = 12'haaa;
rom[23808] = 12'ha99;
rom[23809] = 12'haaa;
rom[23810] = 12'haaa;
rom[23811] = 12'h999;
rom[23812] = 12'h999;
rom[23813] = 12'h999;
rom[23814] = 12'h999;
rom[23815] = 12'h999;
rom[23816] = 12'h999;
rom[23817] = 12'h999;
rom[23818] = 12'h999;
rom[23819] = 12'h999;
rom[23820] = 12'h999;
rom[23821] = 12'h999;
rom[23822] = 12'h888;
rom[23823] = 12'h888;
rom[23824] = 12'h888;
rom[23825] = 12'h888;
rom[23826] = 12'h888;
rom[23827] = 12'h888;
rom[23828] = 12'h888;
rom[23829] = 12'h888;
rom[23830] = 12'h888;
rom[23831] = 12'h777;
rom[23832] = 12'h777;
rom[23833] = 12'h777;
rom[23834] = 12'h777;
rom[23835] = 12'h666;
rom[23836] = 12'h666;
rom[23837] = 12'h666;
rom[23838] = 12'h555;
rom[23839] = 12'h555;
rom[23840] = 12'h555;
rom[23841] = 12'h444;
rom[23842] = 12'h444;
rom[23843] = 12'h333;
rom[23844] = 12'h333;
rom[23845] = 12'h333;
rom[23846] = 12'h222;
rom[23847] = 12'h222;
rom[23848] = 12'h222;
rom[23849] = 12'h111;
rom[23850] = 12'h111;
rom[23851] = 12'h111;
rom[23852] = 12'h111;
rom[23853] = 12'h111;
rom[23854] = 12'h111;
rom[23855] = 12'h111;
rom[23856] = 12'h111;
rom[23857] = 12'h111;
rom[23858] = 12'h111;
rom[23859] = 12'h111;
rom[23860] = 12'h111;
rom[23861] = 12'h111;
rom[23862] = 12'h  0;
rom[23863] = 12'h  0;
rom[23864] = 12'h  0;
rom[23865] = 12'h  0;
rom[23866] = 12'h  0;
rom[23867] = 12'h  0;
rom[23868] = 12'h  0;
rom[23869] = 12'h  0;
rom[23870] = 12'h  0;
rom[23871] = 12'h  0;
rom[23872] = 12'h  0;
rom[23873] = 12'h  0;
rom[23874] = 12'h  0;
rom[23875] = 12'h  0;
rom[23876] = 12'h  0;
rom[23877] = 12'h  0;
rom[23878] = 12'h  0;
rom[23879] = 12'h  0;
rom[23880] = 12'h  0;
rom[23881] = 12'h  0;
rom[23882] = 12'h  0;
rom[23883] = 12'h  0;
rom[23884] = 12'h  0;
rom[23885] = 12'h  0;
rom[23886] = 12'h  0;
rom[23887] = 12'h  0;
rom[23888] = 12'h  0;
rom[23889] = 12'h  0;
rom[23890] = 12'h  0;
rom[23891] = 12'h  0;
rom[23892] = 12'h  0;
rom[23893] = 12'h111;
rom[23894] = 12'h111;
rom[23895] = 12'h111;
rom[23896] = 12'h111;
rom[23897] = 12'h111;
rom[23898] = 12'h111;
rom[23899] = 12'h222;
rom[23900] = 12'h222;
rom[23901] = 12'h222;
rom[23902] = 12'h222;
rom[23903] = 12'h333;
rom[23904] = 12'h222;
rom[23905] = 12'h222;
rom[23906] = 12'h333;
rom[23907] = 12'h444;
rom[23908] = 12'h444;
rom[23909] = 12'h444;
rom[23910] = 12'h333;
rom[23911] = 12'h333;
rom[23912] = 12'h333;
rom[23913] = 12'h333;
rom[23914] = 12'h444;
rom[23915] = 12'h444;
rom[23916] = 12'h444;
rom[23917] = 12'h444;
rom[23918] = 12'h444;
rom[23919] = 12'h444;
rom[23920] = 12'h444;
rom[23921] = 12'h444;
rom[23922] = 12'h444;
rom[23923] = 12'h444;
rom[23924] = 12'h555;
rom[23925] = 12'h555;
rom[23926] = 12'h555;
rom[23927] = 12'h555;
rom[23928] = 12'h555;
rom[23929] = 12'h555;
rom[23930] = 12'h555;
rom[23931] = 12'h555;
rom[23932] = 12'h555;
rom[23933] = 12'h666;
rom[23934] = 12'h666;
rom[23935] = 12'h777;
rom[23936] = 12'h888;
rom[23937] = 12'h888;
rom[23938] = 12'h888;
rom[23939] = 12'h999;
rom[23940] = 12'h999;
rom[23941] = 12'h999;
rom[23942] = 12'h999;
rom[23943] = 12'h999;
rom[23944] = 12'h888;
rom[23945] = 12'h888;
rom[23946] = 12'h888;
rom[23947] = 12'h877;
rom[23948] = 12'h777;
rom[23949] = 12'h766;
rom[23950] = 12'h666;
rom[23951] = 12'h655;
rom[23952] = 12'h665;
rom[23953] = 12'h665;
rom[23954] = 12'h665;
rom[23955] = 12'h665;
rom[23956] = 12'h665;
rom[23957] = 12'h666;
rom[23958] = 12'h666;
rom[23959] = 12'h666;
rom[23960] = 12'h666;
rom[23961] = 12'h666;
rom[23962] = 12'h766;
rom[23963] = 12'h766;
rom[23964] = 12'h776;
rom[23965] = 12'h776;
rom[23966] = 12'h776;
rom[23967] = 12'h777;
rom[23968] = 12'h777;
rom[23969] = 12'h777;
rom[23970] = 12'h777;
rom[23971] = 12'h777;
rom[23972] = 12'h777;
rom[23973] = 12'h777;
rom[23974] = 12'h777;
rom[23975] = 12'h777;
rom[23976] = 12'h666;
rom[23977] = 12'h666;
rom[23978] = 12'h666;
rom[23979] = 12'h777;
rom[23980] = 12'h777;
rom[23981] = 12'h777;
rom[23982] = 12'h777;
rom[23983] = 12'h777;
rom[23984] = 12'h777;
rom[23985] = 12'h777;
rom[23986] = 12'h777;
rom[23987] = 12'h777;
rom[23988] = 12'h777;
rom[23989] = 12'h888;
rom[23990] = 12'h888;
rom[23991] = 12'h888;
rom[23992] = 12'h888;
rom[23993] = 12'h888;
rom[23994] = 12'h999;
rom[23995] = 12'h999;
rom[23996] = 12'haaa;
rom[23997] = 12'haaa;
rom[23998] = 12'haaa;
rom[23999] = 12'haaa;
rom[24000] = 12'h777;
rom[24001] = 12'h777;
rom[24002] = 12'h777;
rom[24003] = 12'h777;
rom[24004] = 12'h777;
rom[24005] = 12'h777;
rom[24006] = 12'h777;
rom[24007] = 12'h666;
rom[24008] = 12'h666;
rom[24009] = 12'h666;
rom[24010] = 12'h666;
rom[24011] = 12'h666;
rom[24012] = 12'h666;
rom[24013] = 12'h666;
rom[24014] = 12'h666;
rom[24015] = 12'h666;
rom[24016] = 12'h666;
rom[24017] = 12'h666;
rom[24018] = 12'h666;
rom[24019] = 12'h666;
rom[24020] = 12'h666;
rom[24021] = 12'h666;
rom[24022] = 12'h666;
rom[24023] = 12'h666;
rom[24024] = 12'h666;
rom[24025] = 12'h666;
rom[24026] = 12'h666;
rom[24027] = 12'h666;
rom[24028] = 12'h666;
rom[24029] = 12'h666;
rom[24030] = 12'h666;
rom[24031] = 12'h666;
rom[24032] = 12'h666;
rom[24033] = 12'h666;
rom[24034] = 12'h666;
rom[24035] = 12'h666;
rom[24036] = 12'h777;
rom[24037] = 12'h777;
rom[24038] = 12'h777;
rom[24039] = 12'h777;
rom[24040] = 12'h777;
rom[24041] = 12'h777;
rom[24042] = 12'h777;
rom[24043] = 12'h777;
rom[24044] = 12'h777;
rom[24045] = 12'h777;
rom[24046] = 12'h777;
rom[24047] = 12'h777;
rom[24048] = 12'h777;
rom[24049] = 12'h777;
rom[24050] = 12'h777;
rom[24051] = 12'h777;
rom[24052] = 12'h777;
rom[24053] = 12'h777;
rom[24054] = 12'h777;
rom[24055] = 12'h666;
rom[24056] = 12'h666;
rom[24057] = 12'h666;
rom[24058] = 12'h666;
rom[24059] = 12'h666;
rom[24060] = 12'h666;
rom[24061] = 12'h666;
rom[24062] = 12'h666;
rom[24063] = 12'h666;
rom[24064] = 12'h555;
rom[24065] = 12'h555;
rom[24066] = 12'h555;
rom[24067] = 12'h555;
rom[24068] = 12'h555;
rom[24069] = 12'h555;
rom[24070] = 12'h555;
rom[24071] = 12'h555;
rom[24072] = 12'h555;
rom[24073] = 12'h555;
rom[24074] = 12'h555;
rom[24075] = 12'h555;
rom[24076] = 12'h555;
rom[24077] = 12'h555;
rom[24078] = 12'h444;
rom[24079] = 12'h444;
rom[24080] = 12'h444;
rom[24081] = 12'h444;
rom[24082] = 12'h555;
rom[24083] = 12'h555;
rom[24084] = 12'h555;
rom[24085] = 12'h555;
rom[24086] = 12'h555;
rom[24087] = 12'h555;
rom[24088] = 12'h555;
rom[24089] = 12'h555;
rom[24090] = 12'h444;
rom[24091] = 12'h444;
rom[24092] = 12'h444;
rom[24093] = 12'h444;
rom[24094] = 12'h333;
rom[24095] = 12'h333;
rom[24096] = 12'h222;
rom[24097] = 12'h111;
rom[24098] = 12'h111;
rom[24099] = 12'h100;
rom[24100] = 12'h  0;
rom[24101] = 12'h  0;
rom[24102] = 12'h  0;
rom[24103] = 12'h  0;
rom[24104] = 12'h  0;
rom[24105] = 12'h  0;
rom[24106] = 12'h  0;
rom[24107] = 12'h  0;
rom[24108] = 12'h  0;
rom[24109] = 12'h  0;
rom[24110] = 12'h  0;
rom[24111] = 12'h  0;
rom[24112] = 12'h100;
rom[24113] = 12'h100;
rom[24114] = 12'h100;
rom[24115] = 12'h100;
rom[24116] = 12'h100;
rom[24117] = 12'h100;
rom[24118] = 12'h200;
rom[24119] = 12'h200;
rom[24120] = 12'h310;
rom[24121] = 12'h410;
rom[24122] = 12'h620;
rom[24123] = 12'h720;
rom[24124] = 12'h830;
rom[24125] = 12'h940;
rom[24126] = 12'hb51;
rom[24127] = 12'hc61;
rom[24128] = 12'he71;
rom[24129] = 12'he70;
rom[24130] = 12'hf71;
rom[24131] = 12'hf81;
rom[24132] = 12'hf81;
rom[24133] = 12'hf81;
rom[24134] = 12'hf81;
rom[24135] = 12'hf81;
rom[24136] = 12'hf71;
rom[24137] = 12'he71;
rom[24138] = 12'hd61;
rom[24139] = 12'hb50;
rom[24140] = 12'ha40;
rom[24141] = 12'h830;
rom[24142] = 12'h710;
rom[24143] = 12'h510;
rom[24144] = 12'h500;
rom[24145] = 12'h400;
rom[24146] = 12'h400;
rom[24147] = 12'h300;
rom[24148] = 12'h300;
rom[24149] = 12'h300;
rom[24150] = 12'h300;
rom[24151] = 12'h300;
rom[24152] = 12'h300;
rom[24153] = 12'h300;
rom[24154] = 12'h300;
rom[24155] = 12'h400;
rom[24156] = 12'h400;
rom[24157] = 12'h500;
rom[24158] = 12'h500;
rom[24159] = 12'h600;
rom[24160] = 12'h600;
rom[24161] = 12'h600;
rom[24162] = 12'h700;
rom[24163] = 12'h710;
rom[24164] = 12'h710;
rom[24165] = 12'h710;
rom[24166] = 12'h710;
rom[24167] = 12'h710;
rom[24168] = 12'h710;
rom[24169] = 12'h710;
rom[24170] = 12'h710;
rom[24171] = 12'h610;
rom[24172] = 12'h600;
rom[24173] = 12'h500;
rom[24174] = 12'h500;
rom[24175] = 12'h400;
rom[24176] = 12'h400;
rom[24177] = 12'h300;
rom[24178] = 12'h300;
rom[24179] = 12'h300;
rom[24180] = 12'h300;
rom[24181] = 12'h200;
rom[24182] = 12'h200;
rom[24183] = 12'h100;
rom[24184] = 12'h100;
rom[24185] = 12'h100;
rom[24186] = 12'h100;
rom[24187] = 12'h100;
rom[24188] = 12'h  0;
rom[24189] = 12'h  0;
rom[24190] = 12'h100;
rom[24191] = 12'h111;
rom[24192] = 12'h333;
rom[24193] = 12'h333;
rom[24194] = 12'h333;
rom[24195] = 12'h233;
rom[24196] = 12'h222;
rom[24197] = 12'h222;
rom[24198] = 12'h333;
rom[24199] = 12'h333;
rom[24200] = 12'h333;
rom[24201] = 12'h333;
rom[24202] = 12'h444;
rom[24203] = 12'h555;
rom[24204] = 12'h777;
rom[24205] = 12'h999;
rom[24206] = 12'haaa;
rom[24207] = 12'haaa;
rom[24208] = 12'h999;
rom[24209] = 12'h999;
rom[24210] = 12'haaa;
rom[24211] = 12'h999;
rom[24212] = 12'h999;
rom[24213] = 12'h999;
rom[24214] = 12'h999;
rom[24215] = 12'h999;
rom[24216] = 12'h999;
rom[24217] = 12'h999;
rom[24218] = 12'h999;
rom[24219] = 12'h999;
rom[24220] = 12'h999;
rom[24221] = 12'h999;
rom[24222] = 12'h888;
rom[24223] = 12'h888;
rom[24224] = 12'h888;
rom[24225] = 12'h888;
rom[24226] = 12'h888;
rom[24227] = 12'h888;
rom[24228] = 12'h888;
rom[24229] = 12'h888;
rom[24230] = 12'h888;
rom[24231] = 12'h888;
rom[24232] = 12'h777;
rom[24233] = 12'h777;
rom[24234] = 12'h777;
rom[24235] = 12'h666;
rom[24236] = 12'h666;
rom[24237] = 12'h666;
rom[24238] = 12'h555;
rom[24239] = 12'h555;
rom[24240] = 12'h555;
rom[24241] = 12'h444;
rom[24242] = 12'h444;
rom[24243] = 12'h333;
rom[24244] = 12'h333;
rom[24245] = 12'h333;
rom[24246] = 12'h222;
rom[24247] = 12'h222;
rom[24248] = 12'h222;
rom[24249] = 12'h222;
rom[24250] = 12'h111;
rom[24251] = 12'h111;
rom[24252] = 12'h111;
rom[24253] = 12'h111;
rom[24254] = 12'h111;
rom[24255] = 12'h111;
rom[24256] = 12'h222;
rom[24257] = 12'h111;
rom[24258] = 12'h111;
rom[24259] = 12'h111;
rom[24260] = 12'h111;
rom[24261] = 12'h111;
rom[24262] = 12'h  0;
rom[24263] = 12'h  0;
rom[24264] = 12'h  0;
rom[24265] = 12'h  0;
rom[24266] = 12'h  0;
rom[24267] = 12'h  0;
rom[24268] = 12'h  0;
rom[24269] = 12'h  0;
rom[24270] = 12'h  0;
rom[24271] = 12'h  0;
rom[24272] = 12'h  0;
rom[24273] = 12'h  0;
rom[24274] = 12'h  0;
rom[24275] = 12'h  0;
rom[24276] = 12'h  0;
rom[24277] = 12'h  0;
rom[24278] = 12'h  0;
rom[24279] = 12'h  0;
rom[24280] = 12'h  0;
rom[24281] = 12'h  0;
rom[24282] = 12'h  0;
rom[24283] = 12'h  0;
rom[24284] = 12'h  0;
rom[24285] = 12'h  0;
rom[24286] = 12'h  0;
rom[24287] = 12'h  0;
rom[24288] = 12'h  0;
rom[24289] = 12'h  0;
rom[24290] = 12'h  0;
rom[24291] = 12'h  0;
rom[24292] = 12'h  0;
rom[24293] = 12'h111;
rom[24294] = 12'h111;
rom[24295] = 12'h111;
rom[24296] = 12'h111;
rom[24297] = 12'h111;
rom[24298] = 12'h222;
rom[24299] = 12'h222;
rom[24300] = 12'h222;
rom[24301] = 12'h222;
rom[24302] = 12'h222;
rom[24303] = 12'h222;
rom[24304] = 12'h222;
rom[24305] = 12'h333;
rom[24306] = 12'h333;
rom[24307] = 12'h444;
rom[24308] = 12'h444;
rom[24309] = 12'h444;
rom[24310] = 12'h333;
rom[24311] = 12'h333;
rom[24312] = 12'h444;
rom[24313] = 12'h444;
rom[24314] = 12'h444;
rom[24315] = 12'h444;
rom[24316] = 12'h444;
rom[24317] = 12'h444;
rom[24318] = 12'h444;
rom[24319] = 12'h444;
rom[24320] = 12'h444;
rom[24321] = 12'h444;
rom[24322] = 12'h444;
rom[24323] = 12'h555;
rom[24324] = 12'h555;
rom[24325] = 12'h555;
rom[24326] = 12'h555;
rom[24327] = 12'h555;
rom[24328] = 12'h555;
rom[24329] = 12'h555;
rom[24330] = 12'h555;
rom[24331] = 12'h666;
rom[24332] = 12'h666;
rom[24333] = 12'h777;
rom[24334] = 12'h888;
rom[24335] = 12'h888;
rom[24336] = 12'h999;
rom[24337] = 12'h999;
rom[24338] = 12'h999;
rom[24339] = 12'h999;
rom[24340] = 12'ha99;
rom[24341] = 12'h999;
rom[24342] = 12'h999;
rom[24343] = 12'h999;
rom[24344] = 12'h887;
rom[24345] = 12'h877;
rom[24346] = 12'h877;
rom[24347] = 12'h777;
rom[24348] = 12'h877;
rom[24349] = 12'h777;
rom[24350] = 12'h777;
rom[24351] = 12'h766;
rom[24352] = 12'h766;
rom[24353] = 12'h766;
rom[24354] = 12'h766;
rom[24355] = 12'h766;
rom[24356] = 12'h766;
rom[24357] = 12'h766;
rom[24358] = 12'h766;
rom[24359] = 12'h776;
rom[24360] = 12'h776;
rom[24361] = 12'h776;
rom[24362] = 12'h776;
rom[24363] = 12'h776;
rom[24364] = 12'h776;
rom[24365] = 12'h776;
rom[24366] = 12'h777;
rom[24367] = 12'h777;
rom[24368] = 12'h777;
rom[24369] = 12'h777;
rom[24370] = 12'h777;
rom[24371] = 12'h777;
rom[24372] = 12'h777;
rom[24373] = 12'h777;
rom[24374] = 12'h777;
rom[24375] = 12'h777;
rom[24376] = 12'h777;
rom[24377] = 12'h777;
rom[24378] = 12'h777;
rom[24379] = 12'h777;
rom[24380] = 12'h777;
rom[24381] = 12'h777;
rom[24382] = 12'h777;
rom[24383] = 12'h777;
rom[24384] = 12'h777;
rom[24385] = 12'h777;
rom[24386] = 12'h777;
rom[24387] = 12'h777;
rom[24388] = 12'h777;
rom[24389] = 12'h888;
rom[24390] = 12'h888;
rom[24391] = 12'h888;
rom[24392] = 12'h888;
rom[24393] = 12'h888;
rom[24394] = 12'h999;
rom[24395] = 12'h999;
rom[24396] = 12'haaa;
rom[24397] = 12'haaa;
rom[24398] = 12'haaa;
rom[24399] = 12'haaa;
rom[24400] = 12'h777;
rom[24401] = 12'h777;
rom[24402] = 12'h777;
rom[24403] = 12'h777;
rom[24404] = 12'h777;
rom[24405] = 12'h777;
rom[24406] = 12'h777;
rom[24407] = 12'h666;
rom[24408] = 12'h666;
rom[24409] = 12'h666;
rom[24410] = 12'h666;
rom[24411] = 12'h666;
rom[24412] = 12'h666;
rom[24413] = 12'h666;
rom[24414] = 12'h666;
rom[24415] = 12'h666;
rom[24416] = 12'h666;
rom[24417] = 12'h666;
rom[24418] = 12'h666;
rom[24419] = 12'h666;
rom[24420] = 12'h666;
rom[24421] = 12'h666;
rom[24422] = 12'h666;
rom[24423] = 12'h666;
rom[24424] = 12'h666;
rom[24425] = 12'h666;
rom[24426] = 12'h666;
rom[24427] = 12'h666;
rom[24428] = 12'h666;
rom[24429] = 12'h666;
rom[24430] = 12'h666;
rom[24431] = 12'h666;
rom[24432] = 12'h666;
rom[24433] = 12'h666;
rom[24434] = 12'h666;
rom[24435] = 12'h666;
rom[24436] = 12'h777;
rom[24437] = 12'h777;
rom[24438] = 12'h777;
rom[24439] = 12'h777;
rom[24440] = 12'h777;
rom[24441] = 12'h777;
rom[24442] = 12'h777;
rom[24443] = 12'h777;
rom[24444] = 12'h777;
rom[24445] = 12'h777;
rom[24446] = 12'h777;
rom[24447] = 12'h777;
rom[24448] = 12'h888;
rom[24449] = 12'h888;
rom[24450] = 12'h777;
rom[24451] = 12'h777;
rom[24452] = 12'h777;
rom[24453] = 12'h777;
rom[24454] = 12'h777;
rom[24455] = 12'h777;
rom[24456] = 12'h777;
rom[24457] = 12'h666;
rom[24458] = 12'h666;
rom[24459] = 12'h666;
rom[24460] = 12'h666;
rom[24461] = 12'h666;
rom[24462] = 12'h666;
rom[24463] = 12'h666;
rom[24464] = 12'h555;
rom[24465] = 12'h555;
rom[24466] = 12'h555;
rom[24467] = 12'h555;
rom[24468] = 12'h555;
rom[24469] = 12'h555;
rom[24470] = 12'h555;
rom[24471] = 12'h555;
rom[24472] = 12'h555;
rom[24473] = 12'h555;
rom[24474] = 12'h555;
rom[24475] = 12'h555;
rom[24476] = 12'h555;
rom[24477] = 12'h555;
rom[24478] = 12'h444;
rom[24479] = 12'h444;
rom[24480] = 12'h444;
rom[24481] = 12'h444;
rom[24482] = 12'h444;
rom[24483] = 12'h555;
rom[24484] = 12'h555;
rom[24485] = 12'h555;
rom[24486] = 12'h555;
rom[24487] = 12'h444;
rom[24488] = 12'h444;
rom[24489] = 12'h444;
rom[24490] = 12'h444;
rom[24491] = 12'h444;
rom[24492] = 12'h444;
rom[24493] = 12'h333;
rom[24494] = 12'h333;
rom[24495] = 12'h333;
rom[24496] = 12'h222;
rom[24497] = 12'h222;
rom[24498] = 12'h111;
rom[24499] = 12'h111;
rom[24500] = 12'h100;
rom[24501] = 12'h  0;
rom[24502] = 12'h  0;
rom[24503] = 12'h  0;
rom[24504] = 12'h  0;
rom[24505] = 12'h  0;
rom[24506] = 12'h  0;
rom[24507] = 12'h  0;
rom[24508] = 12'h  0;
rom[24509] = 12'h  0;
rom[24510] = 12'h  0;
rom[24511] = 12'h  0;
rom[24512] = 12'h100;
rom[24513] = 12'h100;
rom[24514] = 12'h100;
rom[24515] = 12'h100;
rom[24516] = 12'h100;
rom[24517] = 12'h100;
rom[24518] = 12'h200;
rom[24519] = 12'h200;
rom[24520] = 12'h310;
rom[24521] = 12'h410;
rom[24522] = 12'h520;
rom[24523] = 12'h620;
rom[24524] = 12'h830;
rom[24525] = 12'h930;
rom[24526] = 12'ha40;
rom[24527] = 12'hb50;
rom[24528] = 12'hd71;
rom[24529] = 12'he70;
rom[24530] = 12'he80;
rom[24531] = 12'hf81;
rom[24532] = 12'hf81;
rom[24533] = 12'hf81;
rom[24534] = 12'hf81;
rom[24535] = 12'hf91;
rom[24536] = 12'hf81;
rom[24537] = 12'hf81;
rom[24538] = 12'he71;
rom[24539] = 12'hd71;
rom[24540] = 12'hc61;
rom[24541] = 12'ha40;
rom[24542] = 12'h930;
rom[24543] = 12'h720;
rom[24544] = 12'h610;
rom[24545] = 12'h510;
rom[24546] = 12'h400;
rom[24547] = 12'h400;
rom[24548] = 12'h400;
rom[24549] = 12'h400;
rom[24550] = 12'h400;
rom[24551] = 12'h300;
rom[24552] = 12'h400;
rom[24553] = 12'h400;
rom[24554] = 12'h400;
rom[24555] = 12'h500;
rom[24556] = 12'h500;
rom[24557] = 12'h600;
rom[24558] = 12'h600;
rom[24559] = 12'h700;
rom[24560] = 12'h700;
rom[24561] = 12'h710;
rom[24562] = 12'h810;
rom[24563] = 12'h810;
rom[24564] = 12'h810;
rom[24565] = 12'h810;
rom[24566] = 12'h810;
rom[24567] = 12'h810;
rom[24568] = 12'h810;
rom[24569] = 12'h810;
rom[24570] = 12'h710;
rom[24571] = 12'h710;
rom[24572] = 12'h600;
rom[24573] = 12'h600;
rom[24574] = 12'h500;
rom[24575] = 12'h500;
rom[24576] = 12'h400;
rom[24577] = 12'h300;
rom[24578] = 12'h300;
rom[24579] = 12'h300;
rom[24580] = 12'h300;
rom[24581] = 12'h200;
rom[24582] = 12'h200;
rom[24583] = 12'h100;
rom[24584] = 12'h100;
rom[24585] = 12'h100;
rom[24586] = 12'h100;
rom[24587] = 12'h100;
rom[24588] = 12'h  0;
rom[24589] = 12'h100;
rom[24590] = 12'h211;
rom[24591] = 12'h212;
rom[24592] = 12'h333;
rom[24593] = 12'h233;
rom[24594] = 12'h222;
rom[24595] = 12'h222;
rom[24596] = 12'h222;
rom[24597] = 12'h222;
rom[24598] = 12'h233;
rom[24599] = 12'h333;
rom[24600] = 12'h333;
rom[24601] = 12'h333;
rom[24602] = 12'h444;
rom[24603] = 12'h555;
rom[24604] = 12'h766;
rom[24605] = 12'h999;
rom[24606] = 12'haaa;
rom[24607] = 12'haaa;
rom[24608] = 12'h999;
rom[24609] = 12'h999;
rom[24610] = 12'h999;
rom[24611] = 12'haaa;
rom[24612] = 12'h999;
rom[24613] = 12'h999;
rom[24614] = 12'h888;
rom[24615] = 12'h999;
rom[24616] = 12'h999;
rom[24617] = 12'h999;
rom[24618] = 12'h999;
rom[24619] = 12'h999;
rom[24620] = 12'h999;
rom[24621] = 12'h999;
rom[24622] = 12'h888;
rom[24623] = 12'h888;
rom[24624] = 12'h888;
rom[24625] = 12'h888;
rom[24626] = 12'h888;
rom[24627] = 12'h888;
rom[24628] = 12'h888;
rom[24629] = 12'h888;
rom[24630] = 12'h888;
rom[24631] = 12'h777;
rom[24632] = 12'h777;
rom[24633] = 12'h777;
rom[24634] = 12'h777;
rom[24635] = 12'h666;
rom[24636] = 12'h666;
rom[24637] = 12'h666;
rom[24638] = 12'h555;
rom[24639] = 12'h555;
rom[24640] = 12'h444;
rom[24641] = 12'h444;
rom[24642] = 12'h444;
rom[24643] = 12'h333;
rom[24644] = 12'h333;
rom[24645] = 12'h333;
rom[24646] = 12'h222;
rom[24647] = 12'h222;
rom[24648] = 12'h222;
rom[24649] = 12'h222;
rom[24650] = 12'h222;
rom[24651] = 12'h222;
rom[24652] = 12'h222;
rom[24653] = 12'h222;
rom[24654] = 12'h222;
rom[24655] = 12'h111;
rom[24656] = 12'h111;
rom[24657] = 12'h111;
rom[24658] = 12'h111;
rom[24659] = 12'h111;
rom[24660] = 12'h111;
rom[24661] = 12'h  0;
rom[24662] = 12'h  0;
rom[24663] = 12'h  0;
rom[24664] = 12'h  0;
rom[24665] = 12'h  0;
rom[24666] = 12'h  0;
rom[24667] = 12'h  0;
rom[24668] = 12'h  0;
rom[24669] = 12'h  0;
rom[24670] = 12'h  0;
rom[24671] = 12'h  0;
rom[24672] = 12'h  0;
rom[24673] = 12'h  0;
rom[24674] = 12'h  0;
rom[24675] = 12'h  0;
rom[24676] = 12'h  0;
rom[24677] = 12'h  0;
rom[24678] = 12'h  0;
rom[24679] = 12'h  0;
rom[24680] = 12'h  0;
rom[24681] = 12'h  0;
rom[24682] = 12'h  0;
rom[24683] = 12'h  0;
rom[24684] = 12'h  0;
rom[24685] = 12'h  0;
rom[24686] = 12'h  0;
rom[24687] = 12'h  0;
rom[24688] = 12'h  0;
rom[24689] = 12'h  0;
rom[24690] = 12'h  0;
rom[24691] = 12'h  0;
rom[24692] = 12'h111;
rom[24693] = 12'h111;
rom[24694] = 12'h111;
rom[24695] = 12'h111;
rom[24696] = 12'h111;
rom[24697] = 12'h111;
rom[24698] = 12'h222;
rom[24699] = 12'h222;
rom[24700] = 12'h222;
rom[24701] = 12'h222;
rom[24702] = 12'h222;
rom[24703] = 12'h222;
rom[24704] = 12'h222;
rom[24705] = 12'h333;
rom[24706] = 12'h444;
rom[24707] = 12'h444;
rom[24708] = 12'h444;
rom[24709] = 12'h444;
rom[24710] = 12'h333;
rom[24711] = 12'h333;
rom[24712] = 12'h444;
rom[24713] = 12'h444;
rom[24714] = 12'h444;
rom[24715] = 12'h444;
rom[24716] = 12'h444;
rom[24717] = 12'h444;
rom[24718] = 12'h444;
rom[24719] = 12'h444;
rom[24720] = 12'h444;
rom[24721] = 12'h555;
rom[24722] = 12'h555;
rom[24723] = 12'h555;
rom[24724] = 12'h555;
rom[24725] = 12'h555;
rom[24726] = 12'h555;
rom[24727] = 12'h555;
rom[24728] = 12'h666;
rom[24729] = 12'h666;
rom[24730] = 12'h666;
rom[24731] = 12'h777;
rom[24732] = 12'h888;
rom[24733] = 12'h888;
rom[24734] = 12'h999;
rom[24735] = 12'h999;
rom[24736] = 12'haaa;
rom[24737] = 12'haaa;
rom[24738] = 12'haaa;
rom[24739] = 12'haaa;
rom[24740] = 12'ha99;
rom[24741] = 12'h999;
rom[24742] = 12'h999;
rom[24743] = 12'h988;
rom[24744] = 12'h888;
rom[24745] = 12'h877;
rom[24746] = 12'h877;
rom[24747] = 12'h877;
rom[24748] = 12'h877;
rom[24749] = 12'h888;
rom[24750] = 12'h888;
rom[24751] = 12'h888;
rom[24752] = 12'h877;
rom[24753] = 12'h777;
rom[24754] = 12'h777;
rom[24755] = 12'h777;
rom[24756] = 12'h777;
rom[24757] = 12'h777;
rom[24758] = 12'h777;
rom[24759] = 12'h777;
rom[24760] = 12'h776;
rom[24761] = 12'h776;
rom[24762] = 12'h776;
rom[24763] = 12'h777;
rom[24764] = 12'h777;
rom[24765] = 12'h777;
rom[24766] = 12'h777;
rom[24767] = 12'h777;
rom[24768] = 12'h777;
rom[24769] = 12'h777;
rom[24770] = 12'h888;
rom[24771] = 12'h888;
rom[24772] = 12'h888;
rom[24773] = 12'h888;
rom[24774] = 12'h888;
rom[24775] = 12'h888;
rom[24776] = 12'h888;
rom[24777] = 12'h888;
rom[24778] = 12'h777;
rom[24779] = 12'h777;
rom[24780] = 12'h777;
rom[24781] = 12'h777;
rom[24782] = 12'h777;
rom[24783] = 12'h777;
rom[24784] = 12'h777;
rom[24785] = 12'h777;
rom[24786] = 12'h777;
rom[24787] = 12'h777;
rom[24788] = 12'h888;
rom[24789] = 12'h888;
rom[24790] = 12'h888;
rom[24791] = 12'h888;
rom[24792] = 12'h888;
rom[24793] = 12'h888;
rom[24794] = 12'h999;
rom[24795] = 12'h999;
rom[24796] = 12'haaa;
rom[24797] = 12'haaa;
rom[24798] = 12'haaa;
rom[24799] = 12'haaa;
rom[24800] = 12'h777;
rom[24801] = 12'h777;
rom[24802] = 12'h777;
rom[24803] = 12'h777;
rom[24804] = 12'h777;
rom[24805] = 12'h777;
rom[24806] = 12'h777;
rom[24807] = 12'h777;
rom[24808] = 12'h666;
rom[24809] = 12'h666;
rom[24810] = 12'h666;
rom[24811] = 12'h666;
rom[24812] = 12'h666;
rom[24813] = 12'h666;
rom[24814] = 12'h666;
rom[24815] = 12'h666;
rom[24816] = 12'h666;
rom[24817] = 12'h666;
rom[24818] = 12'h666;
rom[24819] = 12'h666;
rom[24820] = 12'h666;
rom[24821] = 12'h666;
rom[24822] = 12'h666;
rom[24823] = 12'h666;
rom[24824] = 12'h666;
rom[24825] = 12'h666;
rom[24826] = 12'h666;
rom[24827] = 12'h666;
rom[24828] = 12'h666;
rom[24829] = 12'h666;
rom[24830] = 12'h666;
rom[24831] = 12'h666;
rom[24832] = 12'h777;
rom[24833] = 12'h777;
rom[24834] = 12'h777;
rom[24835] = 12'h777;
rom[24836] = 12'h777;
rom[24837] = 12'h777;
rom[24838] = 12'h777;
rom[24839] = 12'h777;
rom[24840] = 12'h888;
rom[24841] = 12'h777;
rom[24842] = 12'h777;
rom[24843] = 12'h777;
rom[24844] = 12'h777;
rom[24845] = 12'h777;
rom[24846] = 12'h777;
rom[24847] = 12'h888;
rom[24848] = 12'h888;
rom[24849] = 12'h888;
rom[24850] = 12'h888;
rom[24851] = 12'h888;
rom[24852] = 12'h777;
rom[24853] = 12'h777;
rom[24854] = 12'h777;
rom[24855] = 12'h777;
rom[24856] = 12'h777;
rom[24857] = 12'h666;
rom[24858] = 12'h666;
rom[24859] = 12'h666;
rom[24860] = 12'h666;
rom[24861] = 12'h666;
rom[24862] = 12'h666;
rom[24863] = 12'h666;
rom[24864] = 12'h555;
rom[24865] = 12'h555;
rom[24866] = 12'h555;
rom[24867] = 12'h555;
rom[24868] = 12'h555;
rom[24869] = 12'h555;
rom[24870] = 12'h555;
rom[24871] = 12'h555;
rom[24872] = 12'h555;
rom[24873] = 12'h555;
rom[24874] = 12'h555;
rom[24875] = 12'h555;
rom[24876] = 12'h555;
rom[24877] = 12'h555;
rom[24878] = 12'h444;
rom[24879] = 12'h444;
rom[24880] = 12'h444;
rom[24881] = 12'h444;
rom[24882] = 12'h444;
rom[24883] = 12'h444;
rom[24884] = 12'h444;
rom[24885] = 12'h444;
rom[24886] = 12'h444;
rom[24887] = 12'h444;
rom[24888] = 12'h444;
rom[24889] = 12'h444;
rom[24890] = 12'h444;
rom[24891] = 12'h444;
rom[24892] = 12'h444;
rom[24893] = 12'h333;
rom[24894] = 12'h333;
rom[24895] = 12'h333;
rom[24896] = 12'h322;
rom[24897] = 12'h222;
rom[24898] = 12'h222;
rom[24899] = 12'h111;
rom[24900] = 12'h111;
rom[24901] = 12'h100;
rom[24902] = 12'h  0;
rom[24903] = 12'h  0;
rom[24904] = 12'h  0;
rom[24905] = 12'h  0;
rom[24906] = 12'h  0;
rom[24907] = 12'h  0;
rom[24908] = 12'h  0;
rom[24909] = 12'h  0;
rom[24910] = 12'h  0;
rom[24911] = 12'h  0;
rom[24912] = 12'h100;
rom[24913] = 12'h100;
rom[24914] = 12'h100;
rom[24915] = 12'h100;
rom[24916] = 12'h100;
rom[24917] = 12'h100;
rom[24918] = 12'h100;
rom[24919] = 12'h200;
rom[24920] = 12'h200;
rom[24921] = 12'h310;
rom[24922] = 12'h510;
rom[24923] = 12'h620;
rom[24924] = 12'h720;
rom[24925] = 12'h830;
rom[24926] = 12'h930;
rom[24927] = 12'ha40;
rom[24928] = 12'hc60;
rom[24929] = 12'hd70;
rom[24930] = 12'he70;
rom[24931] = 12'hf80;
rom[24932] = 12'hf81;
rom[24933] = 12'hf91;
rom[24934] = 12'hf91;
rom[24935] = 12'hf91;
rom[24936] = 12'hf91;
rom[24937] = 12'hf81;
rom[24938] = 12'hf82;
rom[24939] = 12'he82;
rom[24940] = 12'hd72;
rom[24941] = 12'hc61;
rom[24942] = 12'hb51;
rom[24943] = 12'ha41;
rom[24944] = 12'h831;
rom[24945] = 12'h720;
rom[24946] = 12'h610;
rom[24947] = 12'h510;
rom[24948] = 12'h510;
rom[24949] = 12'h510;
rom[24950] = 12'h510;
rom[24951] = 12'h410;
rom[24952] = 12'h510;
rom[24953] = 12'h510;
rom[24954] = 12'h610;
rom[24955] = 12'h610;
rom[24956] = 12'h710;
rom[24957] = 12'h710;
rom[24958] = 12'h710;
rom[24959] = 12'h810;
rom[24960] = 12'h810;
rom[24961] = 12'h810;
rom[24962] = 12'h810;
rom[24963] = 12'h910;
rom[24964] = 12'h910;
rom[24965] = 12'h910;
rom[24966] = 12'h910;
rom[24967] = 12'h810;
rom[24968] = 12'h810;
rom[24969] = 12'h810;
rom[24970] = 12'h710;
rom[24971] = 12'h710;
rom[24972] = 12'h610;
rom[24973] = 12'h600;
rom[24974] = 12'h500;
rom[24975] = 12'h500;
rom[24976] = 12'h400;
rom[24977] = 12'h400;
rom[24978] = 12'h300;
rom[24979] = 12'h300;
rom[24980] = 12'h300;
rom[24981] = 12'h200;
rom[24982] = 12'h200;
rom[24983] = 12'h100;
rom[24984] = 12'h100;
rom[24985] = 12'h100;
rom[24986] = 12'h100;
rom[24987] = 12'h100;
rom[24988] = 12'h100;
rom[24989] = 12'h100;
rom[24990] = 12'h211;
rom[24991] = 12'h322;
rom[24992] = 12'h233;
rom[24993] = 12'h222;
rom[24994] = 12'h122;
rom[24995] = 12'h122;
rom[24996] = 12'h222;
rom[24997] = 12'h232;
rom[24998] = 12'h333;
rom[24999] = 12'h233;
rom[25000] = 12'h333;
rom[25001] = 12'h333;
rom[25002] = 12'h444;
rom[25003] = 12'h544;
rom[25004] = 12'h766;
rom[25005] = 12'h988;
rom[25006] = 12'ha9a;
rom[25007] = 12'ha99;
rom[25008] = 12'h999;
rom[25009] = 12'h999;
rom[25010] = 12'h999;
rom[25011] = 12'haaa;
rom[25012] = 12'h999;
rom[25013] = 12'h999;
rom[25014] = 12'h888;
rom[25015] = 12'h999;
rom[25016] = 12'h999;
rom[25017] = 12'h999;
rom[25018] = 12'h999;
rom[25019] = 12'h888;
rom[25020] = 12'h888;
rom[25021] = 12'h888;
rom[25022] = 12'h888;
rom[25023] = 12'h888;
rom[25024] = 12'h888;
rom[25025] = 12'h888;
rom[25026] = 12'h888;
rom[25027] = 12'h888;
rom[25028] = 12'h888;
rom[25029] = 12'h888;
rom[25030] = 12'h777;
rom[25031] = 12'h777;
rom[25032] = 12'h777;
rom[25033] = 12'h777;
rom[25034] = 12'h777;
rom[25035] = 12'h666;
rom[25036] = 12'h666;
rom[25037] = 12'h666;
rom[25038] = 12'h555;
rom[25039] = 12'h555;
rom[25040] = 12'h444;
rom[25041] = 12'h444;
rom[25042] = 12'h444;
rom[25043] = 12'h333;
rom[25044] = 12'h333;
rom[25045] = 12'h333;
rom[25046] = 12'h222;
rom[25047] = 12'h222;
rom[25048] = 12'h222;
rom[25049] = 12'h222;
rom[25050] = 12'h222;
rom[25051] = 12'h222;
rom[25052] = 12'h222;
rom[25053] = 12'h222;
rom[25054] = 12'h222;
rom[25055] = 12'h222;
rom[25056] = 12'h111;
rom[25057] = 12'h111;
rom[25058] = 12'h  0;
rom[25059] = 12'h  0;
rom[25060] = 12'h  0;
rom[25061] = 12'h  0;
rom[25062] = 12'h  0;
rom[25063] = 12'h  0;
rom[25064] = 12'h  0;
rom[25065] = 12'h  0;
rom[25066] = 12'h  0;
rom[25067] = 12'h  0;
rom[25068] = 12'h  0;
rom[25069] = 12'h  0;
rom[25070] = 12'h  0;
rom[25071] = 12'h  0;
rom[25072] = 12'h  0;
rom[25073] = 12'h  0;
rom[25074] = 12'h  0;
rom[25075] = 12'h  0;
rom[25076] = 12'h  0;
rom[25077] = 12'h  0;
rom[25078] = 12'h  0;
rom[25079] = 12'h  0;
rom[25080] = 12'h  0;
rom[25081] = 12'h  0;
rom[25082] = 12'h  0;
rom[25083] = 12'h  0;
rom[25084] = 12'h  0;
rom[25085] = 12'h  0;
rom[25086] = 12'h  0;
rom[25087] = 12'h  0;
rom[25088] = 12'h  0;
rom[25089] = 12'h  0;
rom[25090] = 12'h  0;
rom[25091] = 12'h  0;
rom[25092] = 12'h111;
rom[25093] = 12'h111;
rom[25094] = 12'h111;
rom[25095] = 12'h111;
rom[25096] = 12'h111;
rom[25097] = 12'h111;
rom[25098] = 12'h222;
rom[25099] = 12'h222;
rom[25100] = 12'h222;
rom[25101] = 12'h222;
rom[25102] = 12'h222;
rom[25103] = 12'h222;
rom[25104] = 12'h222;
rom[25105] = 12'h333;
rom[25106] = 12'h444;
rom[25107] = 12'h444;
rom[25108] = 12'h444;
rom[25109] = 12'h333;
rom[25110] = 12'h333;
rom[25111] = 12'h444;
rom[25112] = 12'h444;
rom[25113] = 12'h444;
rom[25114] = 12'h444;
rom[25115] = 12'h444;
rom[25116] = 12'h444;
rom[25117] = 12'h444;
rom[25118] = 12'h444;
rom[25119] = 12'h444;
rom[25120] = 12'h555;
rom[25121] = 12'h555;
rom[25122] = 12'h555;
rom[25123] = 12'h555;
rom[25124] = 12'h666;
rom[25125] = 12'h666;
rom[25126] = 12'h666;
rom[25127] = 12'h666;
rom[25128] = 12'h777;
rom[25129] = 12'h777;
rom[25130] = 12'h888;
rom[25131] = 12'h999;
rom[25132] = 12'h999;
rom[25133] = 12'haaa;
rom[25134] = 12'haaa;
rom[25135] = 12'hbbb;
rom[25136] = 12'hbbb;
rom[25137] = 12'hbbb;
rom[25138] = 12'hbba;
rom[25139] = 12'haaa;
rom[25140] = 12'haaa;
rom[25141] = 12'ha99;
rom[25142] = 12'h999;
rom[25143] = 12'h999;
rom[25144] = 12'h999;
rom[25145] = 12'h988;
rom[25146] = 12'h888;
rom[25147] = 12'h888;
rom[25148] = 12'h888;
rom[25149] = 12'h888;
rom[25150] = 12'h888;
rom[25151] = 12'h888;
rom[25152] = 12'h877;
rom[25153] = 12'h777;
rom[25154] = 12'h777;
rom[25155] = 12'h776;
rom[25156] = 12'h776;
rom[25157] = 12'h766;
rom[25158] = 12'h766;
rom[25159] = 12'h766;
rom[25160] = 12'h766;
rom[25161] = 12'h766;
rom[25162] = 12'h776;
rom[25163] = 12'h776;
rom[25164] = 12'h776;
rom[25165] = 12'h777;
rom[25166] = 12'h777;
rom[25167] = 12'h777;
rom[25168] = 12'h777;
rom[25169] = 12'h777;
rom[25170] = 12'h777;
rom[25171] = 12'h888;
rom[25172] = 12'h888;
rom[25173] = 12'h888;
rom[25174] = 12'h888;
rom[25175] = 12'h888;
rom[25176] = 12'h888;
rom[25177] = 12'h888;
rom[25178] = 12'h888;
rom[25179] = 12'h888;
rom[25180] = 12'h888;
rom[25181] = 12'h888;
rom[25182] = 12'h777;
rom[25183] = 12'h777;
rom[25184] = 12'h777;
rom[25185] = 12'h777;
rom[25186] = 12'h777;
rom[25187] = 12'h888;
rom[25188] = 12'h888;
rom[25189] = 12'h888;
rom[25190] = 12'h888;
rom[25191] = 12'h888;
rom[25192] = 12'h888;
rom[25193] = 12'h888;
rom[25194] = 12'h999;
rom[25195] = 12'h999;
rom[25196] = 12'haaa;
rom[25197] = 12'haaa;
rom[25198] = 12'haaa;
rom[25199] = 12'haaa;
rom[25200] = 12'h777;
rom[25201] = 12'h777;
rom[25202] = 12'h777;
rom[25203] = 12'h777;
rom[25204] = 12'h777;
rom[25205] = 12'h777;
rom[25206] = 12'h777;
rom[25207] = 12'h777;
rom[25208] = 12'h777;
rom[25209] = 12'h777;
rom[25210] = 12'h666;
rom[25211] = 12'h666;
rom[25212] = 12'h666;
rom[25213] = 12'h666;
rom[25214] = 12'h666;
rom[25215] = 12'h666;
rom[25216] = 12'h666;
rom[25217] = 12'h666;
rom[25218] = 12'h666;
rom[25219] = 12'h666;
rom[25220] = 12'h666;
rom[25221] = 12'h777;
rom[25222] = 12'h777;
rom[25223] = 12'h777;
rom[25224] = 12'h777;
rom[25225] = 12'h777;
rom[25226] = 12'h777;
rom[25227] = 12'h777;
rom[25228] = 12'h777;
rom[25229] = 12'h777;
rom[25230] = 12'h777;
rom[25231] = 12'h777;
rom[25232] = 12'h777;
rom[25233] = 12'h777;
rom[25234] = 12'h777;
rom[25235] = 12'h777;
rom[25236] = 12'h777;
rom[25237] = 12'h777;
rom[25238] = 12'h777;
rom[25239] = 12'h777;
rom[25240] = 12'h888;
rom[25241] = 12'h888;
rom[25242] = 12'h777;
rom[25243] = 12'h777;
rom[25244] = 12'h777;
rom[25245] = 12'h777;
rom[25246] = 12'h888;
rom[25247] = 12'h888;
rom[25248] = 12'h888;
rom[25249] = 12'h888;
rom[25250] = 12'h888;
rom[25251] = 12'h888;
rom[25252] = 12'h888;
rom[25253] = 12'h777;
rom[25254] = 12'h777;
rom[25255] = 12'h777;
rom[25256] = 12'h777;
rom[25257] = 12'h666;
rom[25258] = 12'h666;
rom[25259] = 12'h666;
rom[25260] = 12'h666;
rom[25261] = 12'h666;
rom[25262] = 12'h666;
rom[25263] = 12'h666;
rom[25264] = 12'h555;
rom[25265] = 12'h555;
rom[25266] = 12'h555;
rom[25267] = 12'h555;
rom[25268] = 12'h555;
rom[25269] = 12'h555;
rom[25270] = 12'h555;
rom[25271] = 12'h555;
rom[25272] = 12'h555;
rom[25273] = 12'h555;
rom[25274] = 12'h555;
rom[25275] = 12'h555;
rom[25276] = 12'h555;
rom[25277] = 12'h555;
rom[25278] = 12'h444;
rom[25279] = 12'h444;
rom[25280] = 12'h444;
rom[25281] = 12'h444;
rom[25282] = 12'h444;
rom[25283] = 12'h444;
rom[25284] = 12'h444;
rom[25285] = 12'h444;
rom[25286] = 12'h444;
rom[25287] = 12'h444;
rom[25288] = 12'h444;
rom[25289] = 12'h444;
rom[25290] = 12'h444;
rom[25291] = 12'h444;
rom[25292] = 12'h333;
rom[25293] = 12'h333;
rom[25294] = 12'h222;
rom[25295] = 12'h222;
rom[25296] = 12'h333;
rom[25297] = 12'h222;
rom[25298] = 12'h222;
rom[25299] = 12'h111;
rom[25300] = 12'h111;
rom[25301] = 12'h100;
rom[25302] = 12'h  0;
rom[25303] = 12'h  0;
rom[25304] = 12'h  0;
rom[25305] = 12'h  0;
rom[25306] = 12'h  0;
rom[25307] = 12'h  0;
rom[25308] = 12'h  0;
rom[25309] = 12'h  0;
rom[25310] = 12'h  0;
rom[25311] = 12'h  0;
rom[25312] = 12'h  0;
rom[25313] = 12'h100;
rom[25314] = 12'h100;
rom[25315] = 12'h  0;
rom[25316] = 12'h  0;
rom[25317] = 12'h100;
rom[25318] = 12'h100;
rom[25319] = 12'h200;
rom[25320] = 12'h200;
rom[25321] = 12'h300;
rom[25322] = 12'h410;
rom[25323] = 12'h510;
rom[25324] = 12'h610;
rom[25325] = 12'h720;
rom[25326] = 12'h820;
rom[25327] = 12'h930;
rom[25328] = 12'hb50;
rom[25329] = 12'hc60;
rom[25330] = 12'hd70;
rom[25331] = 12'he81;
rom[25332] = 12'hf81;
rom[25333] = 12'hf81;
rom[25334] = 12'hf81;
rom[25335] = 12'hf91;
rom[25336] = 12'hf91;
rom[25337] = 12'hf91;
rom[25338] = 12'hf91;
rom[25339] = 12'hf82;
rom[25340] = 12'hf82;
rom[25341] = 12'he82;
rom[25342] = 12'he72;
rom[25343] = 12'hd72;
rom[25344] = 12'hb51;
rom[25345] = 12'ha41;
rom[25346] = 12'h830;
rom[25347] = 12'h820;
rom[25348] = 12'h720;
rom[25349] = 12'h720;
rom[25350] = 12'h720;
rom[25351] = 12'h720;
rom[25352] = 12'h720;
rom[25353] = 12'h720;
rom[25354] = 12'h820;
rom[25355] = 12'h820;
rom[25356] = 12'h810;
rom[25357] = 12'h810;
rom[25358] = 12'h810;
rom[25359] = 12'h910;
rom[25360] = 12'h910;
rom[25361] = 12'h910;
rom[25362] = 12'h910;
rom[25363] = 12'ha20;
rom[25364] = 12'h920;
rom[25365] = 12'h920;
rom[25366] = 12'h920;
rom[25367] = 12'h920;
rom[25368] = 12'h810;
rom[25369] = 12'h810;
rom[25370] = 12'h710;
rom[25371] = 12'h710;
rom[25372] = 12'h610;
rom[25373] = 12'h610;
rom[25374] = 12'h500;
rom[25375] = 12'h500;
rom[25376] = 12'h400;
rom[25377] = 12'h400;
rom[25378] = 12'h300;
rom[25379] = 12'h300;
rom[25380] = 12'h300;
rom[25381] = 12'h200;
rom[25382] = 12'h200;
rom[25383] = 12'h100;
rom[25384] = 12'h100;
rom[25385] = 12'h100;
rom[25386] = 12'h100;
rom[25387] = 12'h100;
rom[25388] = 12'h100;
rom[25389] = 12'h101;
rom[25390] = 12'h212;
rom[25391] = 12'h323;
rom[25392] = 12'h222;
rom[25393] = 12'h122;
rom[25394] = 12'h111;
rom[25395] = 12'h111;
rom[25396] = 12'h222;
rom[25397] = 12'h233;
rom[25398] = 12'h333;
rom[25399] = 12'h222;
rom[25400] = 12'h333;
rom[25401] = 12'h333;
rom[25402] = 12'h444;
rom[25403] = 12'h444;
rom[25404] = 12'h666;
rom[25405] = 12'h988;
rom[25406] = 12'ha99;
rom[25407] = 12'h999;
rom[25408] = 12'h999;
rom[25409] = 12'h999;
rom[25410] = 12'h999;
rom[25411] = 12'haaa;
rom[25412] = 12'h999;
rom[25413] = 12'h888;
rom[25414] = 12'h888;
rom[25415] = 12'h999;
rom[25416] = 12'h999;
rom[25417] = 12'h999;
rom[25418] = 12'h888;
rom[25419] = 12'h888;
rom[25420] = 12'h888;
rom[25421] = 12'h888;
rom[25422] = 12'h888;
rom[25423] = 12'h888;
rom[25424] = 12'h888;
rom[25425] = 12'h888;
rom[25426] = 12'h888;
rom[25427] = 12'h888;
rom[25428] = 12'h888;
rom[25429] = 12'h777;
rom[25430] = 12'h777;
rom[25431] = 12'h777;
rom[25432] = 12'h777;
rom[25433] = 12'h666;
rom[25434] = 12'h666;
rom[25435] = 12'h666;
rom[25436] = 12'h666;
rom[25437] = 12'h555;
rom[25438] = 12'h555;
rom[25439] = 12'h555;
rom[25440] = 12'h444;
rom[25441] = 12'h444;
rom[25442] = 12'h444;
rom[25443] = 12'h333;
rom[25444] = 12'h333;
rom[25445] = 12'h333;
rom[25446] = 12'h222;
rom[25447] = 12'h222;
rom[25448] = 12'h222;
rom[25449] = 12'h222;
rom[25450] = 12'h222;
rom[25451] = 12'h222;
rom[25452] = 12'h222;
rom[25453] = 12'h222;
rom[25454] = 12'h222;
rom[25455] = 12'h222;
rom[25456] = 12'h111;
rom[25457] = 12'h111;
rom[25458] = 12'h  0;
rom[25459] = 12'h  0;
rom[25460] = 12'h  0;
rom[25461] = 12'h  0;
rom[25462] = 12'h  0;
rom[25463] = 12'h  0;
rom[25464] = 12'h  0;
rom[25465] = 12'h  0;
rom[25466] = 12'h  0;
rom[25467] = 12'h  0;
rom[25468] = 12'h  0;
rom[25469] = 12'h  0;
rom[25470] = 12'h  0;
rom[25471] = 12'h  0;
rom[25472] = 12'h  0;
rom[25473] = 12'h  0;
rom[25474] = 12'h  0;
rom[25475] = 12'h  0;
rom[25476] = 12'h  0;
rom[25477] = 12'h  0;
rom[25478] = 12'h  0;
rom[25479] = 12'h  0;
rom[25480] = 12'h  0;
rom[25481] = 12'h  0;
rom[25482] = 12'h  0;
rom[25483] = 12'h  0;
rom[25484] = 12'h  0;
rom[25485] = 12'h  0;
rom[25486] = 12'h  0;
rom[25487] = 12'h  0;
rom[25488] = 12'h  0;
rom[25489] = 12'h  0;
rom[25490] = 12'h  0;
rom[25491] = 12'h  0;
rom[25492] = 12'h111;
rom[25493] = 12'h111;
rom[25494] = 12'h111;
rom[25495] = 12'h111;
rom[25496] = 12'h111;
rom[25497] = 12'h111;
rom[25498] = 12'h222;
rom[25499] = 12'h222;
rom[25500] = 12'h222;
rom[25501] = 12'h222;
rom[25502] = 12'h222;
rom[25503] = 12'h222;
rom[25504] = 12'h222;
rom[25505] = 12'h344;
rom[25506] = 12'h545;
rom[25507] = 12'h444;
rom[25508] = 12'h444;
rom[25509] = 12'h333;
rom[25510] = 12'h333;
rom[25511] = 12'h444;
rom[25512] = 12'h444;
rom[25513] = 12'h444;
rom[25514] = 12'h444;
rom[25515] = 12'h444;
rom[25516] = 12'h444;
rom[25517] = 12'h455;
rom[25518] = 12'h555;
rom[25519] = 12'h455;
rom[25520] = 12'h555;
rom[25521] = 12'h555;
rom[25522] = 12'h566;
rom[25523] = 12'h666;
rom[25524] = 12'h666;
rom[25525] = 12'h677;
rom[25526] = 12'h777;
rom[25527] = 12'h777;
rom[25528] = 12'h888;
rom[25529] = 12'h898;
rom[25530] = 12'h999;
rom[25531] = 12'haaa;
rom[25532] = 12'hbbb;
rom[25533] = 12'hbbb;
rom[25534] = 12'hccb;
rom[25535] = 12'hccb;
rom[25536] = 12'hbbb;
rom[25537] = 12'hbbb;
rom[25538] = 12'hbbb;
rom[25539] = 12'hbba;
rom[25540] = 12'hbaa;
rom[25541] = 12'hbaa;
rom[25542] = 12'hbaa;
rom[25543] = 12'hba9;
rom[25544] = 12'hba9;
rom[25545] = 12'ha98;
rom[25546] = 12'ha98;
rom[25547] = 12'h987;
rom[25548] = 12'h987;
rom[25549] = 12'h977;
rom[25550] = 12'h876;
rom[25551] = 12'h876;
rom[25552] = 12'h876;
rom[25553] = 12'h776;
rom[25554] = 12'h765;
rom[25555] = 12'h765;
rom[25556] = 12'h765;
rom[25557] = 12'h665;
rom[25558] = 12'h665;
rom[25559] = 12'h665;
rom[25560] = 12'h765;
rom[25561] = 12'h765;
rom[25562] = 12'h765;
rom[25563] = 12'h766;
rom[25564] = 12'h776;
rom[25565] = 12'h776;
rom[25566] = 12'h776;
rom[25567] = 12'h777;
rom[25568] = 12'h776;
rom[25569] = 12'h777;
rom[25570] = 12'h777;
rom[25571] = 12'h777;
rom[25572] = 12'h787;
rom[25573] = 12'h887;
rom[25574] = 12'h777;
rom[25575] = 12'h777;
rom[25576] = 12'h888;
rom[25577] = 12'h888;
rom[25578] = 12'h888;
rom[25579] = 12'h888;
rom[25580] = 12'h888;
rom[25581] = 12'h888;
rom[25582] = 12'h888;
rom[25583] = 12'h889;
rom[25584] = 12'h888;
rom[25585] = 12'h888;
rom[25586] = 12'h888;
rom[25587] = 12'h888;
rom[25588] = 12'h888;
rom[25589] = 12'h888;
rom[25590] = 12'h888;
rom[25591] = 12'h888;
rom[25592] = 12'h888;
rom[25593] = 12'h888;
rom[25594] = 12'h999;
rom[25595] = 12'h999;
rom[25596] = 12'haaa;
rom[25597] = 12'haaa;
rom[25598] = 12'haaa;
rom[25599] = 12'haaa;
rom[25600] = 12'h666;
rom[25601] = 12'h666;
rom[25602] = 12'h666;
rom[25603] = 12'h666;
rom[25604] = 12'h666;
rom[25605] = 12'h666;
rom[25606] = 12'h666;
rom[25607] = 12'h666;
rom[25608] = 12'h666;
rom[25609] = 12'h666;
rom[25610] = 12'h666;
rom[25611] = 12'h666;
rom[25612] = 12'h666;
rom[25613] = 12'h666;
rom[25614] = 12'h666;
rom[25615] = 12'h666;
rom[25616] = 12'h777;
rom[25617] = 12'h777;
rom[25618] = 12'h777;
rom[25619] = 12'h777;
rom[25620] = 12'h777;
rom[25621] = 12'h777;
rom[25622] = 12'h777;
rom[25623] = 12'h777;
rom[25624] = 12'h777;
rom[25625] = 12'h777;
rom[25626] = 12'h777;
rom[25627] = 12'h777;
rom[25628] = 12'h777;
rom[25629] = 12'h777;
rom[25630] = 12'h777;
rom[25631] = 12'h777;
rom[25632] = 12'h777;
rom[25633] = 12'h777;
rom[25634] = 12'h777;
rom[25635] = 12'h777;
rom[25636] = 12'h777;
rom[25637] = 12'h777;
rom[25638] = 12'h777;
rom[25639] = 12'h888;
rom[25640] = 12'h888;
rom[25641] = 12'h888;
rom[25642] = 12'h777;
rom[25643] = 12'h777;
rom[25644] = 12'h777;
rom[25645] = 12'h777;
rom[25646] = 12'h777;
rom[25647] = 12'h777;
rom[25648] = 12'h777;
rom[25649] = 12'h888;
rom[25650] = 12'h888;
rom[25651] = 12'h888;
rom[25652] = 12'h888;
rom[25653] = 12'h888;
rom[25654] = 12'h777;
rom[25655] = 12'h777;
rom[25656] = 12'h777;
rom[25657] = 12'h777;
rom[25658] = 12'h666;
rom[25659] = 12'h666;
rom[25660] = 12'h666;
rom[25661] = 12'h666;
rom[25662] = 12'h555;
rom[25663] = 12'h555;
rom[25664] = 12'h666;
rom[25665] = 12'h555;
rom[25666] = 12'h555;
rom[25667] = 12'h555;
rom[25668] = 12'h555;
rom[25669] = 12'h555;
rom[25670] = 12'h555;
rom[25671] = 12'h555;
rom[25672] = 12'h555;
rom[25673] = 12'h555;
rom[25674] = 12'h555;
rom[25675] = 12'h555;
rom[25676] = 12'h555;
rom[25677] = 12'h444;
rom[25678] = 12'h444;
rom[25679] = 12'h444;
rom[25680] = 12'h444;
rom[25681] = 12'h444;
rom[25682] = 12'h444;
rom[25683] = 12'h444;
rom[25684] = 12'h333;
rom[25685] = 12'h333;
rom[25686] = 12'h444;
rom[25687] = 12'h444;
rom[25688] = 12'h444;
rom[25689] = 12'h444;
rom[25690] = 12'h333;
rom[25691] = 12'h333;
rom[25692] = 12'h333;
rom[25693] = 12'h333;
rom[25694] = 12'h222;
rom[25695] = 12'h222;
rom[25696] = 12'h222;
rom[25697] = 12'h222;
rom[25698] = 12'h111;
rom[25699] = 12'h111;
rom[25700] = 12'h111;
rom[25701] = 12'h111;
rom[25702] = 12'h  0;
rom[25703] = 12'h  0;
rom[25704] = 12'h  0;
rom[25705] = 12'h  0;
rom[25706] = 12'h  0;
rom[25707] = 12'h  0;
rom[25708] = 12'h  0;
rom[25709] = 12'h  0;
rom[25710] = 12'h  0;
rom[25711] = 12'h  0;
rom[25712] = 12'h  0;
rom[25713] = 12'h  0;
rom[25714] = 12'h  0;
rom[25715] = 12'h  0;
rom[25716] = 12'h100;
rom[25717] = 12'h100;
rom[25718] = 12'h100;
rom[25719] = 12'h200;
rom[25720] = 12'h200;
rom[25721] = 12'h300;
rom[25722] = 12'h300;
rom[25723] = 12'h400;
rom[25724] = 12'h510;
rom[25725] = 12'h610;
rom[25726] = 12'h720;
rom[25727] = 12'h820;
rom[25728] = 12'ha40;
rom[25729] = 12'hb50;
rom[25730] = 12'hc60;
rom[25731] = 12'hd71;
rom[25732] = 12'he71;
rom[25733] = 12'hf81;
rom[25734] = 12'hf81;
rom[25735] = 12'hf81;
rom[25736] = 12'hf81;
rom[25737] = 12'hf80;
rom[25738] = 12'hf80;
rom[25739] = 12'hf80;
rom[25740] = 12'hf81;
rom[25741] = 12'hf81;
rom[25742] = 12'hf81;
rom[25743] = 12'hf81;
rom[25744] = 12'he72;
rom[25745] = 12'hd72;
rom[25746] = 12'hd61;
rom[25747] = 12'hc60;
rom[25748] = 12'hc50;
rom[25749] = 12'hb40;
rom[25750] = 12'hb40;
rom[25751] = 12'ha30;
rom[25752] = 12'hb30;
rom[25753] = 12'ha30;
rom[25754] = 12'ha30;
rom[25755] = 12'ha20;
rom[25756] = 12'ha20;
rom[25757] = 12'ha20;
rom[25758] = 12'ha20;
rom[25759] = 12'ha20;
rom[25760] = 12'ha20;
rom[25761] = 12'ha20;
rom[25762] = 12'ha20;
rom[25763] = 12'ha20;
rom[25764] = 12'ha20;
rom[25765] = 12'ha20;
rom[25766] = 12'ha20;
rom[25767] = 12'h920;
rom[25768] = 12'h820;
rom[25769] = 12'h810;
rom[25770] = 12'h710;
rom[25771] = 12'h710;
rom[25772] = 12'h610;
rom[25773] = 12'h600;
rom[25774] = 12'h500;
rom[25775] = 12'h400;
rom[25776] = 12'h400;
rom[25777] = 12'h300;
rom[25778] = 12'h300;
rom[25779] = 12'h300;
rom[25780] = 12'h300;
rom[25781] = 12'h200;
rom[25782] = 12'h200;
rom[25783] = 12'h200;
rom[25784] = 12'h100;
rom[25785] = 12'h200;
rom[25786] = 12'h100;
rom[25787] = 12'h  0;
rom[25788] = 12'h100;
rom[25789] = 12'h222;
rom[25790] = 12'h323;
rom[25791] = 12'h222;
rom[25792] = 12'h112;
rom[25793] = 12'h111;
rom[25794] = 12'h122;
rom[25795] = 12'h222;
rom[25796] = 12'h222;
rom[25797] = 12'h222;
rom[25798] = 12'h222;
rom[25799] = 12'h222;
rom[25800] = 12'h333;
rom[25801] = 12'h333;
rom[25802] = 12'h333;
rom[25803] = 12'h444;
rom[25804] = 12'h666;
rom[25805] = 12'h888;
rom[25806] = 12'h999;
rom[25807] = 12'h999;
rom[25808] = 12'h888;
rom[25809] = 12'h999;
rom[25810] = 12'h999;
rom[25811] = 12'h999;
rom[25812] = 12'h999;
rom[25813] = 12'h999;
rom[25814] = 12'h888;
rom[25815] = 12'h888;
rom[25816] = 12'h888;
rom[25817] = 12'h888;
rom[25818] = 12'h888;
rom[25819] = 12'h888;
rom[25820] = 12'h888;
rom[25821] = 12'h888;
rom[25822] = 12'h888;
rom[25823] = 12'h888;
rom[25824] = 12'h888;
rom[25825] = 12'h888;
rom[25826] = 12'h888;
rom[25827] = 12'h888;
rom[25828] = 12'h888;
rom[25829] = 12'h888;
rom[25830] = 12'h777;
rom[25831] = 12'h777;
rom[25832] = 12'h777;
rom[25833] = 12'h777;
rom[25834] = 12'h666;
rom[25835] = 12'h666;
rom[25836] = 12'h666;
rom[25837] = 12'h555;
rom[25838] = 12'h555;
rom[25839] = 12'h555;
rom[25840] = 12'h444;
rom[25841] = 12'h444;
rom[25842] = 12'h444;
rom[25843] = 12'h333;
rom[25844] = 12'h333;
rom[25845] = 12'h222;
rom[25846] = 12'h222;
rom[25847] = 12'h222;
rom[25848] = 12'h222;
rom[25849] = 12'h222;
rom[25850] = 12'h222;
rom[25851] = 12'h222;
rom[25852] = 12'h222;
rom[25853] = 12'h222;
rom[25854] = 12'h111;
rom[25855] = 12'h  0;
rom[25856] = 12'h111;
rom[25857] = 12'h  0;
rom[25858] = 12'h  0;
rom[25859] = 12'h  0;
rom[25860] = 12'h  0;
rom[25861] = 12'h  0;
rom[25862] = 12'h  0;
rom[25863] = 12'h  0;
rom[25864] = 12'h  0;
rom[25865] = 12'h  0;
rom[25866] = 12'h  0;
rom[25867] = 12'h  0;
rom[25868] = 12'h  0;
rom[25869] = 12'h  0;
rom[25870] = 12'h  0;
rom[25871] = 12'h  0;
rom[25872] = 12'h  0;
rom[25873] = 12'h  0;
rom[25874] = 12'h  0;
rom[25875] = 12'h  0;
rom[25876] = 12'h  0;
rom[25877] = 12'h  0;
rom[25878] = 12'h  0;
rom[25879] = 12'h  0;
rom[25880] = 12'h  0;
rom[25881] = 12'h  0;
rom[25882] = 12'h  0;
rom[25883] = 12'h  0;
rom[25884] = 12'h  0;
rom[25885] = 12'h  0;
rom[25886] = 12'h  0;
rom[25887] = 12'h  0;
rom[25888] = 12'h  0;
rom[25889] = 12'h  0;
rom[25890] = 12'h  0;
rom[25891] = 12'h  0;
rom[25892] = 12'h111;
rom[25893] = 12'h111;
rom[25894] = 12'h111;
rom[25895] = 12'h111;
rom[25896] = 12'h111;
rom[25897] = 12'h222;
rom[25898] = 12'h222;
rom[25899] = 12'h222;
rom[25900] = 12'h222;
rom[25901] = 12'h222;
rom[25902] = 12'h222;
rom[25903] = 12'h222;
rom[25904] = 12'h233;
rom[25905] = 12'h334;
rom[25906] = 12'h444;
rom[25907] = 12'h444;
rom[25908] = 12'h344;
rom[25909] = 12'h344;
rom[25910] = 12'h444;
rom[25911] = 12'h444;
rom[25912] = 12'h444;
rom[25913] = 12'h444;
rom[25914] = 12'h445;
rom[25915] = 12'h455;
rom[25916] = 12'h555;
rom[25917] = 12'h555;
rom[25918] = 12'h666;
rom[25919] = 12'h666;
rom[25920] = 12'h677;
rom[25921] = 12'h666;
rom[25922] = 12'h566;
rom[25923] = 12'h667;
rom[25924] = 12'h777;
rom[25925] = 12'h788;
rom[25926] = 12'h888;
rom[25927] = 12'h888;
rom[25928] = 12'h999;
rom[25929] = 12'haaa;
rom[25930] = 12'hbbb;
rom[25931] = 12'hccc;
rom[25932] = 12'hccc;
rom[25933] = 12'hccc;
rom[25934] = 12'hdcc;
rom[25935] = 12'hdcc;
rom[25936] = 12'hddc;
rom[25937] = 12'hdcb;
rom[25938] = 12'hccb;
rom[25939] = 12'hdcb;
rom[25940] = 12'hdcb;
rom[25941] = 12'hcba;
rom[25942] = 12'hba8;
rom[25943] = 12'hb97;
rom[25944] = 12'ha86;
rom[25945] = 12'ha75;
rom[25946] = 12'h964;
rom[25947] = 12'h964;
rom[25948] = 12'h864;
rom[25949] = 12'h853;
rom[25950] = 12'h853;
rom[25951] = 12'h742;
rom[25952] = 12'h742;
rom[25953] = 12'h742;
rom[25954] = 12'h752;
rom[25955] = 12'h652;
rom[25956] = 12'h642;
rom[25957] = 12'h642;
rom[25958] = 12'h652;
rom[25959] = 12'h653;
rom[25960] = 12'h653;
rom[25961] = 12'h753;
rom[25962] = 12'h754;
rom[25963] = 12'h754;
rom[25964] = 12'h754;
rom[25965] = 12'h665;
rom[25966] = 12'h765;
rom[25967] = 12'h766;
rom[25968] = 12'h776;
rom[25969] = 12'h776;
rom[25970] = 12'h777;
rom[25971] = 12'h877;
rom[25972] = 12'h777;
rom[25973] = 12'h777;
rom[25974] = 12'h888;
rom[25975] = 12'h888;
rom[25976] = 12'h888;
rom[25977] = 12'h888;
rom[25978] = 12'h888;
rom[25979] = 12'h888;
rom[25980] = 12'h888;
rom[25981] = 12'h888;
rom[25982] = 12'h888;
rom[25983] = 12'h889;
rom[25984] = 12'h999;
rom[25985] = 12'h999;
rom[25986] = 12'h888;
rom[25987] = 12'h888;
rom[25988] = 12'h888;
rom[25989] = 12'h888;
rom[25990] = 12'h888;
rom[25991] = 12'h888;
rom[25992] = 12'h888;
rom[25993] = 12'h999;
rom[25994] = 12'h999;
rom[25995] = 12'h999;
rom[25996] = 12'haaa;
rom[25997] = 12'haaa;
rom[25998] = 12'haaa;
rom[25999] = 12'haaa;
rom[26000] = 12'h555;
rom[26001] = 12'h555;
rom[26002] = 12'h555;
rom[26003] = 12'h555;
rom[26004] = 12'h555;
rom[26005] = 12'h666;
rom[26006] = 12'h666;
rom[26007] = 12'h666;
rom[26008] = 12'h666;
rom[26009] = 12'h666;
rom[26010] = 12'h666;
rom[26011] = 12'h666;
rom[26012] = 12'h666;
rom[26013] = 12'h666;
rom[26014] = 12'h666;
rom[26015] = 12'h666;
rom[26016] = 12'h666;
rom[26017] = 12'h666;
rom[26018] = 12'h666;
rom[26019] = 12'h666;
rom[26020] = 12'h666;
rom[26021] = 12'h777;
rom[26022] = 12'h777;
rom[26023] = 12'h777;
rom[26024] = 12'h777;
rom[26025] = 12'h777;
rom[26026] = 12'h777;
rom[26027] = 12'h777;
rom[26028] = 12'h777;
rom[26029] = 12'h777;
rom[26030] = 12'h777;
rom[26031] = 12'h777;
rom[26032] = 12'h777;
rom[26033] = 12'h777;
rom[26034] = 12'h777;
rom[26035] = 12'h777;
rom[26036] = 12'h777;
rom[26037] = 12'h777;
rom[26038] = 12'h777;
rom[26039] = 12'h888;
rom[26040] = 12'h888;
rom[26041] = 12'h888;
rom[26042] = 12'h888;
rom[26043] = 12'h777;
rom[26044] = 12'h777;
rom[26045] = 12'h777;
rom[26046] = 12'h777;
rom[26047] = 12'h777;
rom[26048] = 12'h777;
rom[26049] = 12'h888;
rom[26050] = 12'h888;
rom[26051] = 12'h888;
rom[26052] = 12'h888;
rom[26053] = 12'h888;
rom[26054] = 12'h888;
rom[26055] = 12'h777;
rom[26056] = 12'h777;
rom[26057] = 12'h777;
rom[26058] = 12'h777;
rom[26059] = 12'h666;
rom[26060] = 12'h666;
rom[26061] = 12'h666;
rom[26062] = 12'h666;
rom[26063] = 12'h666;
rom[26064] = 12'h666;
rom[26065] = 12'h555;
rom[26066] = 12'h555;
rom[26067] = 12'h555;
rom[26068] = 12'h555;
rom[26069] = 12'h555;
rom[26070] = 12'h555;
rom[26071] = 12'h555;
rom[26072] = 12'h555;
rom[26073] = 12'h555;
rom[26074] = 12'h555;
rom[26075] = 12'h555;
rom[26076] = 12'h444;
rom[26077] = 12'h444;
rom[26078] = 12'h444;
rom[26079] = 12'h444;
rom[26080] = 12'h444;
rom[26081] = 12'h444;
rom[26082] = 12'h444;
rom[26083] = 12'h333;
rom[26084] = 12'h333;
rom[26085] = 12'h333;
rom[26086] = 12'h444;
rom[26087] = 12'h444;
rom[26088] = 12'h444;
rom[26089] = 12'h333;
rom[26090] = 12'h333;
rom[26091] = 12'h333;
rom[26092] = 12'h333;
rom[26093] = 12'h333;
rom[26094] = 12'h222;
rom[26095] = 12'h222;
rom[26096] = 12'h111;
rom[26097] = 12'h111;
rom[26098] = 12'h111;
rom[26099] = 12'h111;
rom[26100] = 12'h111;
rom[26101] = 12'h111;
rom[26102] = 12'h  0;
rom[26103] = 12'h  0;
rom[26104] = 12'h  0;
rom[26105] = 12'h  0;
rom[26106] = 12'h  0;
rom[26107] = 12'h  0;
rom[26108] = 12'h  0;
rom[26109] = 12'h  0;
rom[26110] = 12'h  0;
rom[26111] = 12'h  0;
rom[26112] = 12'h  0;
rom[26113] = 12'h  0;
rom[26114] = 12'h  0;
rom[26115] = 12'h  0;
rom[26116] = 12'h  0;
rom[26117] = 12'h100;
rom[26118] = 12'h100;
rom[26119] = 12'h200;
rom[26120] = 12'h200;
rom[26121] = 12'h300;
rom[26122] = 12'h300;
rom[26123] = 12'h400;
rom[26124] = 12'h510;
rom[26125] = 12'h510;
rom[26126] = 12'h611;
rom[26127] = 12'h720;
rom[26128] = 12'h930;
rom[26129] = 12'ha40;
rom[26130] = 12'hb50;
rom[26131] = 12'hc61;
rom[26132] = 12'hd71;
rom[26133] = 12'he71;
rom[26134] = 12'hf81;
rom[26135] = 12'hf81;
rom[26136] = 12'hf80;
rom[26137] = 12'hf80;
rom[26138] = 12'hf80;
rom[26139] = 12'hf80;
rom[26140] = 12'hf80;
rom[26141] = 12'hf80;
rom[26142] = 12'hf80;
rom[26143] = 12'hf80;
rom[26144] = 12'hf81;
rom[26145] = 12'hf71;
rom[26146] = 12'he71;
rom[26147] = 12'he71;
rom[26148] = 12'he60;
rom[26149] = 12'he60;
rom[26150] = 12'he50;
rom[26151] = 12'hd50;
rom[26152] = 12'hd50;
rom[26153] = 12'hd40;
rom[26154] = 12'hc40;
rom[26155] = 12'hc40;
rom[26156] = 12'hc30;
rom[26157] = 12'hc30;
rom[26158] = 12'hc30;
rom[26159] = 12'hb30;
rom[26160] = 12'hb30;
rom[26161] = 12'hb30;
rom[26162] = 12'hb30;
rom[26163] = 12'hb30;
rom[26164] = 12'ha30;
rom[26165] = 12'ha20;
rom[26166] = 12'h920;
rom[26167] = 12'h920;
rom[26168] = 12'h810;
rom[26169] = 12'h710;
rom[26170] = 12'h710;
rom[26171] = 12'h610;
rom[26172] = 12'h600;
rom[26173] = 12'h500;
rom[26174] = 12'h500;
rom[26175] = 12'h400;
rom[26176] = 12'h400;
rom[26177] = 12'h300;
rom[26178] = 12'h300;
rom[26179] = 12'h300;
rom[26180] = 12'h300;
rom[26181] = 12'h200;
rom[26182] = 12'h200;
rom[26183] = 12'h200;
rom[26184] = 12'h200;
rom[26185] = 12'h100;
rom[26186] = 12'h100;
rom[26187] = 12'h100;
rom[26188] = 12'h111;
rom[26189] = 12'h222;
rom[26190] = 12'h323;
rom[26191] = 12'h212;
rom[26192] = 12'h211;
rom[26193] = 12'h111;
rom[26194] = 12'h111;
rom[26195] = 12'h222;
rom[26196] = 12'h222;
rom[26197] = 12'h222;
rom[26198] = 12'h222;
rom[26199] = 12'h222;
rom[26200] = 12'h333;
rom[26201] = 12'h333;
rom[26202] = 12'h333;
rom[26203] = 12'h444;
rom[26204] = 12'h666;
rom[26205] = 12'h777;
rom[26206] = 12'h999;
rom[26207] = 12'h999;
rom[26208] = 12'h888;
rom[26209] = 12'h888;
rom[26210] = 12'h999;
rom[26211] = 12'h999;
rom[26212] = 12'h999;
rom[26213] = 12'h888;
rom[26214] = 12'h888;
rom[26215] = 12'h888;
rom[26216] = 12'h888;
rom[26217] = 12'h888;
rom[26218] = 12'h888;
rom[26219] = 12'h888;
rom[26220] = 12'h888;
rom[26221] = 12'h888;
rom[26222] = 12'h888;
rom[26223] = 12'h888;
rom[26224] = 12'h888;
rom[26225] = 12'h888;
rom[26226] = 12'h888;
rom[26227] = 12'h777;
rom[26228] = 12'h888;
rom[26229] = 12'h888;
rom[26230] = 12'h777;
rom[26231] = 12'h777;
rom[26232] = 12'h777;
rom[26233] = 12'h777;
rom[26234] = 12'h666;
rom[26235] = 12'h666;
rom[26236] = 12'h666;
rom[26237] = 12'h555;
rom[26238] = 12'h555;
rom[26239] = 12'h555;
rom[26240] = 12'h444;
rom[26241] = 12'h444;
rom[26242] = 12'h333;
rom[26243] = 12'h333;
rom[26244] = 12'h333;
rom[26245] = 12'h222;
rom[26246] = 12'h222;
rom[26247] = 12'h222;
rom[26248] = 12'h222;
rom[26249] = 12'h222;
rom[26250] = 12'h222;
rom[26251] = 12'h222;
rom[26252] = 12'h222;
rom[26253] = 12'h222;
rom[26254] = 12'h111;
rom[26255] = 12'h  0;
rom[26256] = 12'h  0;
rom[26257] = 12'h  0;
rom[26258] = 12'h  0;
rom[26259] = 12'h  0;
rom[26260] = 12'h  0;
rom[26261] = 12'h  0;
rom[26262] = 12'h  0;
rom[26263] = 12'h  0;
rom[26264] = 12'h  0;
rom[26265] = 12'h  0;
rom[26266] = 12'h  0;
rom[26267] = 12'h  0;
rom[26268] = 12'h  0;
rom[26269] = 12'h  0;
rom[26270] = 12'h  0;
rom[26271] = 12'h  0;
rom[26272] = 12'h  0;
rom[26273] = 12'h  0;
rom[26274] = 12'h  0;
rom[26275] = 12'h  0;
rom[26276] = 12'h  0;
rom[26277] = 12'h  0;
rom[26278] = 12'h  0;
rom[26279] = 12'h  0;
rom[26280] = 12'h  0;
rom[26281] = 12'h  0;
rom[26282] = 12'h  0;
rom[26283] = 12'h  0;
rom[26284] = 12'h  0;
rom[26285] = 12'h  0;
rom[26286] = 12'h  0;
rom[26287] = 12'h  0;
rom[26288] = 12'h  0;
rom[26289] = 12'h  0;
rom[26290] = 12'h  0;
rom[26291] = 12'h111;
rom[26292] = 12'h111;
rom[26293] = 12'h111;
rom[26294] = 12'h111;
rom[26295] = 12'h111;
rom[26296] = 12'h222;
rom[26297] = 12'h222;
rom[26298] = 12'h222;
rom[26299] = 12'h222;
rom[26300] = 12'h222;
rom[26301] = 12'h222;
rom[26302] = 12'h222;
rom[26303] = 12'h222;
rom[26304] = 12'h333;
rom[26305] = 12'h344;
rom[26306] = 12'h445;
rom[26307] = 12'h444;
rom[26308] = 12'h444;
rom[26309] = 12'h444;
rom[26310] = 12'h444;
rom[26311] = 12'h444;
rom[26312] = 12'h455;
rom[26313] = 12'h555;
rom[26314] = 12'h555;
rom[26315] = 12'h555;
rom[26316] = 12'h555;
rom[26317] = 12'h556;
rom[26318] = 12'h666;
rom[26319] = 12'h666;
rom[26320] = 12'h667;
rom[26321] = 12'h677;
rom[26322] = 12'h778;
rom[26323] = 12'h778;
rom[26324] = 12'h788;
rom[26325] = 12'h788;
rom[26326] = 12'h899;
rom[26327] = 12'haaa;
rom[26328] = 12'haba;
rom[26329] = 12'hbbb;
rom[26330] = 12'hccc;
rom[26331] = 12'hddc;
rom[26332] = 12'hddc;
rom[26333] = 12'hddc;
rom[26334] = 12'hedc;
rom[26335] = 12'heed;
rom[26336] = 12'hddc;
rom[26337] = 12'hccb;
rom[26338] = 12'hba9;
rom[26339] = 12'ha98;
rom[26340] = 12'ha87;
rom[26341] = 12'h976;
rom[26342] = 12'h965;
rom[26343] = 12'h964;
rom[26344] = 12'h852;
rom[26345] = 12'h842;
rom[26346] = 12'h841;
rom[26347] = 12'h841;
rom[26348] = 12'h841;
rom[26349] = 12'h841;
rom[26350] = 12'h741;
rom[26351] = 12'h731;
rom[26352] = 12'h741;
rom[26353] = 12'h741;
rom[26354] = 12'h741;
rom[26355] = 12'h641;
rom[26356] = 12'h641;
rom[26357] = 12'h641;
rom[26358] = 12'h641;
rom[26359] = 12'h642;
rom[26360] = 12'h752;
rom[26361] = 12'h752;
rom[26362] = 12'h753;
rom[26363] = 12'h653;
rom[26364] = 12'h643;
rom[26365] = 12'h654;
rom[26366] = 12'h654;
rom[26367] = 12'h665;
rom[26368] = 12'h665;
rom[26369] = 12'h765;
rom[26370] = 12'h776;
rom[26371] = 12'h776;
rom[26372] = 12'h777;
rom[26373] = 12'h777;
rom[26374] = 12'h777;
rom[26375] = 12'h788;
rom[26376] = 12'h888;
rom[26377] = 12'h888;
rom[26378] = 12'h888;
rom[26379] = 12'h888;
rom[26380] = 12'h888;
rom[26381] = 12'h888;
rom[26382] = 12'h888;
rom[26383] = 12'h888;
rom[26384] = 12'h999;
rom[26385] = 12'h999;
rom[26386] = 12'h888;
rom[26387] = 12'h888;
rom[26388] = 12'h888;
rom[26389] = 12'h888;
rom[26390] = 12'h888;
rom[26391] = 12'h888;
rom[26392] = 12'h888;
rom[26393] = 12'h999;
rom[26394] = 12'h999;
rom[26395] = 12'h999;
rom[26396] = 12'haaa;
rom[26397] = 12'haaa;
rom[26398] = 12'haaa;
rom[26399] = 12'haaa;
rom[26400] = 12'h555;
rom[26401] = 12'h555;
rom[26402] = 12'h555;
rom[26403] = 12'h555;
rom[26404] = 12'h555;
rom[26405] = 12'h555;
rom[26406] = 12'h555;
rom[26407] = 12'h555;
rom[26408] = 12'h555;
rom[26409] = 12'h666;
rom[26410] = 12'h666;
rom[26411] = 12'h666;
rom[26412] = 12'h666;
rom[26413] = 12'h666;
rom[26414] = 12'h666;
rom[26415] = 12'h666;
rom[26416] = 12'h666;
rom[26417] = 12'h666;
rom[26418] = 12'h666;
rom[26419] = 12'h666;
rom[26420] = 12'h666;
rom[26421] = 12'h666;
rom[26422] = 12'h666;
rom[26423] = 12'h666;
rom[26424] = 12'h777;
rom[26425] = 12'h777;
rom[26426] = 12'h777;
rom[26427] = 12'h777;
rom[26428] = 12'h777;
rom[26429] = 12'h777;
rom[26430] = 12'h777;
rom[26431] = 12'h777;
rom[26432] = 12'h777;
rom[26433] = 12'h777;
rom[26434] = 12'h777;
rom[26435] = 12'h777;
rom[26436] = 12'h777;
rom[26437] = 12'h777;
rom[26438] = 12'h888;
rom[26439] = 12'h888;
rom[26440] = 12'h888;
rom[26441] = 12'h888;
rom[26442] = 12'h888;
rom[26443] = 12'h777;
rom[26444] = 12'h777;
rom[26445] = 12'h777;
rom[26446] = 12'h777;
rom[26447] = 12'h777;
rom[26448] = 12'h777;
rom[26449] = 12'h888;
rom[26450] = 12'h888;
rom[26451] = 12'h888;
rom[26452] = 12'h888;
rom[26453] = 12'h888;
rom[26454] = 12'h888;
rom[26455] = 12'h888;
rom[26456] = 12'h777;
rom[26457] = 12'h777;
rom[26458] = 12'h777;
rom[26459] = 12'h666;
rom[26460] = 12'h666;
rom[26461] = 12'h666;
rom[26462] = 12'h666;
rom[26463] = 12'h666;
rom[26464] = 12'h555;
rom[26465] = 12'h555;
rom[26466] = 12'h555;
rom[26467] = 12'h555;
rom[26468] = 12'h555;
rom[26469] = 12'h555;
rom[26470] = 12'h555;
rom[26471] = 12'h555;
rom[26472] = 12'h555;
rom[26473] = 12'h555;
rom[26474] = 12'h555;
rom[26475] = 12'h444;
rom[26476] = 12'h444;
rom[26477] = 12'h444;
rom[26478] = 12'h444;
rom[26479] = 12'h444;
rom[26480] = 12'h444;
rom[26481] = 12'h444;
rom[26482] = 12'h333;
rom[26483] = 12'h333;
rom[26484] = 12'h333;
rom[26485] = 12'h333;
rom[26486] = 12'h333;
rom[26487] = 12'h444;
rom[26488] = 12'h444;
rom[26489] = 12'h333;
rom[26490] = 12'h222;
rom[26491] = 12'h222;
rom[26492] = 12'h222;
rom[26493] = 12'h222;
rom[26494] = 12'h222;
rom[26495] = 12'h222;
rom[26496] = 12'h111;
rom[26497] = 12'h111;
rom[26498] = 12'h111;
rom[26499] = 12'h111;
rom[26500] = 12'h111;
rom[26501] = 12'h  0;
rom[26502] = 12'h  0;
rom[26503] = 12'h  0;
rom[26504] = 12'h  0;
rom[26505] = 12'h  0;
rom[26506] = 12'h  0;
rom[26507] = 12'h  0;
rom[26508] = 12'h  0;
rom[26509] = 12'h  0;
rom[26510] = 12'h  0;
rom[26511] = 12'h  0;
rom[26512] = 12'h  0;
rom[26513] = 12'h  0;
rom[26514] = 12'h  0;
rom[26515] = 12'h  0;
rom[26516] = 12'h  0;
rom[26517] = 12'h100;
rom[26518] = 12'h100;
rom[26519] = 12'h100;
rom[26520] = 12'h200;
rom[26521] = 12'h200;
rom[26522] = 12'h300;
rom[26523] = 12'h300;
rom[26524] = 12'h400;
rom[26525] = 12'h510;
rom[26526] = 12'h510;
rom[26527] = 12'h610;
rom[26528] = 12'h820;
rom[26529] = 12'h930;
rom[26530] = 12'ha40;
rom[26531] = 12'hb50;
rom[26532] = 12'hc60;
rom[26533] = 12'hd60;
rom[26534] = 12'he70;
rom[26535] = 12'he70;
rom[26536] = 12'hf80;
rom[26537] = 12'hf80;
rom[26538] = 12'hf80;
rom[26539] = 12'hf80;
rom[26540] = 12'hf80;
rom[26541] = 12'hf80;
rom[26542] = 12'hf80;
rom[26543] = 12'hf70;
rom[26544] = 12'hf81;
rom[26545] = 12'hf71;
rom[26546] = 12'hf71;
rom[26547] = 12'hf71;
rom[26548] = 12'hf71;
rom[26549] = 12'hf71;
rom[26550] = 12'hf61;
rom[26551] = 12'hf61;
rom[26552] = 12'he51;
rom[26553] = 12'he51;
rom[26554] = 12'he51;
rom[26555] = 12'hd51;
rom[26556] = 12'hd41;
rom[26557] = 12'hd41;
rom[26558] = 12'hd41;
rom[26559] = 12'hc41;
rom[26560] = 12'hc31;
rom[26561] = 12'hc30;
rom[26562] = 12'hb30;
rom[26563] = 12'hb30;
rom[26564] = 12'ha30;
rom[26565] = 12'ha20;
rom[26566] = 12'h920;
rom[26567] = 12'h820;
rom[26568] = 12'h810;
rom[26569] = 12'h710;
rom[26570] = 12'h610;
rom[26571] = 12'h610;
rom[26572] = 12'h500;
rom[26573] = 12'h500;
rom[26574] = 12'h500;
rom[26575] = 12'h400;
rom[26576] = 12'h300;
rom[26577] = 12'h300;
rom[26578] = 12'h300;
rom[26579] = 12'h300;
rom[26580] = 12'h300;
rom[26581] = 12'h200;
rom[26582] = 12'h200;
rom[26583] = 12'h200;
rom[26584] = 12'h200;
rom[26585] = 12'h100;
rom[26586] = 12'h100;
rom[26587] = 12'h101;
rom[26588] = 12'h222;
rom[26589] = 12'h322;
rom[26590] = 12'h222;
rom[26591] = 12'h111;
rom[26592] = 12'h111;
rom[26593] = 12'h111;
rom[26594] = 12'h111;
rom[26595] = 12'h222;
rom[26596] = 12'h222;
rom[26597] = 12'h222;
rom[26598] = 12'h222;
rom[26599] = 12'h222;
rom[26600] = 12'h333;
rom[26601] = 12'h333;
rom[26602] = 12'h333;
rom[26603] = 12'h444;
rom[26604] = 12'h555;
rom[26605] = 12'h777;
rom[26606] = 12'h888;
rom[26607] = 12'h999;
rom[26608] = 12'h888;
rom[26609] = 12'h888;
rom[26610] = 12'h999;
rom[26611] = 12'h999;
rom[26612] = 12'h999;
rom[26613] = 12'h888;
rom[26614] = 12'h888;
rom[26615] = 12'h888;
rom[26616] = 12'h888;
rom[26617] = 12'h888;
rom[26618] = 12'h888;
rom[26619] = 12'h888;
rom[26620] = 12'h888;
rom[26621] = 12'h888;
rom[26622] = 12'h888;
rom[26623] = 12'h888;
rom[26624] = 12'h888;
rom[26625] = 12'h888;
rom[26626] = 12'h777;
rom[26627] = 12'h777;
rom[26628] = 12'h777;
rom[26629] = 12'h777;
rom[26630] = 12'h777;
rom[26631] = 12'h777;
rom[26632] = 12'h777;
rom[26633] = 12'h777;
rom[26634] = 12'h666;
rom[26635] = 12'h666;
rom[26636] = 12'h666;
rom[26637] = 12'h555;
rom[26638] = 12'h555;
rom[26639] = 12'h555;
rom[26640] = 12'h444;
rom[26641] = 12'h444;
rom[26642] = 12'h333;
rom[26643] = 12'h333;
rom[26644] = 12'h333;
rom[26645] = 12'h333;
rom[26646] = 12'h333;
rom[26647] = 12'h333;
rom[26648] = 12'h222;
rom[26649] = 12'h222;
rom[26650] = 12'h222;
rom[26651] = 12'h222;
rom[26652] = 12'h222;
rom[26653] = 12'h111;
rom[26654] = 12'h111;
rom[26655] = 12'h  0;
rom[26656] = 12'h  0;
rom[26657] = 12'h  0;
rom[26658] = 12'h  0;
rom[26659] = 12'h  0;
rom[26660] = 12'h  0;
rom[26661] = 12'h  0;
rom[26662] = 12'h  0;
rom[26663] = 12'h  0;
rom[26664] = 12'h  0;
rom[26665] = 12'h  0;
rom[26666] = 12'h  0;
rom[26667] = 12'h  0;
rom[26668] = 12'h  0;
rom[26669] = 12'h  0;
rom[26670] = 12'h  0;
rom[26671] = 12'h  0;
rom[26672] = 12'h  0;
rom[26673] = 12'h  0;
rom[26674] = 12'h  0;
rom[26675] = 12'h  0;
rom[26676] = 12'h  0;
rom[26677] = 12'h  0;
rom[26678] = 12'h  0;
rom[26679] = 12'h  0;
rom[26680] = 12'h  0;
rom[26681] = 12'h  0;
rom[26682] = 12'h  0;
rom[26683] = 12'h  0;
rom[26684] = 12'h  0;
rom[26685] = 12'h  0;
rom[26686] = 12'h  0;
rom[26687] = 12'h  0;
rom[26688] = 12'h  0;
rom[26689] = 12'h  0;
rom[26690] = 12'h  0;
rom[26691] = 12'h111;
rom[26692] = 12'h111;
rom[26693] = 12'h111;
rom[26694] = 12'h111;
rom[26695] = 12'h111;
rom[26696] = 12'h222;
rom[26697] = 12'h222;
rom[26698] = 12'h222;
rom[26699] = 12'h222;
rom[26700] = 12'h222;
rom[26701] = 12'h222;
rom[26702] = 12'h222;
rom[26703] = 12'h233;
rom[26704] = 12'h334;
rom[26705] = 12'h444;
rom[26706] = 12'h445;
rom[26707] = 12'h445;
rom[26708] = 12'h444;
rom[26709] = 12'h444;
rom[26710] = 12'h445;
rom[26711] = 12'h455;
rom[26712] = 12'h555;
rom[26713] = 12'h555;
rom[26714] = 12'h555;
rom[26715] = 12'h556;
rom[26716] = 12'h556;
rom[26717] = 12'h666;
rom[26718] = 12'h666;
rom[26719] = 12'h667;
rom[26720] = 12'h778;
rom[26721] = 12'h888;
rom[26722] = 12'h899;
rom[26723] = 12'h999;
rom[26724] = 12'h999;
rom[26725] = 12'h9aa;
rom[26726] = 12'hbbb;
rom[26727] = 12'hccc;
rom[26728] = 12'hddc;
rom[26729] = 12'heed;
rom[26730] = 12'heee;
rom[26731] = 12'hfee;
rom[26732] = 12'heed;
rom[26733] = 12'hddc;
rom[26734] = 12'hdcb;
rom[26735] = 12'hcbb;
rom[26736] = 12'hba9;
rom[26737] = 12'ha98;
rom[26738] = 12'h876;
rom[26739] = 12'h754;
rom[26740] = 12'h643;
rom[26741] = 12'h642;
rom[26742] = 12'h631;
rom[26743] = 12'h631;
rom[26744] = 12'h630;
rom[26745] = 12'h620;
rom[26746] = 12'h720;
rom[26747] = 12'h730;
rom[26748] = 12'h730;
rom[26749] = 12'h830;
rom[26750] = 12'h730;
rom[26751] = 12'h730;
rom[26752] = 12'h730;
rom[26753] = 12'h730;
rom[26754] = 12'h730;
rom[26755] = 12'h630;
rom[26756] = 12'h630;
rom[26757] = 12'h630;
rom[26758] = 12'h641;
rom[26759] = 12'h641;
rom[26760] = 12'h742;
rom[26761] = 12'h742;
rom[26762] = 12'h742;
rom[26763] = 12'h642;
rom[26764] = 12'h642;
rom[26765] = 12'h543;
rom[26766] = 12'h543;
rom[26767] = 12'h553;
rom[26768] = 12'h654;
rom[26769] = 12'h654;
rom[26770] = 12'h765;
rom[26771] = 12'h766;
rom[26772] = 12'h776;
rom[26773] = 12'h777;
rom[26774] = 12'h777;
rom[26775] = 12'h777;
rom[26776] = 12'h788;
rom[26777] = 12'h888;
rom[26778] = 12'h888;
rom[26779] = 12'h888;
rom[26780] = 12'h888;
rom[26781] = 12'h888;
rom[26782] = 12'h888;
rom[26783] = 12'h888;
rom[26784] = 12'h889;
rom[26785] = 12'h999;
rom[26786] = 12'h999;
rom[26787] = 12'h999;
rom[26788] = 12'h999;
rom[26789] = 12'h888;
rom[26790] = 12'h888;
rom[26791] = 12'h888;
rom[26792] = 12'h888;
rom[26793] = 12'h999;
rom[26794] = 12'h999;
rom[26795] = 12'h999;
rom[26796] = 12'haaa;
rom[26797] = 12'haaa;
rom[26798] = 12'haaa;
rom[26799] = 12'haaa;
rom[26800] = 12'h555;
rom[26801] = 12'h555;
rom[26802] = 12'h555;
rom[26803] = 12'h555;
rom[26804] = 12'h555;
rom[26805] = 12'h555;
rom[26806] = 12'h555;
rom[26807] = 12'h555;
rom[26808] = 12'h555;
rom[26809] = 12'h555;
rom[26810] = 12'h555;
rom[26811] = 12'h555;
rom[26812] = 12'h666;
rom[26813] = 12'h666;
rom[26814] = 12'h666;
rom[26815] = 12'h666;
rom[26816] = 12'h666;
rom[26817] = 12'h666;
rom[26818] = 12'h666;
rom[26819] = 12'h666;
rom[26820] = 12'h666;
rom[26821] = 12'h666;
rom[26822] = 12'h666;
rom[26823] = 12'h666;
rom[26824] = 12'h666;
rom[26825] = 12'h777;
rom[26826] = 12'h777;
rom[26827] = 12'h777;
rom[26828] = 12'h777;
rom[26829] = 12'h777;
rom[26830] = 12'h777;
rom[26831] = 12'h777;
rom[26832] = 12'h777;
rom[26833] = 12'h777;
rom[26834] = 12'h777;
rom[26835] = 12'h777;
rom[26836] = 12'h777;
rom[26837] = 12'h777;
rom[26838] = 12'h888;
rom[26839] = 12'h888;
rom[26840] = 12'h888;
rom[26841] = 12'h888;
rom[26842] = 12'h888;
rom[26843] = 12'h888;
rom[26844] = 12'h777;
rom[26845] = 12'h777;
rom[26846] = 12'h777;
rom[26847] = 12'h777;
rom[26848] = 12'h777;
rom[26849] = 12'h777;
rom[26850] = 12'h777;
rom[26851] = 12'h777;
rom[26852] = 12'h888;
rom[26853] = 12'h888;
rom[26854] = 12'h888;
rom[26855] = 12'h888;
rom[26856] = 12'h888;
rom[26857] = 12'h888;
rom[26858] = 12'h777;
rom[26859] = 12'h777;
rom[26860] = 12'h666;
rom[26861] = 12'h666;
rom[26862] = 12'h666;
rom[26863] = 12'h666;
rom[26864] = 12'h555;
rom[26865] = 12'h555;
rom[26866] = 12'h555;
rom[26867] = 12'h555;
rom[26868] = 12'h555;
rom[26869] = 12'h555;
rom[26870] = 12'h555;
rom[26871] = 12'h555;
rom[26872] = 12'h555;
rom[26873] = 12'h555;
rom[26874] = 12'h555;
rom[26875] = 12'h444;
rom[26876] = 12'h444;
rom[26877] = 12'h444;
rom[26878] = 12'h444;
rom[26879] = 12'h444;
rom[26880] = 12'h444;
rom[26881] = 12'h333;
rom[26882] = 12'h333;
rom[26883] = 12'h333;
rom[26884] = 12'h333;
rom[26885] = 12'h333;
rom[26886] = 12'h333;
rom[26887] = 12'h333;
rom[26888] = 12'h333;
rom[26889] = 12'h333;
rom[26890] = 12'h222;
rom[26891] = 12'h222;
rom[26892] = 12'h222;
rom[26893] = 12'h222;
rom[26894] = 12'h222;
rom[26895] = 12'h222;
rom[26896] = 12'h111;
rom[26897] = 12'h111;
rom[26898] = 12'h111;
rom[26899] = 12'h  0;
rom[26900] = 12'h  0;
rom[26901] = 12'h  0;
rom[26902] = 12'h  0;
rom[26903] = 12'h  0;
rom[26904] = 12'h  0;
rom[26905] = 12'h  0;
rom[26906] = 12'h  0;
rom[26907] = 12'h  0;
rom[26908] = 12'h  0;
rom[26909] = 12'h  0;
rom[26910] = 12'h  0;
rom[26911] = 12'h  0;
rom[26912] = 12'h  0;
rom[26913] = 12'h  0;
rom[26914] = 12'h  0;
rom[26915] = 12'h  0;
rom[26916] = 12'h  0;
rom[26917] = 12'h  0;
rom[26918] = 12'h100;
rom[26919] = 12'h100;
rom[26920] = 12'h200;
rom[26921] = 12'h200;
rom[26922] = 12'h300;
rom[26923] = 12'h300;
rom[26924] = 12'h400;
rom[26925] = 12'h400;
rom[26926] = 12'h510;
rom[26927] = 12'h510;
rom[26928] = 12'h720;
rom[26929] = 12'h820;
rom[26930] = 12'h830;
rom[26931] = 12'h940;
rom[26932] = 12'ha50;
rom[26933] = 12'hb50;
rom[26934] = 12'hc60;
rom[26935] = 12'hd70;
rom[26936] = 12'he70;
rom[26937] = 12'he70;
rom[26938] = 12'he70;
rom[26939] = 12'he70;
rom[26940] = 12'hf70;
rom[26941] = 12'hf70;
rom[26942] = 12'hf70;
rom[26943] = 12'hf70;
rom[26944] = 12'hf71;
rom[26945] = 12'hf71;
rom[26946] = 12'hf61;
rom[26947] = 12'hf61;
rom[26948] = 12'hf61;
rom[26949] = 12'hf61;
rom[26950] = 12'hf61;
rom[26951] = 12'hf61;
rom[26952] = 12'hf51;
rom[26953] = 12'he51;
rom[26954] = 12'he51;
rom[26955] = 12'he51;
rom[26956] = 12'he51;
rom[26957] = 12'he51;
rom[26958] = 12'hd41;
rom[26959] = 12'hd41;
rom[26960] = 12'hc41;
rom[26961] = 12'hb31;
rom[26962] = 12'hb30;
rom[26963] = 12'ha30;
rom[26964] = 12'ha20;
rom[26965] = 12'h920;
rom[26966] = 12'h820;
rom[26967] = 12'h810;
rom[26968] = 12'h710;
rom[26969] = 12'h610;
rom[26970] = 12'h610;
rom[26971] = 12'h500;
rom[26972] = 12'h500;
rom[26973] = 12'h400;
rom[26974] = 12'h400;
rom[26975] = 12'h400;
rom[26976] = 12'h300;
rom[26977] = 12'h300;
rom[26978] = 12'h300;
rom[26979] = 12'h300;
rom[26980] = 12'h200;
rom[26981] = 12'h200;
rom[26982] = 12'h200;
rom[26983] = 12'h200;
rom[26984] = 12'h100;
rom[26985] = 12'h100;
rom[26986] = 12'h100;
rom[26987] = 12'h211;
rom[26988] = 12'h322;
rom[26989] = 12'h222;
rom[26990] = 12'h212;
rom[26991] = 12'h111;
rom[26992] = 12'h111;
rom[26993] = 12'h111;
rom[26994] = 12'h111;
rom[26995] = 12'h111;
rom[26996] = 12'h222;
rom[26997] = 12'h222;
rom[26998] = 12'h222;
rom[26999] = 12'h222;
rom[27000] = 12'h222;
rom[27001] = 12'h333;
rom[27002] = 12'h333;
rom[27003] = 12'h444;
rom[27004] = 12'h555;
rom[27005] = 12'h777;
rom[27006] = 12'h888;
rom[27007] = 12'h999;
rom[27008] = 12'h888;
rom[27009] = 12'h888;
rom[27010] = 12'h999;
rom[27011] = 12'h999;
rom[27012] = 12'h999;
rom[27013] = 12'h888;
rom[27014] = 12'h888;
rom[27015] = 12'h888;
rom[27016] = 12'h888;
rom[27017] = 12'h888;
rom[27018] = 12'h777;
rom[27019] = 12'h888;
rom[27020] = 12'h888;
rom[27021] = 12'h888;
rom[27022] = 12'h888;
rom[27023] = 12'h777;
rom[27024] = 12'h777;
rom[27025] = 12'h777;
rom[27026] = 12'h777;
rom[27027] = 12'h777;
rom[27028] = 12'h777;
rom[27029] = 12'h777;
rom[27030] = 12'h777;
rom[27031] = 12'h777;
rom[27032] = 12'h777;
rom[27033] = 12'h777;
rom[27034] = 12'h666;
rom[27035] = 12'h666;
rom[27036] = 12'h666;
rom[27037] = 12'h555;
rom[27038] = 12'h555;
rom[27039] = 12'h555;
rom[27040] = 12'h444;
rom[27041] = 12'h444;
rom[27042] = 12'h333;
rom[27043] = 12'h333;
rom[27044] = 12'h333;
rom[27045] = 12'h333;
rom[27046] = 12'h333;
rom[27047] = 12'h333;
rom[27048] = 12'h333;
rom[27049] = 12'h222;
rom[27050] = 12'h222;
rom[27051] = 12'h111;
rom[27052] = 12'h111;
rom[27053] = 12'h111;
rom[27054] = 12'h111;
rom[27055] = 12'h  0;
rom[27056] = 12'h  0;
rom[27057] = 12'h  0;
rom[27058] = 12'h  0;
rom[27059] = 12'h  0;
rom[27060] = 12'h  0;
rom[27061] = 12'h  0;
rom[27062] = 12'h  0;
rom[27063] = 12'h  0;
rom[27064] = 12'h  0;
rom[27065] = 12'h  0;
rom[27066] = 12'h  0;
rom[27067] = 12'h  0;
rom[27068] = 12'h  0;
rom[27069] = 12'h  0;
rom[27070] = 12'h  0;
rom[27071] = 12'h  0;
rom[27072] = 12'h  0;
rom[27073] = 12'h  0;
rom[27074] = 12'h  0;
rom[27075] = 12'h  0;
rom[27076] = 12'h  0;
rom[27077] = 12'h  0;
rom[27078] = 12'h  0;
rom[27079] = 12'h  0;
rom[27080] = 12'h  0;
rom[27081] = 12'h  0;
rom[27082] = 12'h  0;
rom[27083] = 12'h  0;
rom[27084] = 12'h  0;
rom[27085] = 12'h  0;
rom[27086] = 12'h  0;
rom[27087] = 12'h  0;
rom[27088] = 12'h  0;
rom[27089] = 12'h  0;
rom[27090] = 12'h  0;
rom[27091] = 12'h111;
rom[27092] = 12'h111;
rom[27093] = 12'h111;
rom[27094] = 12'h111;
rom[27095] = 12'h111;
rom[27096] = 12'h222;
rom[27097] = 12'h222;
rom[27098] = 12'h222;
rom[27099] = 12'h222;
rom[27100] = 12'h222;
rom[27101] = 12'h222;
rom[27102] = 12'h222;
rom[27103] = 12'h333;
rom[27104] = 12'h444;
rom[27105] = 12'h445;
rom[27106] = 12'h455;
rom[27107] = 12'h445;
rom[27108] = 12'h444;
rom[27109] = 12'h455;
rom[27110] = 12'h555;
rom[27111] = 12'h555;
rom[27112] = 12'h555;
rom[27113] = 12'h555;
rom[27114] = 12'h556;
rom[27115] = 12'h666;
rom[27116] = 12'h666;
rom[27117] = 12'h677;
rom[27118] = 12'h777;
rom[27119] = 12'h888;
rom[27120] = 12'h999;
rom[27121] = 12'h999;
rom[27122] = 12'h999;
rom[27123] = 12'haaa;
rom[27124] = 12'hbbb;
rom[27125] = 12'hccc;
rom[27126] = 12'hddd;
rom[27127] = 12'hddd;
rom[27128] = 12'hfff;
rom[27129] = 12'hffe;
rom[27130] = 12'hffe;
rom[27131] = 12'heed;
rom[27132] = 12'hdcb;
rom[27133] = 12'hba9;
rom[27134] = 12'h977;
rom[27135] = 12'h765;
rom[27136] = 12'h654;
rom[27137] = 12'h543;
rom[27138] = 12'h532;
rom[27139] = 12'h531;
rom[27140] = 12'h521;
rom[27141] = 12'h521;
rom[27142] = 12'h620;
rom[27143] = 12'h620;
rom[27144] = 12'h730;
rom[27145] = 12'h730;
rom[27146] = 12'h730;
rom[27147] = 12'h830;
rom[27148] = 12'h830;
rom[27149] = 12'h931;
rom[27150] = 12'h830;
rom[27151] = 12'h830;
rom[27152] = 12'h830;
rom[27153] = 12'h840;
rom[27154] = 12'h740;
rom[27155] = 12'h730;
rom[27156] = 12'h630;
rom[27157] = 12'h640;
rom[27158] = 12'h741;
rom[27159] = 12'h752;
rom[27160] = 12'h852;
rom[27161] = 12'h752;
rom[27162] = 12'h742;
rom[27163] = 12'h742;
rom[27164] = 12'h642;
rom[27165] = 12'h642;
rom[27166] = 12'h542;
rom[27167] = 12'h542;
rom[27168] = 12'h543;
rom[27169] = 12'h653;
rom[27170] = 12'h654;
rom[27171] = 12'h765;
rom[27172] = 12'h766;
rom[27173] = 12'h776;
rom[27174] = 12'h777;
rom[27175] = 12'h877;
rom[27176] = 12'h888;
rom[27177] = 12'h888;
rom[27178] = 12'h888;
rom[27179] = 12'h888;
rom[27180] = 12'h888;
rom[27181] = 12'h888;
rom[27182] = 12'h888;
rom[27183] = 12'h888;
rom[27184] = 12'h888;
rom[27185] = 12'h888;
rom[27186] = 12'h999;
rom[27187] = 12'h999;
rom[27188] = 12'h999;
rom[27189] = 12'h999;
rom[27190] = 12'h999;
rom[27191] = 12'h888;
rom[27192] = 12'h888;
rom[27193] = 12'h999;
rom[27194] = 12'h999;
rom[27195] = 12'h999;
rom[27196] = 12'haaa;
rom[27197] = 12'haaa;
rom[27198] = 12'haaa;
rom[27199] = 12'haaa;
rom[27200] = 12'h666;
rom[27201] = 12'h666;
rom[27202] = 12'h666;
rom[27203] = 12'h555;
rom[27204] = 12'h555;
rom[27205] = 12'h555;
rom[27206] = 12'h555;
rom[27207] = 12'h555;
rom[27208] = 12'h555;
rom[27209] = 12'h555;
rom[27210] = 12'h555;
rom[27211] = 12'h555;
rom[27212] = 12'h555;
rom[27213] = 12'h555;
rom[27214] = 12'h555;
rom[27215] = 12'h555;
rom[27216] = 12'h666;
rom[27217] = 12'h666;
rom[27218] = 12'h666;
rom[27219] = 12'h666;
rom[27220] = 12'h666;
rom[27221] = 12'h666;
rom[27222] = 12'h666;
rom[27223] = 12'h666;
rom[27224] = 12'h666;
rom[27225] = 12'h666;
rom[27226] = 12'h666;
rom[27227] = 12'h666;
rom[27228] = 12'h777;
rom[27229] = 12'h777;
rom[27230] = 12'h777;
rom[27231] = 12'h777;
rom[27232] = 12'h777;
rom[27233] = 12'h777;
rom[27234] = 12'h777;
rom[27235] = 12'h777;
rom[27236] = 12'h777;
rom[27237] = 12'h888;
rom[27238] = 12'h888;
rom[27239] = 12'h888;
rom[27240] = 12'h888;
rom[27241] = 12'h888;
rom[27242] = 12'h888;
rom[27243] = 12'h888;
rom[27244] = 12'h777;
rom[27245] = 12'h777;
rom[27246] = 12'h777;
rom[27247] = 12'h777;
rom[27248] = 12'h777;
rom[27249] = 12'h777;
rom[27250] = 12'h777;
rom[27251] = 12'h777;
rom[27252] = 12'h777;
rom[27253] = 12'h888;
rom[27254] = 12'h888;
rom[27255] = 12'h888;
rom[27256] = 12'h888;
rom[27257] = 12'h888;
rom[27258] = 12'h888;
rom[27259] = 12'h777;
rom[27260] = 12'h777;
rom[27261] = 12'h666;
rom[27262] = 12'h666;
rom[27263] = 12'h666;
rom[27264] = 12'h666;
rom[27265] = 12'h555;
rom[27266] = 12'h555;
rom[27267] = 12'h555;
rom[27268] = 12'h555;
rom[27269] = 12'h555;
rom[27270] = 12'h555;
rom[27271] = 12'h555;
rom[27272] = 12'h555;
rom[27273] = 12'h555;
rom[27274] = 12'h555;
rom[27275] = 12'h444;
rom[27276] = 12'h444;
rom[27277] = 12'h444;
rom[27278] = 12'h444;
rom[27279] = 12'h444;
rom[27280] = 12'h444;
rom[27281] = 12'h333;
rom[27282] = 12'h333;
rom[27283] = 12'h333;
rom[27284] = 12'h333;
rom[27285] = 12'h333;
rom[27286] = 12'h333;
rom[27287] = 12'h333;
rom[27288] = 12'h333;
rom[27289] = 12'h333;
rom[27290] = 12'h222;
rom[27291] = 12'h222;
rom[27292] = 12'h222;
rom[27293] = 12'h222;
rom[27294] = 12'h222;
rom[27295] = 12'h222;
rom[27296] = 12'h111;
rom[27297] = 12'h111;
rom[27298] = 12'h111;
rom[27299] = 12'h  0;
rom[27300] = 12'h  0;
rom[27301] = 12'h  0;
rom[27302] = 12'h  0;
rom[27303] = 12'h  0;
rom[27304] = 12'h  0;
rom[27305] = 12'h  0;
rom[27306] = 12'h  0;
rom[27307] = 12'h  0;
rom[27308] = 12'h  0;
rom[27309] = 12'h  0;
rom[27310] = 12'h  0;
rom[27311] = 12'h  0;
rom[27312] = 12'h  0;
rom[27313] = 12'h  0;
rom[27314] = 12'h  0;
rom[27315] = 12'h  0;
rom[27316] = 12'h  0;
rom[27317] = 12'h  0;
rom[27318] = 12'h100;
rom[27319] = 12'h100;
rom[27320] = 12'h100;
rom[27321] = 12'h200;
rom[27322] = 12'h200;
rom[27323] = 12'h300;
rom[27324] = 12'h300;
rom[27325] = 12'h400;
rom[27326] = 12'h400;
rom[27327] = 12'h510;
rom[27328] = 12'h510;
rom[27329] = 12'h620;
rom[27330] = 12'h720;
rom[27331] = 12'h830;
rom[27332] = 12'h940;
rom[27333] = 12'ha40;
rom[27334] = 12'hb50;
rom[27335] = 12'hc60;
rom[27336] = 12'hd60;
rom[27337] = 12'hd60;
rom[27338] = 12'he60;
rom[27339] = 12'he70;
rom[27340] = 12'he70;
rom[27341] = 12'he70;
rom[27342] = 12'he60;
rom[27343] = 12'he60;
rom[27344] = 12'hf61;
rom[27345] = 12'he61;
rom[27346] = 12'he60;
rom[27347] = 12'he60;
rom[27348] = 12'hf61;
rom[27349] = 12'hf61;
rom[27350] = 12'hf51;
rom[27351] = 12'hf51;
rom[27352] = 12'hf51;
rom[27353] = 12'he51;
rom[27354] = 12'he51;
rom[27355] = 12'he41;
rom[27356] = 12'he41;
rom[27357] = 12'hd41;
rom[27358] = 12'hd41;
rom[27359] = 12'hd41;
rom[27360] = 12'hb30;
rom[27361] = 12'hb30;
rom[27362] = 12'ha20;
rom[27363] = 12'h920;
rom[27364] = 12'h920;
rom[27365] = 12'h820;
rom[27366] = 12'h810;
rom[27367] = 12'h710;
rom[27368] = 12'h610;
rom[27369] = 12'h610;
rom[27370] = 12'h500;
rom[27371] = 12'h500;
rom[27372] = 12'h400;
rom[27373] = 12'h400;
rom[27374] = 12'h400;
rom[27375] = 12'h300;
rom[27376] = 12'h300;
rom[27377] = 12'h300;
rom[27378] = 12'h300;
rom[27379] = 12'h200;
rom[27380] = 12'h200;
rom[27381] = 12'h200;
rom[27382] = 12'h200;
rom[27383] = 12'h100;
rom[27384] = 12'h100;
rom[27385] = 12'h100;
rom[27386] = 12'h211;
rom[27387] = 12'h322;
rom[27388] = 12'h222;
rom[27389] = 12'h111;
rom[27390] = 12'h111;
rom[27391] = 12'h111;
rom[27392] = 12'h111;
rom[27393] = 12'h111;
rom[27394] = 12'h111;
rom[27395] = 12'h111;
rom[27396] = 12'h222;
rom[27397] = 12'h222;
rom[27398] = 12'h222;
rom[27399] = 12'h222;
rom[27400] = 12'h222;
rom[27401] = 12'h333;
rom[27402] = 12'h333;
rom[27403] = 12'h444;
rom[27404] = 12'h555;
rom[27405] = 12'h777;
rom[27406] = 12'h888;
rom[27407] = 12'h888;
rom[27408] = 12'h888;
rom[27409] = 12'h888;
rom[27410] = 12'h999;
rom[27411] = 12'h999;
rom[27412] = 12'h999;
rom[27413] = 12'h888;
rom[27414] = 12'h888;
rom[27415] = 12'h888;
rom[27416] = 12'h777;
rom[27417] = 12'h777;
rom[27418] = 12'h777;
rom[27419] = 12'h777;
rom[27420] = 12'h777;
rom[27421] = 12'h777;
rom[27422] = 12'h777;
rom[27423] = 12'h777;
rom[27424] = 12'h777;
rom[27425] = 12'h777;
rom[27426] = 12'h777;
rom[27427] = 12'h777;
rom[27428] = 12'h777;
rom[27429] = 12'h777;
rom[27430] = 12'h777;
rom[27431] = 12'h777;
rom[27432] = 12'h777;
rom[27433] = 12'h777;
rom[27434] = 12'h666;
rom[27435] = 12'h666;
rom[27436] = 12'h666;
rom[27437] = 12'h555;
rom[27438] = 12'h555;
rom[27439] = 12'h555;
rom[27440] = 12'h444;
rom[27441] = 12'h444;
rom[27442] = 12'h444;
rom[27443] = 12'h444;
rom[27444] = 12'h444;
rom[27445] = 12'h333;
rom[27446] = 12'h333;
rom[27447] = 12'h333;
rom[27448] = 12'h333;
rom[27449] = 12'h222;
rom[27450] = 12'h222;
rom[27451] = 12'h111;
rom[27452] = 12'h111;
rom[27453] = 12'h111;
rom[27454] = 12'h111;
rom[27455] = 12'h  0;
rom[27456] = 12'h  0;
rom[27457] = 12'h  0;
rom[27458] = 12'h  0;
rom[27459] = 12'h  0;
rom[27460] = 12'h  0;
rom[27461] = 12'h  0;
rom[27462] = 12'h  0;
rom[27463] = 12'h  0;
rom[27464] = 12'h  0;
rom[27465] = 12'h  0;
rom[27466] = 12'h  0;
rom[27467] = 12'h  0;
rom[27468] = 12'h  0;
rom[27469] = 12'h  0;
rom[27470] = 12'h  0;
rom[27471] = 12'h  0;
rom[27472] = 12'h  0;
rom[27473] = 12'h  0;
rom[27474] = 12'h  0;
rom[27475] = 12'h  0;
rom[27476] = 12'h  0;
rom[27477] = 12'h  0;
rom[27478] = 12'h  0;
rom[27479] = 12'h  0;
rom[27480] = 12'h  0;
rom[27481] = 12'h  0;
rom[27482] = 12'h  0;
rom[27483] = 12'h  0;
rom[27484] = 12'h  0;
rom[27485] = 12'h  0;
rom[27486] = 12'h  0;
rom[27487] = 12'h  0;
rom[27488] = 12'h  0;
rom[27489] = 12'h  0;
rom[27490] = 12'h111;
rom[27491] = 12'h111;
rom[27492] = 12'h111;
rom[27493] = 12'h111;
rom[27494] = 12'h111;
rom[27495] = 12'h222;
rom[27496] = 12'h222;
rom[27497] = 12'h222;
rom[27498] = 12'h222;
rom[27499] = 12'h222;
rom[27500] = 12'h222;
rom[27501] = 12'h222;
rom[27502] = 12'h333;
rom[27503] = 12'h333;
rom[27504] = 12'h444;
rom[27505] = 12'h555;
rom[27506] = 12'h455;
rom[27507] = 12'h444;
rom[27508] = 12'h455;
rom[27509] = 12'h555;
rom[27510] = 12'h555;
rom[27511] = 12'h555;
rom[27512] = 12'h566;
rom[27513] = 12'h666;
rom[27514] = 12'h666;
rom[27515] = 12'h666;
rom[27516] = 12'h777;
rom[27517] = 12'h788;
rom[27518] = 12'h888;
rom[27519] = 12'h999;
rom[27520] = 12'h999;
rom[27521] = 12'haaa;
rom[27522] = 12'hbba;
rom[27523] = 12'hccb;
rom[27524] = 12'hddd;
rom[27525] = 12'hffe;
rom[27526] = 12'hfff;
rom[27527] = 12'hffe;
rom[27528] = 12'hffe;
rom[27529] = 12'hedd;
rom[27530] = 12'hcba;
rom[27531] = 12'ha98;
rom[27532] = 12'h977;
rom[27533] = 12'h755;
rom[27534] = 12'h533;
rom[27535] = 12'h421;
rom[27536] = 12'h310;
rom[27537] = 12'h310;
rom[27538] = 12'h410;
rom[27539] = 12'h420;
rom[27540] = 12'h521;
rom[27541] = 12'h621;
rom[27542] = 12'h621;
rom[27543] = 12'h720;
rom[27544] = 12'h720;
rom[27545] = 12'h830;
rom[27546] = 12'h830;
rom[27547] = 12'h930;
rom[27548] = 12'h930;
rom[27549] = 12'h930;
rom[27550] = 12'h930;
rom[27551] = 12'h930;
rom[27552] = 12'h940;
rom[27553] = 12'h940;
rom[27554] = 12'h840;
rom[27555] = 12'h840;
rom[27556] = 12'h740;
rom[27557] = 12'h740;
rom[27558] = 12'h851;
rom[27559] = 12'h852;
rom[27560] = 12'h852;
rom[27561] = 12'h852;
rom[27562] = 12'h852;
rom[27563] = 12'h852;
rom[27564] = 12'h742;
rom[27565] = 12'h642;
rom[27566] = 12'h642;
rom[27567] = 12'h542;
rom[27568] = 12'h542;
rom[27569] = 12'h542;
rom[27570] = 12'h653;
rom[27571] = 12'h654;
rom[27572] = 12'h765;
rom[27573] = 12'h766;
rom[27574] = 12'h776;
rom[27575] = 12'h777;
rom[27576] = 12'h877;
rom[27577] = 12'h888;
rom[27578] = 12'h888;
rom[27579] = 12'h888;
rom[27580] = 12'h888;
rom[27581] = 12'h888;
rom[27582] = 12'h888;
rom[27583] = 12'h888;
rom[27584] = 12'h888;
rom[27585] = 12'h888;
rom[27586] = 12'h888;
rom[27587] = 12'h999;
rom[27588] = 12'h999;
rom[27589] = 12'h999;
rom[27590] = 12'h999;
rom[27591] = 12'h999;
rom[27592] = 12'h888;
rom[27593] = 12'h999;
rom[27594] = 12'h999;
rom[27595] = 12'h999;
rom[27596] = 12'haaa;
rom[27597] = 12'haaa;
rom[27598] = 12'haaa;
rom[27599] = 12'haaa;
rom[27600] = 12'h666;
rom[27601] = 12'h666;
rom[27602] = 12'h666;
rom[27603] = 12'h555;
rom[27604] = 12'h555;
rom[27605] = 12'h555;
rom[27606] = 12'h555;
rom[27607] = 12'h555;
rom[27608] = 12'h666;
rom[27609] = 12'h555;
rom[27610] = 12'h555;
rom[27611] = 12'h555;
rom[27612] = 12'h555;
rom[27613] = 12'h555;
rom[27614] = 12'h555;
rom[27615] = 12'h555;
rom[27616] = 12'h666;
rom[27617] = 12'h555;
rom[27618] = 12'h555;
rom[27619] = 12'h666;
rom[27620] = 12'h666;
rom[27621] = 12'h666;
rom[27622] = 12'h666;
rom[27623] = 12'h666;
rom[27624] = 12'h666;
rom[27625] = 12'h666;
rom[27626] = 12'h666;
rom[27627] = 12'h666;
rom[27628] = 12'h666;
rom[27629] = 12'h777;
rom[27630] = 12'h777;
rom[27631] = 12'h777;
rom[27632] = 12'h777;
rom[27633] = 12'h777;
rom[27634] = 12'h777;
rom[27635] = 12'h777;
rom[27636] = 12'h888;
rom[27637] = 12'h888;
rom[27638] = 12'h888;
rom[27639] = 12'h888;
rom[27640] = 12'h888;
rom[27641] = 12'h888;
rom[27642] = 12'h888;
rom[27643] = 12'h888;
rom[27644] = 12'h777;
rom[27645] = 12'h777;
rom[27646] = 12'h777;
rom[27647] = 12'h777;
rom[27648] = 12'h777;
rom[27649] = 12'h777;
rom[27650] = 12'h777;
rom[27651] = 12'h777;
rom[27652] = 12'h777;
rom[27653] = 12'h777;
rom[27654] = 12'h888;
rom[27655] = 12'h888;
rom[27656] = 12'h888;
rom[27657] = 12'h888;
rom[27658] = 12'h888;
rom[27659] = 12'h888;
rom[27660] = 12'h777;
rom[27661] = 12'h666;
rom[27662] = 12'h666;
rom[27663] = 12'h666;
rom[27664] = 12'h666;
rom[27665] = 12'h555;
rom[27666] = 12'h555;
rom[27667] = 12'h555;
rom[27668] = 12'h555;
rom[27669] = 12'h555;
rom[27670] = 12'h555;
rom[27671] = 12'h555;
rom[27672] = 12'h555;
rom[27673] = 12'h555;
rom[27674] = 12'h555;
rom[27675] = 12'h444;
rom[27676] = 12'h444;
rom[27677] = 12'h444;
rom[27678] = 12'h444;
rom[27679] = 12'h444;
rom[27680] = 12'h333;
rom[27681] = 12'h333;
rom[27682] = 12'h333;
rom[27683] = 12'h333;
rom[27684] = 12'h333;
rom[27685] = 12'h333;
rom[27686] = 12'h333;
rom[27687] = 12'h333;
rom[27688] = 12'h333;
rom[27689] = 12'h333;
rom[27690] = 12'h222;
rom[27691] = 12'h222;
rom[27692] = 12'h222;
rom[27693] = 12'h222;
rom[27694] = 12'h222;
rom[27695] = 12'h111;
rom[27696] = 12'h111;
rom[27697] = 12'h111;
rom[27698] = 12'h111;
rom[27699] = 12'h111;
rom[27700] = 12'h  0;
rom[27701] = 12'h  0;
rom[27702] = 12'h  0;
rom[27703] = 12'h  0;
rom[27704] = 12'h  0;
rom[27705] = 12'h  0;
rom[27706] = 12'h  0;
rom[27707] = 12'h  0;
rom[27708] = 12'h  0;
rom[27709] = 12'h  0;
rom[27710] = 12'h  0;
rom[27711] = 12'h  0;
rom[27712] = 12'h  0;
rom[27713] = 12'h  0;
rom[27714] = 12'h  0;
rom[27715] = 12'h  0;
rom[27716] = 12'h  0;
rom[27717] = 12'h  0;
rom[27718] = 12'h  0;
rom[27719] = 12'h100;
rom[27720] = 12'h100;
rom[27721] = 12'h100;
rom[27722] = 12'h200;
rom[27723] = 12'h200;
rom[27724] = 12'h300;
rom[27725] = 12'h300;
rom[27726] = 12'h300;
rom[27727] = 12'h400;
rom[27728] = 12'h410;
rom[27729] = 12'h510;
rom[27730] = 12'h620;
rom[27731] = 12'h720;
rom[27732] = 12'h830;
rom[27733] = 12'h940;
rom[27734] = 12'ha40;
rom[27735] = 12'hb50;
rom[27736] = 12'hc50;
rom[27737] = 12'hc60;
rom[27738] = 12'hd60;
rom[27739] = 12'hd60;
rom[27740] = 12'he60;
rom[27741] = 12'he60;
rom[27742] = 12'he60;
rom[27743] = 12'he60;
rom[27744] = 12'he60;
rom[27745] = 12'he50;
rom[27746] = 12'he50;
rom[27747] = 12'he50;
rom[27748] = 12'he51;
rom[27749] = 12'hf51;
rom[27750] = 12'hf51;
rom[27751] = 12'he51;
rom[27752] = 12'he51;
rom[27753] = 12'he41;
rom[27754] = 12'he41;
rom[27755] = 12'hd41;
rom[27756] = 12'hd41;
rom[27757] = 12'hd30;
rom[27758] = 12'hc30;
rom[27759] = 12'hc30;
rom[27760] = 12'ha20;
rom[27761] = 12'h920;
rom[27762] = 12'h920;
rom[27763] = 12'h810;
rom[27764] = 12'h810;
rom[27765] = 12'h710;
rom[27766] = 12'h710;
rom[27767] = 12'h610;
rom[27768] = 12'h600;
rom[27769] = 12'h500;
rom[27770] = 12'h400;
rom[27771] = 12'h400;
rom[27772] = 12'h400;
rom[27773] = 12'h300;
rom[27774] = 12'h300;
rom[27775] = 12'h300;
rom[27776] = 12'h300;
rom[27777] = 12'h200;
rom[27778] = 12'h200;
rom[27779] = 12'h200;
rom[27780] = 12'h200;
rom[27781] = 12'h200;
rom[27782] = 12'h100;
rom[27783] = 12'h100;
rom[27784] = 12'h100;
rom[27785] = 12'h100;
rom[27786] = 12'h222;
rom[27787] = 12'h322;
rom[27788] = 12'h212;
rom[27789] = 12'h101;
rom[27790] = 12'h101;
rom[27791] = 12'h111;
rom[27792] = 12'h111;
rom[27793] = 12'h111;
rom[27794] = 12'h111;
rom[27795] = 12'h111;
rom[27796] = 12'h111;
rom[27797] = 12'h222;
rom[27798] = 12'h222;
rom[27799] = 12'h222;
rom[27800] = 12'h222;
rom[27801] = 12'h333;
rom[27802] = 12'h333;
rom[27803] = 12'h444;
rom[27804] = 12'h555;
rom[27805] = 12'h666;
rom[27806] = 12'h888;
rom[27807] = 12'h888;
rom[27808] = 12'h888;
rom[27809] = 12'h888;
rom[27810] = 12'h888;
rom[27811] = 12'h999;
rom[27812] = 12'h888;
rom[27813] = 12'h888;
rom[27814] = 12'h888;
rom[27815] = 12'h888;
rom[27816] = 12'h777;
rom[27817] = 12'h777;
rom[27818] = 12'h777;
rom[27819] = 12'h777;
rom[27820] = 12'h777;
rom[27821] = 12'h777;
rom[27822] = 12'h777;
rom[27823] = 12'h777;
rom[27824] = 12'h777;
rom[27825] = 12'h777;
rom[27826] = 12'h777;
rom[27827] = 12'h777;
rom[27828] = 12'h777;
rom[27829] = 12'h777;
rom[27830] = 12'h777;
rom[27831] = 12'h777;
rom[27832] = 12'h777;
rom[27833] = 12'h777;
rom[27834] = 12'h666;
rom[27835] = 12'h666;
rom[27836] = 12'h666;
rom[27837] = 12'h555;
rom[27838] = 12'h555;
rom[27839] = 12'h555;
rom[27840] = 12'h444;
rom[27841] = 12'h444;
rom[27842] = 12'h444;
rom[27843] = 12'h444;
rom[27844] = 12'h444;
rom[27845] = 12'h333;
rom[27846] = 12'h333;
rom[27847] = 12'h222;
rom[27848] = 12'h222;
rom[27849] = 12'h222;
rom[27850] = 12'h111;
rom[27851] = 12'h111;
rom[27852] = 12'h111;
rom[27853] = 12'h111;
rom[27854] = 12'h  0;
rom[27855] = 12'h  0;
rom[27856] = 12'h  0;
rom[27857] = 12'h  0;
rom[27858] = 12'h  0;
rom[27859] = 12'h  0;
rom[27860] = 12'h  0;
rom[27861] = 12'h  0;
rom[27862] = 12'h  0;
rom[27863] = 12'h  0;
rom[27864] = 12'h  0;
rom[27865] = 12'h  0;
rom[27866] = 12'h  0;
rom[27867] = 12'h  0;
rom[27868] = 12'h  0;
rom[27869] = 12'h  0;
rom[27870] = 12'h  0;
rom[27871] = 12'h  0;
rom[27872] = 12'h  0;
rom[27873] = 12'h  0;
rom[27874] = 12'h  0;
rom[27875] = 12'h  0;
rom[27876] = 12'h  0;
rom[27877] = 12'h  0;
rom[27878] = 12'h  0;
rom[27879] = 12'h  0;
rom[27880] = 12'h  0;
rom[27881] = 12'h  0;
rom[27882] = 12'h  0;
rom[27883] = 12'h  0;
rom[27884] = 12'h  0;
rom[27885] = 12'h  0;
rom[27886] = 12'h  0;
rom[27887] = 12'h  0;
rom[27888] = 12'h  0;
rom[27889] = 12'h111;
rom[27890] = 12'h111;
rom[27891] = 12'h111;
rom[27892] = 12'h111;
rom[27893] = 12'h111;
rom[27894] = 12'h111;
rom[27895] = 12'h222;
rom[27896] = 12'h222;
rom[27897] = 12'h222;
rom[27898] = 12'h222;
rom[27899] = 12'h222;
rom[27900] = 12'h222;
rom[27901] = 12'h333;
rom[27902] = 12'h333;
rom[27903] = 12'h444;
rom[27904] = 12'h555;
rom[27905] = 12'h555;
rom[27906] = 12'h555;
rom[27907] = 12'h445;
rom[27908] = 12'h555;
rom[27909] = 12'h555;
rom[27910] = 12'h666;
rom[27911] = 12'h666;
rom[27912] = 12'h666;
rom[27913] = 12'h666;
rom[27914] = 12'h666;
rom[27915] = 12'h777;
rom[27916] = 12'h777;
rom[27917] = 12'h888;
rom[27918] = 12'h999;
rom[27919] = 12'h999;
rom[27920] = 12'haaa;
rom[27921] = 12'hcbb;
rom[27922] = 12'hddd;
rom[27923] = 12'heee;
rom[27924] = 12'hffe;
rom[27925] = 12'hfff;
rom[27926] = 12'hfff;
rom[27927] = 12'hffe;
rom[27928] = 12'hcbb;
rom[27929] = 12'ha98;
rom[27930] = 12'h755;
rom[27931] = 12'h532;
rom[27932] = 12'h421;
rom[27933] = 12'h421;
rom[27934] = 12'h411;
rom[27935] = 12'h410;
rom[27936] = 12'h421;
rom[27937] = 12'h410;
rom[27938] = 12'h410;
rom[27939] = 12'h520;
rom[27940] = 12'h521;
rom[27941] = 12'h621;
rom[27942] = 12'h720;
rom[27943] = 12'h720;
rom[27944] = 12'h720;
rom[27945] = 12'h820;
rom[27946] = 12'h920;
rom[27947] = 12'h930;
rom[27948] = 12'ha30;
rom[27949] = 12'ha30;
rom[27950] = 12'ha30;
rom[27951] = 12'ha30;
rom[27952] = 12'ha30;
rom[27953] = 12'h930;
rom[27954] = 12'h930;
rom[27955] = 12'h830;
rom[27956] = 12'h830;
rom[27957] = 12'h840;
rom[27958] = 12'h851;
rom[27959] = 12'h952;
rom[27960] = 12'h952;
rom[27961] = 12'h952;
rom[27962] = 12'h852;
rom[27963] = 12'h852;
rom[27964] = 12'h742;
rom[27965] = 12'h741;
rom[27966] = 12'h641;
rom[27967] = 12'h531;
rom[27968] = 12'h531;
rom[27969] = 12'h532;
rom[27970] = 12'h642;
rom[27971] = 12'h643;
rom[27972] = 12'h654;
rom[27973] = 12'h654;
rom[27974] = 12'h765;
rom[27975] = 12'h766;
rom[27976] = 12'h777;
rom[27977] = 12'h877;
rom[27978] = 12'h888;
rom[27979] = 12'h888;
rom[27980] = 12'h888;
rom[27981] = 12'h888;
rom[27982] = 12'h888;
rom[27983] = 12'h888;
rom[27984] = 12'h888;
rom[27985] = 12'h888;
rom[27986] = 12'h888;
rom[27987] = 12'h888;
rom[27988] = 12'h999;
rom[27989] = 12'h999;
rom[27990] = 12'h999;
rom[27991] = 12'h999;
rom[27992] = 12'h999;
rom[27993] = 12'h999;
rom[27994] = 12'h999;
rom[27995] = 12'h999;
rom[27996] = 12'haaa;
rom[27997] = 12'haaa;
rom[27998] = 12'haaa;
rom[27999] = 12'haaa;
rom[28000] = 12'h666;
rom[28001] = 12'h666;
rom[28002] = 12'h666;
rom[28003] = 12'h555;
rom[28004] = 12'h555;
rom[28005] = 12'h555;
rom[28006] = 12'h555;
rom[28007] = 12'h555;
rom[28008] = 12'h666;
rom[28009] = 12'h666;
rom[28010] = 12'h666;
rom[28011] = 12'h666;
rom[28012] = 12'h666;
rom[28013] = 12'h555;
rom[28014] = 12'h555;
rom[28015] = 12'h555;
rom[28016] = 12'h666;
rom[28017] = 12'h555;
rom[28018] = 12'h555;
rom[28019] = 12'h666;
rom[28020] = 12'h666;
rom[28021] = 12'h666;
rom[28022] = 12'h666;
rom[28023] = 12'h666;
rom[28024] = 12'h666;
rom[28025] = 12'h666;
rom[28026] = 12'h666;
rom[28027] = 12'h666;
rom[28028] = 12'h666;
rom[28029] = 12'h777;
rom[28030] = 12'h777;
rom[28031] = 12'h777;
rom[28032] = 12'h777;
rom[28033] = 12'h777;
rom[28034] = 12'h777;
rom[28035] = 12'h888;
rom[28036] = 12'h888;
rom[28037] = 12'h888;
rom[28038] = 12'h888;
rom[28039] = 12'h888;
rom[28040] = 12'h888;
rom[28041] = 12'h888;
rom[28042] = 12'h888;
rom[28043] = 12'h888;
rom[28044] = 12'h777;
rom[28045] = 12'h777;
rom[28046] = 12'h777;
rom[28047] = 12'h777;
rom[28048] = 12'h777;
rom[28049] = 12'h777;
rom[28050] = 12'h666;
rom[28051] = 12'h666;
rom[28052] = 12'h666;
rom[28053] = 12'h777;
rom[28054] = 12'h777;
rom[28055] = 12'h777;
rom[28056] = 12'h888;
rom[28057] = 12'h888;
rom[28058] = 12'h888;
rom[28059] = 12'h888;
rom[28060] = 12'h888;
rom[28061] = 12'h777;
rom[28062] = 12'h666;
rom[28063] = 12'h666;
rom[28064] = 12'h666;
rom[28065] = 12'h666;
rom[28066] = 12'h555;
rom[28067] = 12'h555;
rom[28068] = 12'h555;
rom[28069] = 12'h555;
rom[28070] = 12'h555;
rom[28071] = 12'h555;
rom[28072] = 12'h555;
rom[28073] = 12'h555;
rom[28074] = 12'h555;
rom[28075] = 12'h444;
rom[28076] = 12'h444;
rom[28077] = 12'h444;
rom[28078] = 12'h444;
rom[28079] = 12'h444;
rom[28080] = 12'h333;
rom[28081] = 12'h333;
rom[28082] = 12'h333;
rom[28083] = 12'h333;
rom[28084] = 12'h222;
rom[28085] = 12'h222;
rom[28086] = 12'h333;
rom[28087] = 12'h333;
rom[28088] = 12'h333;
rom[28089] = 12'h333;
rom[28090] = 12'h222;
rom[28091] = 12'h222;
rom[28092] = 12'h222;
rom[28093] = 12'h222;
rom[28094] = 12'h111;
rom[28095] = 12'h111;
rom[28096] = 12'h111;
rom[28097] = 12'h111;
rom[28098] = 12'h111;
rom[28099] = 12'h111;
rom[28100] = 12'h  0;
rom[28101] = 12'h  0;
rom[28102] = 12'h  0;
rom[28103] = 12'h  0;
rom[28104] = 12'h  0;
rom[28105] = 12'h  0;
rom[28106] = 12'h  0;
rom[28107] = 12'h  0;
rom[28108] = 12'h  0;
rom[28109] = 12'h  0;
rom[28110] = 12'h  0;
rom[28111] = 12'h  0;
rom[28112] = 12'h  0;
rom[28113] = 12'h  0;
rom[28114] = 12'h  0;
rom[28115] = 12'h  0;
rom[28116] = 12'h  0;
rom[28117] = 12'h  0;
rom[28118] = 12'h  0;
rom[28119] = 12'h  0;
rom[28120] = 12'h100;
rom[28121] = 12'h100;
rom[28122] = 12'h100;
rom[28123] = 12'h200;
rom[28124] = 12'h200;
rom[28125] = 12'h200;
rom[28126] = 12'h300;
rom[28127] = 12'h300;
rom[28128] = 12'h410;
rom[28129] = 12'h410;
rom[28130] = 12'h510;
rom[28131] = 12'h620;
rom[28132] = 12'h620;
rom[28133] = 12'h730;
rom[28134] = 12'h830;
rom[28135] = 12'h940;
rom[28136] = 12'ha40;
rom[28137] = 12'hb40;
rom[28138] = 12'hc50;
rom[28139] = 12'hc50;
rom[28140] = 12'hd50;
rom[28141] = 12'hd50;
rom[28142] = 12'hd50;
rom[28143] = 12'hd50;
rom[28144] = 12'he50;
rom[28145] = 12'he50;
rom[28146] = 12'he50;
rom[28147] = 12'he50;
rom[28148] = 12'he50;
rom[28149] = 12'he51;
rom[28150] = 12'he41;
rom[28151] = 12'he41;
rom[28152] = 12'he41;
rom[28153] = 12'hd40;
rom[28154] = 12'hd30;
rom[28155] = 12'hd30;
rom[28156] = 12'hc30;
rom[28157] = 12'hc20;
rom[28158] = 12'hb20;
rom[28159] = 12'hb20;
rom[28160] = 12'h920;
rom[28161] = 12'h810;
rom[28162] = 12'h810;
rom[28163] = 12'h710;
rom[28164] = 12'h710;
rom[28165] = 12'h610;
rom[28166] = 12'h600;
rom[28167] = 12'h500;
rom[28168] = 12'h500;
rom[28169] = 12'h400;
rom[28170] = 12'h400;
rom[28171] = 12'h300;
rom[28172] = 12'h300;
rom[28173] = 12'h300;
rom[28174] = 12'h200;
rom[28175] = 12'h200;
rom[28176] = 12'h200;
rom[28177] = 12'h200;
rom[28178] = 12'h200;
rom[28179] = 12'h200;
rom[28180] = 12'h200;
rom[28181] = 12'h100;
rom[28182] = 12'h100;
rom[28183] = 12'h100;
rom[28184] = 12'h100;
rom[28185] = 12'h211;
rom[28186] = 12'h322;
rom[28187] = 12'h222;
rom[28188] = 12'h111;
rom[28189] = 12'h  0;
rom[28190] = 12'h  0;
rom[28191] = 12'h111;
rom[28192] = 12'h111;
rom[28193] = 12'h111;
rom[28194] = 12'h111;
rom[28195] = 12'h111;
rom[28196] = 12'h111;
rom[28197] = 12'h222;
rom[28198] = 12'h222;
rom[28199] = 12'h222;
rom[28200] = 12'h222;
rom[28201] = 12'h333;
rom[28202] = 12'h333;
rom[28203] = 12'h333;
rom[28204] = 12'h555;
rom[28205] = 12'h666;
rom[28206] = 12'h777;
rom[28207] = 12'h888;
rom[28208] = 12'h888;
rom[28209] = 12'h888;
rom[28210] = 12'h888;
rom[28211] = 12'h888;
rom[28212] = 12'h888;
rom[28213] = 12'h888;
rom[28214] = 12'h888;
rom[28215] = 12'h777;
rom[28216] = 12'h777;
rom[28217] = 12'h777;
rom[28218] = 12'h777;
rom[28219] = 12'h777;
rom[28220] = 12'h777;
rom[28221] = 12'h777;
rom[28222] = 12'h777;
rom[28223] = 12'h777;
rom[28224] = 12'h777;
rom[28225] = 12'h777;
rom[28226] = 12'h777;
rom[28227] = 12'h777;
rom[28228] = 12'h777;
rom[28229] = 12'h777;
rom[28230] = 12'h777;
rom[28231] = 12'h777;
rom[28232] = 12'h777;
rom[28233] = 12'h777;
rom[28234] = 12'h666;
rom[28235] = 12'h666;
rom[28236] = 12'h666;
rom[28237] = 12'h555;
rom[28238] = 12'h555;
rom[28239] = 12'h555;
rom[28240] = 12'h555;
rom[28241] = 12'h555;
rom[28242] = 12'h444;
rom[28243] = 12'h444;
rom[28244] = 12'h333;
rom[28245] = 12'h333;
rom[28246] = 12'h222;
rom[28247] = 12'h222;
rom[28248] = 12'h222;
rom[28249] = 12'h111;
rom[28250] = 12'h111;
rom[28251] = 12'h111;
rom[28252] = 12'h111;
rom[28253] = 12'h111;
rom[28254] = 12'h  0;
rom[28255] = 12'h  0;
rom[28256] = 12'h111;
rom[28257] = 12'h  0;
rom[28258] = 12'h  0;
rom[28259] = 12'h  0;
rom[28260] = 12'h  0;
rom[28261] = 12'h  0;
rom[28262] = 12'h  0;
rom[28263] = 12'h  0;
rom[28264] = 12'h  0;
rom[28265] = 12'h  0;
rom[28266] = 12'h  0;
rom[28267] = 12'h  0;
rom[28268] = 12'h  0;
rom[28269] = 12'h  0;
rom[28270] = 12'h  0;
rom[28271] = 12'h  0;
rom[28272] = 12'h  0;
rom[28273] = 12'h  0;
rom[28274] = 12'h  0;
rom[28275] = 12'h  0;
rom[28276] = 12'h  0;
rom[28277] = 12'h  0;
rom[28278] = 12'h  0;
rom[28279] = 12'h  0;
rom[28280] = 12'h  0;
rom[28281] = 12'h  0;
rom[28282] = 12'h  0;
rom[28283] = 12'h  0;
rom[28284] = 12'h  0;
rom[28285] = 12'h  0;
rom[28286] = 12'h  0;
rom[28287] = 12'h  0;
rom[28288] = 12'h  0;
rom[28289] = 12'h111;
rom[28290] = 12'h111;
rom[28291] = 12'h111;
rom[28292] = 12'h111;
rom[28293] = 12'h111;
rom[28294] = 12'h222;
rom[28295] = 12'h222;
rom[28296] = 12'h222;
rom[28297] = 12'h222;
rom[28298] = 12'h222;
rom[28299] = 12'h222;
rom[28300] = 12'h333;
rom[28301] = 12'h333;
rom[28302] = 12'h444;
rom[28303] = 12'h444;
rom[28304] = 12'h555;
rom[28305] = 12'h555;
rom[28306] = 12'h555;
rom[28307] = 12'h555;
rom[28308] = 12'h555;
rom[28309] = 12'h666;
rom[28310] = 12'h666;
rom[28311] = 12'h666;
rom[28312] = 12'h666;
rom[28313] = 12'h777;
rom[28314] = 12'h777;
rom[28315] = 12'h777;
rom[28316] = 12'h888;
rom[28317] = 12'h999;
rom[28318] = 12'haaa;
rom[28319] = 12'hbbb;
rom[28320] = 12'hccc;
rom[28321] = 12'heed;
rom[28322] = 12'hfff;
rom[28323] = 12'hffe;
rom[28324] = 12'hfee;
rom[28325] = 12'hedd;
rom[28326] = 12'hcbb;
rom[28327] = 12'haa9;
rom[28328] = 12'h765;
rom[28329] = 12'h643;
rom[28330] = 12'h421;
rom[28331] = 12'h200;
rom[28332] = 12'h200;
rom[28333] = 12'h300;
rom[28334] = 12'h410;
rom[28335] = 12'h410;
rom[28336] = 12'h521;
rom[28337] = 12'h521;
rom[28338] = 12'h510;
rom[28339] = 12'h510;
rom[28340] = 12'h610;
rom[28341] = 12'h620;
rom[28342] = 12'h720;
rom[28343] = 12'h720;
rom[28344] = 12'h820;
rom[28345] = 12'h820;
rom[28346] = 12'h920;
rom[28347] = 12'ha30;
rom[28348] = 12'ha30;
rom[28349] = 12'hb30;
rom[28350] = 12'hb40;
rom[28351] = 12'hb40;
rom[28352] = 12'ha30;
rom[28353] = 12'ha30;
rom[28354] = 12'h930;
rom[28355] = 12'h930;
rom[28356] = 12'h830;
rom[28357] = 12'h840;
rom[28358] = 12'h951;
rom[28359] = 12'h962;
rom[28360] = 12'h952;
rom[28361] = 12'h951;
rom[28362] = 12'h951;
rom[28363] = 12'h841;
rom[28364] = 12'h841;
rom[28365] = 12'h741;
rom[28366] = 12'h641;
rom[28367] = 12'h631;
rom[28368] = 12'h631;
rom[28369] = 12'h542;
rom[28370] = 12'h642;
rom[28371] = 12'h642;
rom[28372] = 12'h643;
rom[28373] = 12'h654;
rom[28374] = 12'h665;
rom[28375] = 12'h765;
rom[28376] = 12'h776;
rom[28377] = 12'h777;
rom[28378] = 12'h887;
rom[28379] = 12'h888;
rom[28380] = 12'h888;
rom[28381] = 12'h888;
rom[28382] = 12'h888;
rom[28383] = 12'h888;
rom[28384] = 12'h888;
rom[28385] = 12'h888;
rom[28386] = 12'h888;
rom[28387] = 12'h888;
rom[28388] = 12'h888;
rom[28389] = 12'h888;
rom[28390] = 12'h888;
rom[28391] = 12'h888;
rom[28392] = 12'h999;
rom[28393] = 12'h999;
rom[28394] = 12'h999;
rom[28395] = 12'h999;
rom[28396] = 12'haaa;
rom[28397] = 12'haaa;
rom[28398] = 12'haaa;
rom[28399] = 12'haaa;
rom[28400] = 12'h666;
rom[28401] = 12'h666;
rom[28402] = 12'h666;
rom[28403] = 12'h555;
rom[28404] = 12'h555;
rom[28405] = 12'h555;
rom[28406] = 12'h555;
rom[28407] = 12'h555;
rom[28408] = 12'h666;
rom[28409] = 12'h666;
rom[28410] = 12'h666;
rom[28411] = 12'h666;
rom[28412] = 12'h666;
rom[28413] = 12'h666;
rom[28414] = 12'h666;
rom[28415] = 12'h666;
rom[28416] = 12'h666;
rom[28417] = 12'h666;
rom[28418] = 12'h666;
rom[28419] = 12'h666;
rom[28420] = 12'h666;
rom[28421] = 12'h666;
rom[28422] = 12'h666;
rom[28423] = 12'h666;
rom[28424] = 12'h666;
rom[28425] = 12'h666;
rom[28426] = 12'h666;
rom[28427] = 12'h666;
rom[28428] = 12'h777;
rom[28429] = 12'h777;
rom[28430] = 12'h777;
rom[28431] = 12'h777;
rom[28432] = 12'h777;
rom[28433] = 12'h777;
rom[28434] = 12'h777;
rom[28435] = 12'h888;
rom[28436] = 12'h888;
rom[28437] = 12'h888;
rom[28438] = 12'h888;
rom[28439] = 12'h888;
rom[28440] = 12'h888;
rom[28441] = 12'h888;
rom[28442] = 12'h888;
rom[28443] = 12'h888;
rom[28444] = 12'h777;
rom[28445] = 12'h777;
rom[28446] = 12'h777;
rom[28447] = 12'h777;
rom[28448] = 12'h777;
rom[28449] = 12'h666;
rom[28450] = 12'h666;
rom[28451] = 12'h666;
rom[28452] = 12'h666;
rom[28453] = 12'h666;
rom[28454] = 12'h777;
rom[28455] = 12'h777;
rom[28456] = 12'h888;
rom[28457] = 12'h888;
rom[28458] = 12'h888;
rom[28459] = 12'h888;
rom[28460] = 12'h888;
rom[28461] = 12'h777;
rom[28462] = 12'h777;
rom[28463] = 12'h666;
rom[28464] = 12'h666;
rom[28465] = 12'h666;
rom[28466] = 12'h555;
rom[28467] = 12'h555;
rom[28468] = 12'h555;
rom[28469] = 12'h555;
rom[28470] = 12'h555;
rom[28471] = 12'h555;
rom[28472] = 12'h555;
rom[28473] = 12'h555;
rom[28474] = 12'h444;
rom[28475] = 12'h444;
rom[28476] = 12'h444;
rom[28477] = 12'h444;
rom[28478] = 12'h444;
rom[28479] = 12'h444;
rom[28480] = 12'h333;
rom[28481] = 12'h333;
rom[28482] = 12'h333;
rom[28483] = 12'h333;
rom[28484] = 12'h222;
rom[28485] = 12'h222;
rom[28486] = 12'h222;
rom[28487] = 12'h333;
rom[28488] = 12'h333;
rom[28489] = 12'h333;
rom[28490] = 12'h222;
rom[28491] = 12'h222;
rom[28492] = 12'h222;
rom[28493] = 12'h111;
rom[28494] = 12'h111;
rom[28495] = 12'h111;
rom[28496] = 12'h111;
rom[28497] = 12'h111;
rom[28498] = 12'h111;
rom[28499] = 12'h111;
rom[28500] = 12'h  0;
rom[28501] = 12'h  0;
rom[28502] = 12'h  0;
rom[28503] = 12'h  0;
rom[28504] = 12'h  0;
rom[28505] = 12'h  0;
rom[28506] = 12'h  0;
rom[28507] = 12'h  0;
rom[28508] = 12'h  0;
rom[28509] = 12'h  0;
rom[28510] = 12'h  0;
rom[28511] = 12'h  0;
rom[28512] = 12'h  0;
rom[28513] = 12'h  0;
rom[28514] = 12'h  0;
rom[28515] = 12'h  0;
rom[28516] = 12'h  0;
rom[28517] = 12'h  0;
rom[28518] = 12'h  0;
rom[28519] = 12'h  0;
rom[28520] = 12'h100;
rom[28521] = 12'h100;
rom[28522] = 12'h100;
rom[28523] = 12'h100;
rom[28524] = 12'h200;
rom[28525] = 12'h200;
rom[28526] = 12'h200;
rom[28527] = 12'h200;
rom[28528] = 12'h300;
rom[28529] = 12'h310;
rom[28530] = 12'h410;
rom[28531] = 12'h520;
rom[28532] = 12'h520;
rom[28533] = 12'h620;
rom[28534] = 12'h730;
rom[28535] = 12'h830;
rom[28536] = 12'h930;
rom[28537] = 12'ha30;
rom[28538] = 12'ha40;
rom[28539] = 12'hb40;
rom[28540] = 12'hc40;
rom[28541] = 12'hc40;
rom[28542] = 12'hc40;
rom[28543] = 12'hc40;
rom[28544] = 12'hd51;
rom[28545] = 12'hd40;
rom[28546] = 12'hd40;
rom[28547] = 12'hd40;
rom[28548] = 12'hd40;
rom[28549] = 12'hd40;
rom[28550] = 12'hd40;
rom[28551] = 12'hd30;
rom[28552] = 12'hc30;
rom[28553] = 12'hc30;
rom[28554] = 12'hc30;
rom[28555] = 12'hc20;
rom[28556] = 12'hb20;
rom[28557] = 12'hb20;
rom[28558] = 12'hb20;
rom[28559] = 12'ha10;
rom[28560] = 12'h810;
rom[28561] = 12'h710;
rom[28562] = 12'h710;
rom[28563] = 12'h710;
rom[28564] = 12'h610;
rom[28565] = 12'h600;
rom[28566] = 12'h500;
rom[28567] = 12'h400;
rom[28568] = 12'h400;
rom[28569] = 12'h400;
rom[28570] = 12'h300;
rom[28571] = 12'h300;
rom[28572] = 12'h200;
rom[28573] = 12'h200;
rom[28574] = 12'h200;
rom[28575] = 12'h200;
rom[28576] = 12'h200;
rom[28577] = 12'h200;
rom[28578] = 12'h200;
rom[28579] = 12'h100;
rom[28580] = 12'h100;
rom[28581] = 12'h100;
rom[28582] = 12'h100;
rom[28583] = 12'h100;
rom[28584] = 12'h100;
rom[28585] = 12'h211;
rom[28586] = 12'h322;
rom[28587] = 12'h222;
rom[28588] = 12'h111;
rom[28589] = 12'h  0;
rom[28590] = 12'h  0;
rom[28591] = 12'h111;
rom[28592] = 12'h111;
rom[28593] = 12'h111;
rom[28594] = 12'h111;
rom[28595] = 12'h111;
rom[28596] = 12'h111;
rom[28597] = 12'h222;
rom[28598] = 12'h222;
rom[28599] = 12'h222;
rom[28600] = 12'h222;
rom[28601] = 12'h333;
rom[28602] = 12'h333;
rom[28603] = 12'h333;
rom[28604] = 12'h444;
rom[28605] = 12'h666;
rom[28606] = 12'h777;
rom[28607] = 12'h888;
rom[28608] = 12'h888;
rom[28609] = 12'h888;
rom[28610] = 12'h888;
rom[28611] = 12'h888;
rom[28612] = 12'h888;
rom[28613] = 12'h777;
rom[28614] = 12'h777;
rom[28615] = 12'h777;
rom[28616] = 12'h777;
rom[28617] = 12'h777;
rom[28618] = 12'h777;
rom[28619] = 12'h777;
rom[28620] = 12'h777;
rom[28621] = 12'h777;
rom[28622] = 12'h777;
rom[28623] = 12'h777;
rom[28624] = 12'h777;
rom[28625] = 12'h777;
rom[28626] = 12'h777;
rom[28627] = 12'h777;
rom[28628] = 12'h777;
rom[28629] = 12'h777;
rom[28630] = 12'h777;
rom[28631] = 12'h777;
rom[28632] = 12'h777;
rom[28633] = 12'h777;
rom[28634] = 12'h666;
rom[28635] = 12'h666;
rom[28636] = 12'h666;
rom[28637] = 12'h555;
rom[28638] = 12'h555;
rom[28639] = 12'h555;
rom[28640] = 12'h555;
rom[28641] = 12'h555;
rom[28642] = 12'h444;
rom[28643] = 12'h333;
rom[28644] = 12'h333;
rom[28645] = 12'h222;
rom[28646] = 12'h222;
rom[28647] = 12'h222;
rom[28648] = 12'h111;
rom[28649] = 12'h111;
rom[28650] = 12'h111;
rom[28651] = 12'h111;
rom[28652] = 12'h111;
rom[28653] = 12'h111;
rom[28654] = 12'h  0;
rom[28655] = 12'h  0;
rom[28656] = 12'h111;
rom[28657] = 12'h  0;
rom[28658] = 12'h  0;
rom[28659] = 12'h  0;
rom[28660] = 12'h  0;
rom[28661] = 12'h  0;
rom[28662] = 12'h  0;
rom[28663] = 12'h  0;
rom[28664] = 12'h  0;
rom[28665] = 12'h  0;
rom[28666] = 12'h  0;
rom[28667] = 12'h  0;
rom[28668] = 12'h  0;
rom[28669] = 12'h  0;
rom[28670] = 12'h  0;
rom[28671] = 12'h  0;
rom[28672] = 12'h  0;
rom[28673] = 12'h  0;
rom[28674] = 12'h  0;
rom[28675] = 12'h  0;
rom[28676] = 12'h  0;
rom[28677] = 12'h  0;
rom[28678] = 12'h  0;
rom[28679] = 12'h  0;
rom[28680] = 12'h  0;
rom[28681] = 12'h  0;
rom[28682] = 12'h  0;
rom[28683] = 12'h  0;
rom[28684] = 12'h  0;
rom[28685] = 12'h  0;
rom[28686] = 12'h  0;
rom[28687] = 12'h  0;
rom[28688] = 12'h  0;
rom[28689] = 12'h111;
rom[28690] = 12'h111;
rom[28691] = 12'h111;
rom[28692] = 12'h111;
rom[28693] = 12'h111;
rom[28694] = 12'h222;
rom[28695] = 12'h222;
rom[28696] = 12'h222;
rom[28697] = 12'h222;
rom[28698] = 12'h333;
rom[28699] = 12'h333;
rom[28700] = 12'h333;
rom[28701] = 12'h333;
rom[28702] = 12'h444;
rom[28703] = 12'h555;
rom[28704] = 12'h555;
rom[28705] = 12'h555;
rom[28706] = 12'h555;
rom[28707] = 12'h555;
rom[28708] = 12'h555;
rom[28709] = 12'h666;
rom[28710] = 12'h777;
rom[28711] = 12'h777;
rom[28712] = 12'h777;
rom[28713] = 12'h888;
rom[28714] = 12'h888;
rom[28715] = 12'h999;
rom[28716] = 12'haaa;
rom[28717] = 12'hbbb;
rom[28718] = 12'hccc;
rom[28719] = 12'hddd;
rom[28720] = 12'hfee;
rom[28721] = 12'hffe;
rom[28722] = 12'hffe;
rom[28723] = 12'heed;
rom[28724] = 12'hddc;
rom[28725] = 12'hbaa;
rom[28726] = 12'h766;
rom[28727] = 12'h432;
rom[28728] = 12'h321;
rom[28729] = 12'h311;
rom[28730] = 12'h310;
rom[28731] = 12'h310;
rom[28732] = 12'h310;
rom[28733] = 12'h310;
rom[28734] = 12'h400;
rom[28735] = 12'h400;
rom[28736] = 12'h400;
rom[28737] = 12'h410;
rom[28738] = 12'h410;
rom[28739] = 12'h510;
rom[28740] = 12'h610;
rom[28741] = 12'h620;
rom[28742] = 12'h710;
rom[28743] = 12'h710;
rom[28744] = 12'h820;
rom[28745] = 12'h920;
rom[28746] = 12'ha20;
rom[28747] = 12'ha30;
rom[28748] = 12'hb30;
rom[28749] = 12'hb30;
rom[28750] = 12'hc40;
rom[28751] = 12'hc40;
rom[28752] = 12'hb40;
rom[28753] = 12'hb40;
rom[28754] = 12'ha40;
rom[28755] = 12'h940;
rom[28756] = 12'h940;
rom[28757] = 12'h940;
rom[28758] = 12'ha51;
rom[28759] = 12'ha62;
rom[28760] = 12'ha62;
rom[28761] = 12'h951;
rom[28762] = 12'h941;
rom[28763] = 12'h840;
rom[28764] = 12'h840;
rom[28765] = 12'h741;
rom[28766] = 12'h741;
rom[28767] = 12'h641;
rom[28768] = 12'h641;
rom[28769] = 12'h642;
rom[28770] = 12'h642;
rom[28771] = 12'h642;
rom[28772] = 12'h643;
rom[28773] = 12'h653;
rom[28774] = 12'h654;
rom[28775] = 12'h765;
rom[28776] = 12'h766;
rom[28777] = 12'h776;
rom[28778] = 12'h777;
rom[28779] = 12'h888;
rom[28780] = 12'h888;
rom[28781] = 12'h888;
rom[28782] = 12'h888;
rom[28783] = 12'h888;
rom[28784] = 12'h999;
rom[28785] = 12'h999;
rom[28786] = 12'h888;
rom[28787] = 12'h888;
rom[28788] = 12'h888;
rom[28789] = 12'h888;
rom[28790] = 12'h888;
rom[28791] = 12'h888;
rom[28792] = 12'h999;
rom[28793] = 12'h999;
rom[28794] = 12'h999;
rom[28795] = 12'haaa;
rom[28796] = 12'haaa;
rom[28797] = 12'haaa;
rom[28798] = 12'haaa;
rom[28799] = 12'haaa;
rom[28800] = 12'h666;
rom[28801] = 12'h666;
rom[28802] = 12'h666;
rom[28803] = 12'h666;
rom[28804] = 12'h666;
rom[28805] = 12'h666;
rom[28806] = 12'h666;
rom[28807] = 12'h666;
rom[28808] = 12'h666;
rom[28809] = 12'h666;
rom[28810] = 12'h666;
rom[28811] = 12'h666;
rom[28812] = 12'h666;
rom[28813] = 12'h666;
rom[28814] = 12'h666;
rom[28815] = 12'h666;
rom[28816] = 12'h666;
rom[28817] = 12'h666;
rom[28818] = 12'h666;
rom[28819] = 12'h666;
rom[28820] = 12'h666;
rom[28821] = 12'h666;
rom[28822] = 12'h666;
rom[28823] = 12'h666;
rom[28824] = 12'h666;
rom[28825] = 12'h666;
rom[28826] = 12'h666;
rom[28827] = 12'h666;
rom[28828] = 12'h777;
rom[28829] = 12'h777;
rom[28830] = 12'h777;
rom[28831] = 12'h777;
rom[28832] = 12'h777;
rom[28833] = 12'h777;
rom[28834] = 12'h777;
rom[28835] = 12'h888;
rom[28836] = 12'h888;
rom[28837] = 12'h888;
rom[28838] = 12'h888;
rom[28839] = 12'h999;
rom[28840] = 12'h888;
rom[28841] = 12'h888;
rom[28842] = 12'h888;
rom[28843] = 12'h888;
rom[28844] = 12'h777;
rom[28845] = 12'h777;
rom[28846] = 12'h777;
rom[28847] = 12'h777;
rom[28848] = 12'h777;
rom[28849] = 12'h666;
rom[28850] = 12'h666;
rom[28851] = 12'h666;
rom[28852] = 12'h666;
rom[28853] = 12'h666;
rom[28854] = 12'h666;
rom[28855] = 12'h777;
rom[28856] = 12'h777;
rom[28857] = 12'h888;
rom[28858] = 12'h888;
rom[28859] = 12'h888;
rom[28860] = 12'h888;
rom[28861] = 12'h888;
rom[28862] = 12'h777;
rom[28863] = 12'h777;
rom[28864] = 12'h666;
rom[28865] = 12'h666;
rom[28866] = 12'h666;
rom[28867] = 12'h555;
rom[28868] = 12'h555;
rom[28869] = 12'h555;
rom[28870] = 12'h555;
rom[28871] = 12'h555;
rom[28872] = 12'h555;
rom[28873] = 12'h444;
rom[28874] = 12'h444;
rom[28875] = 12'h444;
rom[28876] = 12'h444;
rom[28877] = 12'h444;
rom[28878] = 12'h444;
rom[28879] = 12'h333;
rom[28880] = 12'h333;
rom[28881] = 12'h333;
rom[28882] = 12'h333;
rom[28883] = 12'h222;
rom[28884] = 12'h222;
rom[28885] = 12'h222;
rom[28886] = 12'h222;
rom[28887] = 12'h222;
rom[28888] = 12'h222;
rom[28889] = 12'h222;
rom[28890] = 12'h222;
rom[28891] = 12'h222;
rom[28892] = 12'h222;
rom[28893] = 12'h222;
rom[28894] = 12'h111;
rom[28895] = 12'h111;
rom[28896] = 12'h111;
rom[28897] = 12'h111;
rom[28898] = 12'h111;
rom[28899] = 12'h111;
rom[28900] = 12'h  0;
rom[28901] = 12'h  0;
rom[28902] = 12'h  0;
rom[28903] = 12'h  0;
rom[28904] = 12'h  0;
rom[28905] = 12'h  0;
rom[28906] = 12'h  0;
rom[28907] = 12'h  0;
rom[28908] = 12'h  0;
rom[28909] = 12'h  0;
rom[28910] = 12'h  0;
rom[28911] = 12'h  0;
rom[28912] = 12'h  0;
rom[28913] = 12'h  0;
rom[28914] = 12'h  0;
rom[28915] = 12'h  0;
rom[28916] = 12'h  0;
rom[28917] = 12'h  0;
rom[28918] = 12'h  0;
rom[28919] = 12'h  0;
rom[28920] = 12'h  0;
rom[28921] = 12'h  0;
rom[28922] = 12'h100;
rom[28923] = 12'h100;
rom[28924] = 12'h100;
rom[28925] = 12'h100;
rom[28926] = 12'h200;
rom[28927] = 12'h200;
rom[28928] = 12'h200;
rom[28929] = 12'h200;
rom[28930] = 12'h310;
rom[28931] = 12'h410;
rom[28932] = 12'h410;
rom[28933] = 12'h520;
rom[28934] = 12'h620;
rom[28935] = 12'h720;
rom[28936] = 12'h820;
rom[28937] = 12'h830;
rom[28938] = 12'h930;
rom[28939] = 12'ha30;
rom[28940] = 12'ha30;
rom[28941] = 12'hb40;
rom[28942] = 12'hb40;
rom[28943] = 12'hb40;
rom[28944] = 12'hb30;
rom[28945] = 12'hc30;
rom[28946] = 12'hc30;
rom[28947] = 12'hc30;
rom[28948] = 12'hc30;
rom[28949] = 12'hc30;
rom[28950] = 12'hb30;
rom[28951] = 12'hb20;
rom[28952] = 12'hb20;
rom[28953] = 12'hb20;
rom[28954] = 12'ha20;
rom[28955] = 12'ha20;
rom[28956] = 12'ha10;
rom[28957] = 12'ha10;
rom[28958] = 12'h910;
rom[28959] = 12'h910;
rom[28960] = 12'h710;
rom[28961] = 12'h610;
rom[28962] = 12'h610;
rom[28963] = 12'h600;
rom[28964] = 12'h500;
rom[28965] = 12'h500;
rom[28966] = 12'h500;
rom[28967] = 12'h400;
rom[28968] = 12'h300;
rom[28969] = 12'h300;
rom[28970] = 12'h200;
rom[28971] = 12'h200;
rom[28972] = 12'h200;
rom[28973] = 12'h100;
rom[28974] = 12'h100;
rom[28975] = 12'h100;
rom[28976] = 12'h100;
rom[28977] = 12'h100;
rom[28978] = 12'h100;
rom[28979] = 12'h100;
rom[28980] = 12'h100;
rom[28981] = 12'h100;
rom[28982] = 12'h100;
rom[28983] = 12'h100;
rom[28984] = 12'h211;
rom[28985] = 12'h211;
rom[28986] = 12'h211;
rom[28987] = 12'h111;
rom[28988] = 12'h  0;
rom[28989] = 12'h  0;
rom[28990] = 12'h111;
rom[28991] = 12'h111;
rom[28992] = 12'h111;
rom[28993] = 12'h111;
rom[28994] = 12'h111;
rom[28995] = 12'h111;
rom[28996] = 12'h111;
rom[28997] = 12'h111;
rom[28998] = 12'h111;
rom[28999] = 12'h222;
rom[29000] = 12'h222;
rom[29001] = 12'h222;
rom[29002] = 12'h333;
rom[29003] = 12'h333;
rom[29004] = 12'h444;
rom[29005] = 12'h666;
rom[29006] = 12'h777;
rom[29007] = 12'h777;
rom[29008] = 12'h777;
rom[29009] = 12'h888;
rom[29010] = 12'h888;
rom[29011] = 12'h888;
rom[29012] = 12'h888;
rom[29013] = 12'h777;
rom[29014] = 12'h777;
rom[29015] = 12'h666;
rom[29016] = 12'h777;
rom[29017] = 12'h777;
rom[29018] = 12'h777;
rom[29019] = 12'h777;
rom[29020] = 12'h777;
rom[29021] = 12'h777;
rom[29022] = 12'h666;
rom[29023] = 12'h666;
rom[29024] = 12'h666;
rom[29025] = 12'h666;
rom[29026] = 12'h666;
rom[29027] = 12'h777;
rom[29028] = 12'h777;
rom[29029] = 12'h777;
rom[29030] = 12'h777;
rom[29031] = 12'h777;
rom[29032] = 12'h777;
rom[29033] = 12'h777;
rom[29034] = 12'h666;
rom[29035] = 12'h666;
rom[29036] = 12'h666;
rom[29037] = 12'h555;
rom[29038] = 12'h555;
rom[29039] = 12'h555;
rom[29040] = 12'h444;
rom[29041] = 12'h444;
rom[29042] = 12'h333;
rom[29043] = 12'h333;
rom[29044] = 12'h222;
rom[29045] = 12'h222;
rom[29046] = 12'h222;
rom[29047] = 12'h111;
rom[29048] = 12'h111;
rom[29049] = 12'h111;
rom[29050] = 12'h111;
rom[29051] = 12'h111;
rom[29052] = 12'h  0;
rom[29053] = 12'h  0;
rom[29054] = 12'h  0;
rom[29055] = 12'h111;
rom[29056] = 12'h  0;
rom[29057] = 12'h  0;
rom[29058] = 12'h  0;
rom[29059] = 12'h  0;
rom[29060] = 12'h  0;
rom[29061] = 12'h  0;
rom[29062] = 12'h  0;
rom[29063] = 12'h  0;
rom[29064] = 12'h  0;
rom[29065] = 12'h  0;
rom[29066] = 12'h  0;
rom[29067] = 12'h  0;
rom[29068] = 12'h  0;
rom[29069] = 12'h  0;
rom[29070] = 12'h  0;
rom[29071] = 12'h  0;
rom[29072] = 12'h  0;
rom[29073] = 12'h  0;
rom[29074] = 12'h  0;
rom[29075] = 12'h  0;
rom[29076] = 12'h  0;
rom[29077] = 12'h  0;
rom[29078] = 12'h  0;
rom[29079] = 12'h  0;
rom[29080] = 12'h  0;
rom[29081] = 12'h  0;
rom[29082] = 12'h  0;
rom[29083] = 12'h  0;
rom[29084] = 12'h  0;
rom[29085] = 12'h  0;
rom[29086] = 12'h  0;
rom[29087] = 12'h111;
rom[29088] = 12'h  0;
rom[29089] = 12'h111;
rom[29090] = 12'h111;
rom[29091] = 12'h111;
rom[29092] = 12'h111;
rom[29093] = 12'h222;
rom[29094] = 12'h222;
rom[29095] = 12'h222;
rom[29096] = 12'h222;
rom[29097] = 12'h333;
rom[29098] = 12'h333;
rom[29099] = 12'h333;
rom[29100] = 12'h333;
rom[29101] = 12'h333;
rom[29102] = 12'h444;
rom[29103] = 12'h666;
rom[29104] = 12'h666;
rom[29105] = 12'h555;
rom[29106] = 12'h555;
rom[29107] = 12'h666;
rom[29108] = 12'h666;
rom[29109] = 12'h666;
rom[29110] = 12'h777;
rom[29111] = 12'h777;
rom[29112] = 12'h888;
rom[29113] = 12'h999;
rom[29114] = 12'h999;
rom[29115] = 12'hbbb;
rom[29116] = 12'hccc;
rom[29117] = 12'hddd;
rom[29118] = 12'heee;
rom[29119] = 12'hfee;
rom[29120] = 12'hffe;
rom[29121] = 12'hffe;
rom[29122] = 12'heed;
rom[29123] = 12'hcba;
rom[29124] = 12'h877;
rom[29125] = 12'h543;
rom[29126] = 12'h321;
rom[29127] = 12'h210;
rom[29128] = 12'h311;
rom[29129] = 12'h310;
rom[29130] = 12'h310;
rom[29131] = 12'h300;
rom[29132] = 12'h300;
rom[29133] = 12'h300;
rom[29134] = 12'h300;
rom[29135] = 12'h300;
rom[29136] = 12'h300;
rom[29137] = 12'h400;
rom[29138] = 12'h400;
rom[29139] = 12'h410;
rom[29140] = 12'h510;
rom[29141] = 12'h610;
rom[29142] = 12'h710;
rom[29143] = 12'h710;
rom[29144] = 12'h820;
rom[29145] = 12'h920;
rom[29146] = 12'ha20;
rom[29147] = 12'hb30;
rom[29148] = 12'hb30;
rom[29149] = 12'hc40;
rom[29150] = 12'hc40;
rom[29151] = 12'hc40;
rom[29152] = 12'hc40;
rom[29153] = 12'hb40;
rom[29154] = 12'hb40;
rom[29155] = 12'ha40;
rom[29156] = 12'h940;
rom[29157] = 12'h940;
rom[29158] = 12'ha61;
rom[29159] = 12'hb72;
rom[29160] = 12'hb62;
rom[29161] = 12'ha51;
rom[29162] = 12'h940;
rom[29163] = 12'h840;
rom[29164] = 12'h840;
rom[29165] = 12'h740;
rom[29166] = 12'h740;
rom[29167] = 12'h640;
rom[29168] = 12'h641;
rom[29169] = 12'h641;
rom[29170] = 12'h642;
rom[29171] = 12'h642;
rom[29172] = 12'h643;
rom[29173] = 12'h653;
rom[29174] = 12'h654;
rom[29175] = 12'h654;
rom[29176] = 12'h765;
rom[29177] = 12'h766;
rom[29178] = 12'h777;
rom[29179] = 12'h787;
rom[29180] = 12'h787;
rom[29181] = 12'h887;
rom[29182] = 12'h888;
rom[29183] = 12'h888;
rom[29184] = 12'h999;
rom[29185] = 12'h999;
rom[29186] = 12'h999;
rom[29187] = 12'h999;
rom[29188] = 12'h888;
rom[29189] = 12'h888;
rom[29190] = 12'h888;
rom[29191] = 12'h888;
rom[29192] = 12'h888;
rom[29193] = 12'h999;
rom[29194] = 12'h999;
rom[29195] = 12'haaa;
rom[29196] = 12'haaa;
rom[29197] = 12'haaa;
rom[29198] = 12'haaa;
rom[29199] = 12'haaa;
rom[29200] = 12'h666;
rom[29201] = 12'h666;
rom[29202] = 12'h666;
rom[29203] = 12'h555;
rom[29204] = 12'h555;
rom[29205] = 12'h555;
rom[29206] = 12'h555;
rom[29207] = 12'h555;
rom[29208] = 12'h666;
rom[29209] = 12'h666;
rom[29210] = 12'h666;
rom[29211] = 12'h666;
rom[29212] = 12'h666;
rom[29213] = 12'h666;
rom[29214] = 12'h666;
rom[29215] = 12'h666;
rom[29216] = 12'h666;
rom[29217] = 12'h666;
rom[29218] = 12'h666;
rom[29219] = 12'h666;
rom[29220] = 12'h666;
rom[29221] = 12'h666;
rom[29222] = 12'h666;
rom[29223] = 12'h666;
rom[29224] = 12'h666;
rom[29225] = 12'h666;
rom[29226] = 12'h666;
rom[29227] = 12'h777;
rom[29228] = 12'h777;
rom[29229] = 12'h777;
rom[29230] = 12'h777;
rom[29231] = 12'h777;
rom[29232] = 12'h777;
rom[29233] = 12'h777;
rom[29234] = 12'h777;
rom[29235] = 12'h888;
rom[29236] = 12'h888;
rom[29237] = 12'h888;
rom[29238] = 12'h888;
rom[29239] = 12'h999;
rom[29240] = 12'h888;
rom[29241] = 12'h888;
rom[29242] = 12'h888;
rom[29243] = 12'h888;
rom[29244] = 12'h777;
rom[29245] = 12'h777;
rom[29246] = 12'h777;
rom[29247] = 12'h777;
rom[29248] = 12'h777;
rom[29249] = 12'h666;
rom[29250] = 12'h666;
rom[29251] = 12'h666;
rom[29252] = 12'h666;
rom[29253] = 12'h666;
rom[29254] = 12'h666;
rom[29255] = 12'h777;
rom[29256] = 12'h777;
rom[29257] = 12'h777;
rom[29258] = 12'h888;
rom[29259] = 12'h888;
rom[29260] = 12'h888;
rom[29261] = 12'h888;
rom[29262] = 12'h888;
rom[29263] = 12'h777;
rom[29264] = 12'h666;
rom[29265] = 12'h666;
rom[29266] = 12'h666;
rom[29267] = 12'h666;
rom[29268] = 12'h555;
rom[29269] = 12'h555;
rom[29270] = 12'h555;
rom[29271] = 12'h555;
rom[29272] = 12'h555;
rom[29273] = 12'h444;
rom[29274] = 12'h444;
rom[29275] = 12'h444;
rom[29276] = 12'h444;
rom[29277] = 12'h444;
rom[29278] = 12'h444;
rom[29279] = 12'h333;
rom[29280] = 12'h333;
rom[29281] = 12'h333;
rom[29282] = 12'h333;
rom[29283] = 12'h333;
rom[29284] = 12'h222;
rom[29285] = 12'h222;
rom[29286] = 12'h222;
rom[29287] = 12'h222;
rom[29288] = 12'h222;
rom[29289] = 12'h222;
rom[29290] = 12'h222;
rom[29291] = 12'h222;
rom[29292] = 12'h222;
rom[29293] = 12'h111;
rom[29294] = 12'h111;
rom[29295] = 12'h111;
rom[29296] = 12'h  0;
rom[29297] = 12'h  0;
rom[29298] = 12'h  0;
rom[29299] = 12'h  0;
rom[29300] = 12'h  0;
rom[29301] = 12'h  0;
rom[29302] = 12'h  0;
rom[29303] = 12'h  0;
rom[29304] = 12'h  0;
rom[29305] = 12'h  0;
rom[29306] = 12'h  0;
rom[29307] = 12'h  0;
rom[29308] = 12'h  0;
rom[29309] = 12'h  0;
rom[29310] = 12'h  0;
rom[29311] = 12'h  0;
rom[29312] = 12'h  0;
rom[29313] = 12'h  0;
rom[29314] = 12'h  0;
rom[29315] = 12'h  0;
rom[29316] = 12'h  0;
rom[29317] = 12'h  0;
rom[29318] = 12'h  0;
rom[29319] = 12'h  0;
rom[29320] = 12'h  0;
rom[29321] = 12'h  0;
rom[29322] = 12'h  0;
rom[29323] = 12'h100;
rom[29324] = 12'h100;
rom[29325] = 12'h100;
rom[29326] = 12'h100;
rom[29327] = 12'h100;
rom[29328] = 12'h200;
rom[29329] = 12'h200;
rom[29330] = 12'h200;
rom[29331] = 12'h310;
rom[29332] = 12'h410;
rom[29333] = 12'h410;
rom[29334] = 12'h510;
rom[29335] = 12'h620;
rom[29336] = 12'h720;
rom[29337] = 12'h720;
rom[29338] = 12'h820;
rom[29339] = 12'h930;
rom[29340] = 12'h930;
rom[29341] = 12'h930;
rom[29342] = 12'ha30;
rom[29343] = 12'ha30;
rom[29344] = 12'ha30;
rom[29345] = 12'ha30;
rom[29346] = 12'ha30;
rom[29347] = 12'ha30;
rom[29348] = 12'ha30;
rom[29349] = 12'ha20;
rom[29350] = 12'ha20;
rom[29351] = 12'ha20;
rom[29352] = 12'ha20;
rom[29353] = 12'h920;
rom[29354] = 12'h910;
rom[29355] = 12'h910;
rom[29356] = 12'h910;
rom[29357] = 12'h810;
rom[29358] = 12'h810;
rom[29359] = 12'h810;
rom[29360] = 12'h600;
rom[29361] = 12'h500;
rom[29362] = 12'h500;
rom[29363] = 12'h500;
rom[29364] = 12'h400;
rom[29365] = 12'h400;
rom[29366] = 12'h400;
rom[29367] = 12'h300;
rom[29368] = 12'h200;
rom[29369] = 12'h200;
rom[29370] = 12'h200;
rom[29371] = 12'h100;
rom[29372] = 12'h100;
rom[29373] = 12'h100;
rom[29374] = 12'h100;
rom[29375] = 12'h100;
rom[29376] = 12'h100;
rom[29377] = 12'h100;
rom[29378] = 12'h100;
rom[29379] = 12'h100;
rom[29380] = 12'h100;
rom[29381] = 12'h100;
rom[29382] = 12'h100;
rom[29383] = 12'h100;
rom[29384] = 12'h211;
rom[29385] = 12'h211;
rom[29386] = 12'h111;
rom[29387] = 12'h100;
rom[29388] = 12'h  0;
rom[29389] = 12'h111;
rom[29390] = 12'h111;
rom[29391] = 12'h  0;
rom[29392] = 12'h111;
rom[29393] = 12'h111;
rom[29394] = 12'h111;
rom[29395] = 12'h111;
rom[29396] = 12'h111;
rom[29397] = 12'h111;
rom[29398] = 12'h222;
rom[29399] = 12'h222;
rom[29400] = 12'h222;
rom[29401] = 12'h222;
rom[29402] = 12'h333;
rom[29403] = 12'h333;
rom[29404] = 12'h444;
rom[29405] = 12'h666;
rom[29406] = 12'h777;
rom[29407] = 12'h777;
rom[29408] = 12'h777;
rom[29409] = 12'h888;
rom[29410] = 12'h888;
rom[29411] = 12'h888;
rom[29412] = 12'h777;
rom[29413] = 12'h777;
rom[29414] = 12'h777;
rom[29415] = 12'h666;
rom[29416] = 12'h777;
rom[29417] = 12'h777;
rom[29418] = 12'h777;
rom[29419] = 12'h777;
rom[29420] = 12'h777;
rom[29421] = 12'h666;
rom[29422] = 12'h666;
rom[29423] = 12'h666;
rom[29424] = 12'h666;
rom[29425] = 12'h666;
rom[29426] = 12'h666;
rom[29427] = 12'h666;
rom[29428] = 12'h777;
rom[29429] = 12'h777;
rom[29430] = 12'h777;
rom[29431] = 12'h777;
rom[29432] = 12'h777;
rom[29433] = 12'h777;
rom[29434] = 12'h666;
rom[29435] = 12'h666;
rom[29436] = 12'h666;
rom[29437] = 12'h555;
rom[29438] = 12'h555;
rom[29439] = 12'h444;
rom[29440] = 12'h444;
rom[29441] = 12'h333;
rom[29442] = 12'h333;
rom[29443] = 12'h222;
rom[29444] = 12'h222;
rom[29445] = 12'h222;
rom[29446] = 12'h222;
rom[29447] = 12'h111;
rom[29448] = 12'h111;
rom[29449] = 12'h111;
rom[29450] = 12'h111;
rom[29451] = 12'h111;
rom[29452] = 12'h  0;
rom[29453] = 12'h  0;
rom[29454] = 12'h  0;
rom[29455] = 12'h111;
rom[29456] = 12'h  0;
rom[29457] = 12'h  0;
rom[29458] = 12'h  0;
rom[29459] = 12'h  0;
rom[29460] = 12'h  0;
rom[29461] = 12'h  0;
rom[29462] = 12'h  0;
rom[29463] = 12'h  0;
rom[29464] = 12'h  0;
rom[29465] = 12'h  0;
rom[29466] = 12'h  0;
rom[29467] = 12'h  0;
rom[29468] = 12'h  0;
rom[29469] = 12'h  0;
rom[29470] = 12'h  0;
rom[29471] = 12'h  0;
rom[29472] = 12'h  0;
rom[29473] = 12'h  0;
rom[29474] = 12'h  0;
rom[29475] = 12'h  0;
rom[29476] = 12'h  0;
rom[29477] = 12'h  0;
rom[29478] = 12'h  0;
rom[29479] = 12'h  0;
rom[29480] = 12'h  0;
rom[29481] = 12'h  0;
rom[29482] = 12'h  0;
rom[29483] = 12'h  0;
rom[29484] = 12'h  0;
rom[29485] = 12'h  0;
rom[29486] = 12'h  0;
rom[29487] = 12'h111;
rom[29488] = 12'h  0;
rom[29489] = 12'h111;
rom[29490] = 12'h111;
rom[29491] = 12'h111;
rom[29492] = 12'h111;
rom[29493] = 12'h222;
rom[29494] = 12'h222;
rom[29495] = 12'h222;
rom[29496] = 12'h333;
rom[29497] = 12'h333;
rom[29498] = 12'h333;
rom[29499] = 12'h333;
rom[29500] = 12'h333;
rom[29501] = 12'h333;
rom[29502] = 12'h555;
rom[29503] = 12'h666;
rom[29504] = 12'h666;
rom[29505] = 12'h666;
rom[29506] = 12'h666;
rom[29507] = 12'h666;
rom[29508] = 12'h777;
rom[29509] = 12'h777;
rom[29510] = 12'h888;
rom[29511] = 12'h888;
rom[29512] = 12'h999;
rom[29513] = 12'haaa;
rom[29514] = 12'hccc;
rom[29515] = 12'hccc;
rom[29516] = 12'hddd;
rom[29517] = 12'heee;
rom[29518] = 12'hfff;
rom[29519] = 12'hfff;
rom[29520] = 12'hffe;
rom[29521] = 12'hddc;
rom[29522] = 12'ha99;
rom[29523] = 12'h655;
rom[29524] = 12'h332;
rom[29525] = 12'h211;
rom[29526] = 12'h211;
rom[29527] = 12'h311;
rom[29528] = 12'h210;
rom[29529] = 12'h210;
rom[29530] = 12'h200;
rom[29531] = 12'h200;
rom[29532] = 12'h300;
rom[29533] = 12'h300;
rom[29534] = 12'h300;
rom[29535] = 12'h300;
rom[29536] = 12'h300;
rom[29537] = 12'h300;
rom[29538] = 12'h400;
rom[29539] = 12'h400;
rom[29540] = 12'h500;
rom[29541] = 12'h510;
rom[29542] = 12'h610;
rom[29543] = 12'h710;
rom[29544] = 12'h820;
rom[29545] = 12'h920;
rom[29546] = 12'ha20;
rom[29547] = 12'hb30;
rom[29548] = 12'hc30;
rom[29549] = 12'hd40;
rom[29550] = 12'hd40;
rom[29551] = 12'hd40;
rom[29552] = 12'hc40;
rom[29553] = 12'hc40;
rom[29554] = 12'hb40;
rom[29555] = 12'hb40;
rom[29556] = 12'ha40;
rom[29557] = 12'ha50;
rom[29558] = 12'hb61;
rom[29559] = 12'hb72;
rom[29560] = 12'hb61;
rom[29561] = 12'h951;
rom[29562] = 12'h840;
rom[29563] = 12'h840;
rom[29564] = 12'h840;
rom[29565] = 12'h740;
rom[29566] = 12'h740;
rom[29567] = 12'h740;
rom[29568] = 12'h641;
rom[29569] = 12'h641;
rom[29570] = 12'h642;
rom[29571] = 12'h642;
rom[29572] = 12'h642;
rom[29573] = 12'h643;
rom[29574] = 12'h654;
rom[29575] = 12'h654;
rom[29576] = 12'h665;
rom[29577] = 12'h666;
rom[29578] = 12'h776;
rom[29579] = 12'h777;
rom[29580] = 12'h887;
rom[29581] = 12'h888;
rom[29582] = 12'h888;
rom[29583] = 12'h888;
rom[29584] = 12'h999;
rom[29585] = 12'h999;
rom[29586] = 12'h999;
rom[29587] = 12'h999;
rom[29588] = 12'h999;
rom[29589] = 12'h888;
rom[29590] = 12'h888;
rom[29591] = 12'h888;
rom[29592] = 12'h888;
rom[29593] = 12'h999;
rom[29594] = 12'h999;
rom[29595] = 12'haaa;
rom[29596] = 12'haaa;
rom[29597] = 12'haaa;
rom[29598] = 12'haaa;
rom[29599] = 12'haaa;
rom[29600] = 12'h666;
rom[29601] = 12'h666;
rom[29602] = 12'h666;
rom[29603] = 12'h555;
rom[29604] = 12'h555;
rom[29605] = 12'h555;
rom[29606] = 12'h555;
rom[29607] = 12'h666;
rom[29608] = 12'h666;
rom[29609] = 12'h666;
rom[29610] = 12'h666;
rom[29611] = 12'h666;
rom[29612] = 12'h666;
rom[29613] = 12'h666;
rom[29614] = 12'h666;
rom[29615] = 12'h666;
rom[29616] = 12'h666;
rom[29617] = 12'h666;
rom[29618] = 12'h666;
rom[29619] = 12'h666;
rom[29620] = 12'h666;
rom[29621] = 12'h666;
rom[29622] = 12'h666;
rom[29623] = 12'h666;
rom[29624] = 12'h666;
rom[29625] = 12'h666;
rom[29626] = 12'h666;
rom[29627] = 12'h666;
rom[29628] = 12'h777;
rom[29629] = 12'h777;
rom[29630] = 12'h777;
rom[29631] = 12'h777;
rom[29632] = 12'h777;
rom[29633] = 12'h777;
rom[29634] = 12'h888;
rom[29635] = 12'h888;
rom[29636] = 12'h888;
rom[29637] = 12'h888;
rom[29638] = 12'h888;
rom[29639] = 12'h999;
rom[29640] = 12'h888;
rom[29641] = 12'h888;
rom[29642] = 12'h888;
rom[29643] = 12'h888;
rom[29644] = 12'h777;
rom[29645] = 12'h777;
rom[29646] = 12'h777;
rom[29647] = 12'h666;
rom[29648] = 12'h666;
rom[29649] = 12'h666;
rom[29650] = 12'h666;
rom[29651] = 12'h666;
rom[29652] = 12'h666;
rom[29653] = 12'h666;
rom[29654] = 12'h666;
rom[29655] = 12'h666;
rom[29656] = 12'h777;
rom[29657] = 12'h777;
rom[29658] = 12'h888;
rom[29659] = 12'h888;
rom[29660] = 12'h888;
rom[29661] = 12'h888;
rom[29662] = 12'h888;
rom[29663] = 12'h888;
rom[29664] = 12'h777;
rom[29665] = 12'h777;
rom[29666] = 12'h666;
rom[29667] = 12'h666;
rom[29668] = 12'h555;
rom[29669] = 12'h555;
rom[29670] = 12'h555;
rom[29671] = 12'h555;
rom[29672] = 12'h555;
rom[29673] = 12'h444;
rom[29674] = 12'h444;
rom[29675] = 12'h444;
rom[29676] = 12'h444;
rom[29677] = 12'h444;
rom[29678] = 12'h444;
rom[29679] = 12'h333;
rom[29680] = 12'h333;
rom[29681] = 12'h333;
rom[29682] = 12'h333;
rom[29683] = 12'h333;
rom[29684] = 12'h222;
rom[29685] = 12'h222;
rom[29686] = 12'h222;
rom[29687] = 12'h222;
rom[29688] = 12'h222;
rom[29689] = 12'h222;
rom[29690] = 12'h222;
rom[29691] = 12'h222;
rom[29692] = 12'h222;
rom[29693] = 12'h111;
rom[29694] = 12'h111;
rom[29695] = 12'h111;
rom[29696] = 12'h  0;
rom[29697] = 12'h  0;
rom[29698] = 12'h  0;
rom[29699] = 12'h  0;
rom[29700] = 12'h  0;
rom[29701] = 12'h  0;
rom[29702] = 12'h  0;
rom[29703] = 12'h  0;
rom[29704] = 12'h  0;
rom[29705] = 12'h  0;
rom[29706] = 12'h  0;
rom[29707] = 12'h  0;
rom[29708] = 12'h  0;
rom[29709] = 12'h  0;
rom[29710] = 12'h  0;
rom[29711] = 12'h  0;
rom[29712] = 12'h  0;
rom[29713] = 12'h  0;
rom[29714] = 12'h  0;
rom[29715] = 12'h  0;
rom[29716] = 12'h  0;
rom[29717] = 12'h  0;
rom[29718] = 12'h  0;
rom[29719] = 12'h  0;
rom[29720] = 12'h  0;
rom[29721] = 12'h  0;
rom[29722] = 12'h  0;
rom[29723] = 12'h  0;
rom[29724] = 12'h  0;
rom[29725] = 12'h100;
rom[29726] = 12'h100;
rom[29727] = 12'h100;
rom[29728] = 12'h100;
rom[29729] = 12'h200;
rom[29730] = 12'h200;
rom[29731] = 12'h200;
rom[29732] = 12'h300;
rom[29733] = 12'h410;
rom[29734] = 12'h510;
rom[29735] = 12'h510;
rom[29736] = 12'h610;
rom[29737] = 12'h610;
rom[29738] = 12'h720;
rom[29739] = 12'h720;
rom[29740] = 12'h820;
rom[29741] = 12'h820;
rom[29742] = 12'h820;
rom[29743] = 12'h820;
rom[29744] = 12'h820;
rom[29745] = 12'h920;
rom[29746] = 12'h920;
rom[29747] = 12'h920;
rom[29748] = 12'h920;
rom[29749] = 12'h920;
rom[29750] = 12'h920;
rom[29751] = 12'h820;
rom[29752] = 12'h810;
rom[29753] = 12'h810;
rom[29754] = 12'h810;
rom[29755] = 12'h710;
rom[29756] = 12'h710;
rom[29757] = 12'h710;
rom[29758] = 12'h700;
rom[29759] = 12'h600;
rom[29760] = 12'h500;
rom[29761] = 12'h400;
rom[29762] = 12'h400;
rom[29763] = 12'h400;
rom[29764] = 12'h300;
rom[29765] = 12'h300;
rom[29766] = 12'h300;
rom[29767] = 12'h200;
rom[29768] = 12'h200;
rom[29769] = 12'h200;
rom[29770] = 12'h100;
rom[29771] = 12'h100;
rom[29772] = 12'h100;
rom[29773] = 12'h100;
rom[29774] = 12'h  0;
rom[29775] = 12'h  0;
rom[29776] = 12'h100;
rom[29777] = 12'h100;
rom[29778] = 12'h100;
rom[29779] = 12'h100;
rom[29780] = 12'h100;
rom[29781] = 12'h100;
rom[29782] = 12'h100;
rom[29783] = 12'h111;
rom[29784] = 12'h211;
rom[29785] = 12'h111;
rom[29786] = 12'h  0;
rom[29787] = 12'h  0;
rom[29788] = 12'h  0;
rom[29789] = 12'h111;
rom[29790] = 12'h110;
rom[29791] = 12'h  0;
rom[29792] = 12'h  0;
rom[29793] = 12'h  0;
rom[29794] = 12'h111;
rom[29795] = 12'h111;
rom[29796] = 12'h111;
rom[29797] = 12'h111;
rom[29798] = 12'h222;
rom[29799] = 12'h222;
rom[29800] = 12'h222;
rom[29801] = 12'h222;
rom[29802] = 12'h222;
rom[29803] = 12'h333;
rom[29804] = 12'h444;
rom[29805] = 12'h555;
rom[29806] = 12'h666;
rom[29807] = 12'h777;
rom[29808] = 12'h777;
rom[29809] = 12'h888;
rom[29810] = 12'h888;
rom[29811] = 12'h777;
rom[29812] = 12'h777;
rom[29813] = 12'h777;
rom[29814] = 12'h777;
rom[29815] = 12'h666;
rom[29816] = 12'h666;
rom[29817] = 12'h666;
rom[29818] = 12'h666;
rom[29819] = 12'h666;
rom[29820] = 12'h666;
rom[29821] = 12'h666;
rom[29822] = 12'h666;
rom[29823] = 12'h666;
rom[29824] = 12'h666;
rom[29825] = 12'h666;
rom[29826] = 12'h666;
rom[29827] = 12'h666;
rom[29828] = 12'h666;
rom[29829] = 12'h777;
rom[29830] = 12'h777;
rom[29831] = 12'h777;
rom[29832] = 12'h777;
rom[29833] = 12'h666;
rom[29834] = 12'h666;
rom[29835] = 12'h666;
rom[29836] = 12'h666;
rom[29837] = 12'h555;
rom[29838] = 12'h555;
rom[29839] = 12'h444;
rom[29840] = 12'h333;
rom[29841] = 12'h333;
rom[29842] = 12'h222;
rom[29843] = 12'h222;
rom[29844] = 12'h222;
rom[29845] = 12'h222;
rom[29846] = 12'h222;
rom[29847] = 12'h222;
rom[29848] = 12'h111;
rom[29849] = 12'h111;
rom[29850] = 12'h111;
rom[29851] = 12'h111;
rom[29852] = 12'h  0;
rom[29853] = 12'h  0;
rom[29854] = 12'h  0;
rom[29855] = 12'h111;
rom[29856] = 12'h  0;
rom[29857] = 12'h  0;
rom[29858] = 12'h  0;
rom[29859] = 12'h  0;
rom[29860] = 12'h  0;
rom[29861] = 12'h  0;
rom[29862] = 12'h  0;
rom[29863] = 12'h  0;
rom[29864] = 12'h  0;
rom[29865] = 12'h  0;
rom[29866] = 12'h  0;
rom[29867] = 12'h  0;
rom[29868] = 12'h  0;
rom[29869] = 12'h  0;
rom[29870] = 12'h  0;
rom[29871] = 12'h  0;
rom[29872] = 12'h  0;
rom[29873] = 12'h  0;
rom[29874] = 12'h  0;
rom[29875] = 12'h  0;
rom[29876] = 12'h  0;
rom[29877] = 12'h  0;
rom[29878] = 12'h  0;
rom[29879] = 12'h  0;
rom[29880] = 12'h  0;
rom[29881] = 12'h  0;
rom[29882] = 12'h  0;
rom[29883] = 12'h  0;
rom[29884] = 12'h  0;
rom[29885] = 12'h  0;
rom[29886] = 12'h  0;
rom[29887] = 12'h111;
rom[29888] = 12'h111;
rom[29889] = 12'h111;
rom[29890] = 12'h222;
rom[29891] = 12'h111;
rom[29892] = 12'h111;
rom[29893] = 12'h222;
rom[29894] = 12'h222;
rom[29895] = 12'h222;
rom[29896] = 12'h333;
rom[29897] = 12'h333;
rom[29898] = 12'h333;
rom[29899] = 12'h333;
rom[29900] = 12'h444;
rom[29901] = 12'h444;
rom[29902] = 12'h555;
rom[29903] = 12'h666;
rom[29904] = 12'h666;
rom[29905] = 12'h666;
rom[29906] = 12'h777;
rom[29907] = 12'h777;
rom[29908] = 12'h888;
rom[29909] = 12'h888;
rom[29910] = 12'h999;
rom[29911] = 12'ha99;
rom[29912] = 12'haaa;
rom[29913] = 12'hcbb;
rom[29914] = 12'hddd;
rom[29915] = 12'heed;
rom[29916] = 12'hfee;
rom[29917] = 12'hfff;
rom[29918] = 12'hfff;
rom[29919] = 12'hfff;
rom[29920] = 12'hbba;
rom[29921] = 12'h888;
rom[29922] = 12'h544;
rom[29923] = 12'h221;
rom[29924] = 12'h110;
rom[29925] = 12'h110;
rom[29926] = 12'h211;
rom[29927] = 12'h211;
rom[29928] = 12'h210;
rom[29929] = 12'h200;
rom[29930] = 12'h200;
rom[29931] = 12'h200;
rom[29932] = 12'h200;
rom[29933] = 12'h200;
rom[29934] = 12'h300;
rom[29935] = 12'h300;
rom[29936] = 12'h300;
rom[29937] = 12'h300;
rom[29938] = 12'h300;
rom[29939] = 12'h400;
rom[29940] = 12'h400;
rom[29941] = 12'h500;
rom[29942] = 12'h610;
rom[29943] = 12'h610;
rom[29944] = 12'h810;
rom[29945] = 12'h920;
rom[29946] = 12'ha20;
rom[29947] = 12'hb30;
rom[29948] = 12'hc30;
rom[29949] = 12'hd40;
rom[29950] = 12'hd40;
rom[29951] = 12'hd40;
rom[29952] = 12'hd40;
rom[29953] = 12'hc40;
rom[29954] = 12'hc40;
rom[29955] = 12'hb50;
rom[29956] = 12'ha50;
rom[29957] = 12'hb60;
rom[29958] = 12'hb61;
rom[29959] = 12'hb72;
rom[29960] = 12'ha61;
rom[29961] = 12'h950;
rom[29962] = 12'h840;
rom[29963] = 12'h840;
rom[29964] = 12'h840;
rom[29965] = 12'h740;
rom[29966] = 12'h740;
rom[29967] = 12'h640;
rom[29968] = 12'h641;
rom[29969] = 12'h641;
rom[29970] = 12'h642;
rom[29971] = 12'h642;
rom[29972] = 12'h642;
rom[29973] = 12'h643;
rom[29974] = 12'h653;
rom[29975] = 12'h654;
rom[29976] = 12'h654;
rom[29977] = 12'h665;
rom[29978] = 12'h766;
rom[29979] = 12'h777;
rom[29980] = 12'h777;
rom[29981] = 12'h888;
rom[29982] = 12'h888;
rom[29983] = 12'h888;
rom[29984] = 12'h999;
rom[29985] = 12'h999;
rom[29986] = 12'h999;
rom[29987] = 12'h999;
rom[29988] = 12'h999;
rom[29989] = 12'h999;
rom[29990] = 12'h888;
rom[29991] = 12'h888;
rom[29992] = 12'h999;
rom[29993] = 12'h999;
rom[29994] = 12'h999;
rom[29995] = 12'haaa;
rom[29996] = 12'haaa;
rom[29997] = 12'haaa;
rom[29998] = 12'haaa;
rom[29999] = 12'haaa;
rom[30000] = 12'h666;
rom[30001] = 12'h666;
rom[30002] = 12'h666;
rom[30003] = 12'h666;
rom[30004] = 12'h666;
rom[30005] = 12'h666;
rom[30006] = 12'h666;
rom[30007] = 12'h666;
rom[30008] = 12'h666;
rom[30009] = 12'h666;
rom[30010] = 12'h666;
rom[30011] = 12'h666;
rom[30012] = 12'h666;
rom[30013] = 12'h666;
rom[30014] = 12'h666;
rom[30015] = 12'h666;
rom[30016] = 12'h666;
rom[30017] = 12'h666;
rom[30018] = 12'h666;
rom[30019] = 12'h666;
rom[30020] = 12'h666;
rom[30021] = 12'h666;
rom[30022] = 12'h666;
rom[30023] = 12'h666;
rom[30024] = 12'h666;
rom[30025] = 12'h666;
rom[30026] = 12'h666;
rom[30027] = 12'h666;
rom[30028] = 12'h777;
rom[30029] = 12'h777;
rom[30030] = 12'h777;
rom[30031] = 12'h777;
rom[30032] = 12'h777;
rom[30033] = 12'h888;
rom[30034] = 12'h888;
rom[30035] = 12'h888;
rom[30036] = 12'h888;
rom[30037] = 12'h888;
rom[30038] = 12'h888;
rom[30039] = 12'h999;
rom[30040] = 12'h999;
rom[30041] = 12'h888;
rom[30042] = 12'h888;
rom[30043] = 12'h888;
rom[30044] = 12'h777;
rom[30045] = 12'h777;
rom[30046] = 12'h777;
rom[30047] = 12'h666;
rom[30048] = 12'h666;
rom[30049] = 12'h666;
rom[30050] = 12'h666;
rom[30051] = 12'h666;
rom[30052] = 12'h666;
rom[30053] = 12'h666;
rom[30054] = 12'h666;
rom[30055] = 12'h666;
rom[30056] = 12'h777;
rom[30057] = 12'h777;
rom[30058] = 12'h777;
rom[30059] = 12'h888;
rom[30060] = 12'h888;
rom[30061] = 12'h888;
rom[30062] = 12'h888;
rom[30063] = 12'h888;
rom[30064] = 12'h888;
rom[30065] = 12'h777;
rom[30066] = 12'h777;
rom[30067] = 12'h666;
rom[30068] = 12'h666;
rom[30069] = 12'h555;
rom[30070] = 12'h555;
rom[30071] = 12'h555;
rom[30072] = 12'h555;
rom[30073] = 12'h444;
rom[30074] = 12'h444;
rom[30075] = 12'h444;
rom[30076] = 12'h444;
rom[30077] = 12'h444;
rom[30078] = 12'h444;
rom[30079] = 12'h333;
rom[30080] = 12'h333;
rom[30081] = 12'h333;
rom[30082] = 12'h333;
rom[30083] = 12'h333;
rom[30084] = 12'h333;
rom[30085] = 12'h333;
rom[30086] = 12'h222;
rom[30087] = 12'h222;
rom[30088] = 12'h222;
rom[30089] = 12'h222;
rom[30090] = 12'h222;
rom[30091] = 12'h222;
rom[30092] = 12'h222;
rom[30093] = 12'h111;
rom[30094] = 12'h111;
rom[30095] = 12'h  0;
rom[30096] = 12'h  0;
rom[30097] = 12'h  0;
rom[30098] = 12'h  0;
rom[30099] = 12'h  0;
rom[30100] = 12'h  0;
rom[30101] = 12'h  0;
rom[30102] = 12'h  0;
rom[30103] = 12'h  0;
rom[30104] = 12'h  0;
rom[30105] = 12'h  0;
rom[30106] = 12'h  0;
rom[30107] = 12'h  0;
rom[30108] = 12'h  0;
rom[30109] = 12'h  0;
rom[30110] = 12'h  0;
rom[30111] = 12'h  0;
rom[30112] = 12'h  0;
rom[30113] = 12'h  0;
rom[30114] = 12'h  0;
rom[30115] = 12'h  0;
rom[30116] = 12'h  0;
rom[30117] = 12'h  0;
rom[30118] = 12'h  0;
rom[30119] = 12'h  0;
rom[30120] = 12'h  0;
rom[30121] = 12'h  0;
rom[30122] = 12'h  0;
rom[30123] = 12'h  0;
rom[30124] = 12'h  0;
rom[30125] = 12'h  0;
rom[30126] = 12'h100;
rom[30127] = 12'h100;
rom[30128] = 12'h100;
rom[30129] = 12'h100;
rom[30130] = 12'h200;
rom[30131] = 12'h200;
rom[30132] = 12'h300;
rom[30133] = 12'h300;
rom[30134] = 12'h400;
rom[30135] = 12'h410;
rom[30136] = 12'h510;
rom[30137] = 12'h510;
rom[30138] = 12'h610;
rom[30139] = 12'h610;
rom[30140] = 12'h610;
rom[30141] = 12'h620;
rom[30142] = 12'h720;
rom[30143] = 12'h720;
rom[30144] = 12'h720;
rom[30145] = 12'h720;
rom[30146] = 12'h720;
rom[30147] = 12'h720;
rom[30148] = 12'h720;
rom[30149] = 12'h710;
rom[30150] = 12'h710;
rom[30151] = 12'h710;
rom[30152] = 12'h710;
rom[30153] = 12'h710;
rom[30154] = 12'h610;
rom[30155] = 12'h610;
rom[30156] = 12'h600;
rom[30157] = 12'h500;
rom[30158] = 12'h500;
rom[30159] = 12'h500;
rom[30160] = 12'h400;
rom[30161] = 12'h300;
rom[30162] = 12'h300;
rom[30163] = 12'h300;
rom[30164] = 12'h300;
rom[30165] = 12'h200;
rom[30166] = 12'h200;
rom[30167] = 12'h200;
rom[30168] = 12'h100;
rom[30169] = 12'h100;
rom[30170] = 12'h100;
rom[30171] = 12'h100;
rom[30172] = 12'h  0;
rom[30173] = 12'h  0;
rom[30174] = 12'h  0;
rom[30175] = 12'h  0;
rom[30176] = 12'h  0;
rom[30177] = 12'h  0;
rom[30178] = 12'h  0;
rom[30179] = 12'h  0;
rom[30180] = 12'h100;
rom[30181] = 12'h100;
rom[30182] = 12'h111;
rom[30183] = 12'h111;
rom[30184] = 12'h111;
rom[30185] = 12'h100;
rom[30186] = 12'h  0;
rom[30187] = 12'h  0;
rom[30188] = 12'h  0;
rom[30189] = 12'h 10;
rom[30190] = 12'h  0;
rom[30191] = 12'h  0;
rom[30192] = 12'h  0;
rom[30193] = 12'h  0;
rom[30194] = 12'h  0;
rom[30195] = 12'h111;
rom[30196] = 12'h111;
rom[30197] = 12'h111;
rom[30198] = 12'h111;
rom[30199] = 12'h222;
rom[30200] = 12'h222;
rom[30201] = 12'h222;
rom[30202] = 12'h222;
rom[30203] = 12'h333;
rom[30204] = 12'h444;
rom[30205] = 12'h555;
rom[30206] = 12'h666;
rom[30207] = 12'h777;
rom[30208] = 12'h777;
rom[30209] = 12'h888;
rom[30210] = 12'h888;
rom[30211] = 12'h777;
rom[30212] = 12'h777;
rom[30213] = 12'h777;
rom[30214] = 12'h666;
rom[30215] = 12'h666;
rom[30216] = 12'h666;
rom[30217] = 12'h666;
rom[30218] = 12'h666;
rom[30219] = 12'h666;
rom[30220] = 12'h666;
rom[30221] = 12'h666;
rom[30222] = 12'h666;
rom[30223] = 12'h666;
rom[30224] = 12'h666;
rom[30225] = 12'h666;
rom[30226] = 12'h666;
rom[30227] = 12'h666;
rom[30228] = 12'h666;
rom[30229] = 12'h666;
rom[30230] = 12'h777;
rom[30231] = 12'h777;
rom[30232] = 12'h777;
rom[30233] = 12'h666;
rom[30234] = 12'h666;
rom[30235] = 12'h666;
rom[30236] = 12'h666;
rom[30237] = 12'h555;
rom[30238] = 12'h444;
rom[30239] = 12'h444;
rom[30240] = 12'h333;
rom[30241] = 12'h333;
rom[30242] = 12'h222;
rom[30243] = 12'h222;
rom[30244] = 12'h222;
rom[30245] = 12'h222;
rom[30246] = 12'h222;
rom[30247] = 12'h222;
rom[30248] = 12'h111;
rom[30249] = 12'h111;
rom[30250] = 12'h111;
rom[30251] = 12'h  0;
rom[30252] = 12'h  0;
rom[30253] = 12'h  0;
rom[30254] = 12'h  0;
rom[30255] = 12'h111;
rom[30256] = 12'h  0;
rom[30257] = 12'h  0;
rom[30258] = 12'h  0;
rom[30259] = 12'h  0;
rom[30260] = 12'h  0;
rom[30261] = 12'h  0;
rom[30262] = 12'h  0;
rom[30263] = 12'h  0;
rom[30264] = 12'h  0;
rom[30265] = 12'h  0;
rom[30266] = 12'h  0;
rom[30267] = 12'h  0;
rom[30268] = 12'h  0;
rom[30269] = 12'h  0;
rom[30270] = 12'h  0;
rom[30271] = 12'h  0;
rom[30272] = 12'h  0;
rom[30273] = 12'h  0;
rom[30274] = 12'h  0;
rom[30275] = 12'h  0;
rom[30276] = 12'h  0;
rom[30277] = 12'h  0;
rom[30278] = 12'h  0;
rom[30279] = 12'h  0;
rom[30280] = 12'h  0;
rom[30281] = 12'h  0;
rom[30282] = 12'h  0;
rom[30283] = 12'h  0;
rom[30284] = 12'h  0;
rom[30285] = 12'h  0;
rom[30286] = 12'h  0;
rom[30287] = 12'h111;
rom[30288] = 12'h111;
rom[30289] = 12'h111;
rom[30290] = 12'h222;
rom[30291] = 12'h222;
rom[30292] = 12'h222;
rom[30293] = 12'h222;
rom[30294] = 12'h333;
rom[30295] = 12'h333;
rom[30296] = 12'h333;
rom[30297] = 12'h333;
rom[30298] = 12'h333;
rom[30299] = 12'h333;
rom[30300] = 12'h444;
rom[30301] = 12'h555;
rom[30302] = 12'h555;
rom[30303] = 12'h666;
rom[30304] = 12'h666;
rom[30305] = 12'h766;
rom[30306] = 12'h777;
rom[30307] = 12'h888;
rom[30308] = 12'h988;
rom[30309] = 12'h999;
rom[30310] = 12'haaa;
rom[30311] = 12'hbaa;
rom[30312] = 12'hbbb;
rom[30313] = 12'hccc;
rom[30314] = 12'hddd;
rom[30315] = 12'heee;
rom[30316] = 12'hfff;
rom[30317] = 12'hfff;
rom[30318] = 12'heed;
rom[30319] = 12'hbbb;
rom[30320] = 12'h555;
rom[30321] = 12'h443;
rom[30322] = 12'h221;
rom[30323] = 12'h110;
rom[30324] = 12'h211;
rom[30325] = 12'h221;
rom[30326] = 12'h211;
rom[30327] = 12'h110;
rom[30328] = 12'h100;
rom[30329] = 12'h100;
rom[30330] = 12'h100;
rom[30331] = 12'h200;
rom[30332] = 12'h200;
rom[30333] = 12'h200;
rom[30334] = 12'h200;
rom[30335] = 12'h200;
rom[30336] = 12'h200;
rom[30337] = 12'h300;
rom[30338] = 12'h300;
rom[30339] = 12'h300;
rom[30340] = 12'h400;
rom[30341] = 12'h400;
rom[30342] = 12'h500;
rom[30343] = 12'h600;
rom[30344] = 12'h710;
rom[30345] = 12'h810;
rom[30346] = 12'h920;
rom[30347] = 12'ha30;
rom[30348] = 12'hc30;
rom[30349] = 12'hd40;
rom[30350] = 12'hd40;
rom[30351] = 12'hd40;
rom[30352] = 12'hd40;
rom[30353] = 12'hc50;
rom[30354] = 12'hc50;
rom[30355] = 12'hb50;
rom[30356] = 12'hb50;
rom[30357] = 12'hb61;
rom[30358] = 12'hb71;
rom[30359] = 12'hb72;
rom[30360] = 12'ha61;
rom[30361] = 12'h950;
rom[30362] = 12'h840;
rom[30363] = 12'h840;
rom[30364] = 12'h740;
rom[30365] = 12'h740;
rom[30366] = 12'h740;
rom[30367] = 12'h640;
rom[30368] = 12'h641;
rom[30369] = 12'h641;
rom[30370] = 12'h642;
rom[30371] = 12'h642;
rom[30372] = 12'h642;
rom[30373] = 12'h543;
rom[30374] = 12'h543;
rom[30375] = 12'h554;
rom[30376] = 12'h554;
rom[30377] = 12'h655;
rom[30378] = 12'h666;
rom[30379] = 12'h776;
rom[30380] = 12'h777;
rom[30381] = 12'h777;
rom[30382] = 12'h888;
rom[30383] = 12'h888;
rom[30384] = 12'h888;
rom[30385] = 12'h999;
rom[30386] = 12'h999;
rom[30387] = 12'h999;
rom[30388] = 12'h999;
rom[30389] = 12'h999;
rom[30390] = 12'h888;
rom[30391] = 12'h888;
rom[30392] = 12'h999;
rom[30393] = 12'h999;
rom[30394] = 12'h999;
rom[30395] = 12'haaa;
rom[30396] = 12'haaa;
rom[30397] = 12'haaa;
rom[30398] = 12'haaa;
rom[30399] = 12'haaa;
rom[30400] = 12'h777;
rom[30401] = 12'h666;
rom[30402] = 12'h666;
rom[30403] = 12'h666;
rom[30404] = 12'h666;
rom[30405] = 12'h666;
rom[30406] = 12'h666;
rom[30407] = 12'h666;
rom[30408] = 12'h666;
rom[30409] = 12'h666;
rom[30410] = 12'h666;
rom[30411] = 12'h666;
rom[30412] = 12'h666;
rom[30413] = 12'h666;
rom[30414] = 12'h666;
rom[30415] = 12'h666;
rom[30416] = 12'h666;
rom[30417] = 12'h666;
rom[30418] = 12'h666;
rom[30419] = 12'h666;
rom[30420] = 12'h666;
rom[30421] = 12'h666;
rom[30422] = 12'h666;
rom[30423] = 12'h666;
rom[30424] = 12'h666;
rom[30425] = 12'h666;
rom[30426] = 12'h666;
rom[30427] = 12'h777;
rom[30428] = 12'h777;
rom[30429] = 12'h777;
rom[30430] = 12'h777;
rom[30431] = 12'h777;
rom[30432] = 12'h888;
rom[30433] = 12'h888;
rom[30434] = 12'h888;
rom[30435] = 12'h888;
rom[30436] = 12'h888;
rom[30437] = 12'h888;
rom[30438] = 12'h999;
rom[30439] = 12'h999;
rom[30440] = 12'h999;
rom[30441] = 12'h888;
rom[30442] = 12'h888;
rom[30443] = 12'h888;
rom[30444] = 12'h777;
rom[30445] = 12'h777;
rom[30446] = 12'h777;
rom[30447] = 12'h666;
rom[30448] = 12'h666;
rom[30449] = 12'h666;
rom[30450] = 12'h666;
rom[30451] = 12'h666;
rom[30452] = 12'h666;
rom[30453] = 12'h666;
rom[30454] = 12'h666;
rom[30455] = 12'h666;
rom[30456] = 12'h777;
rom[30457] = 12'h777;
rom[30458] = 12'h777;
rom[30459] = 12'h777;
rom[30460] = 12'h888;
rom[30461] = 12'h888;
rom[30462] = 12'h888;
rom[30463] = 12'h888;
rom[30464] = 12'h888;
rom[30465] = 12'h888;
rom[30466] = 12'h777;
rom[30467] = 12'h777;
rom[30468] = 12'h666;
rom[30469] = 12'h666;
rom[30470] = 12'h666;
rom[30471] = 12'h666;
rom[30472] = 12'h555;
rom[30473] = 12'h555;
rom[30474] = 12'h444;
rom[30475] = 12'h444;
rom[30476] = 12'h444;
rom[30477] = 12'h444;
rom[30478] = 12'h444;
rom[30479] = 12'h333;
rom[30480] = 12'h333;
rom[30481] = 12'h333;
rom[30482] = 12'h333;
rom[30483] = 12'h333;
rom[30484] = 12'h333;
rom[30485] = 12'h333;
rom[30486] = 12'h222;
rom[30487] = 12'h222;
rom[30488] = 12'h222;
rom[30489] = 12'h222;
rom[30490] = 12'h222;
rom[30491] = 12'h222;
rom[30492] = 12'h111;
rom[30493] = 12'h111;
rom[30494] = 12'h111;
rom[30495] = 12'h  0;
rom[30496] = 12'h  0;
rom[30497] = 12'h  0;
rom[30498] = 12'h  0;
rom[30499] = 12'h  0;
rom[30500] = 12'h  0;
rom[30501] = 12'h  0;
rom[30502] = 12'h  0;
rom[30503] = 12'h  0;
rom[30504] = 12'h  0;
rom[30505] = 12'h  0;
rom[30506] = 12'h  0;
rom[30507] = 12'h  0;
rom[30508] = 12'h  0;
rom[30509] = 12'h  0;
rom[30510] = 12'h  0;
rom[30511] = 12'h  0;
rom[30512] = 12'h  0;
rom[30513] = 12'h  0;
rom[30514] = 12'h  0;
rom[30515] = 12'h  0;
rom[30516] = 12'h  0;
rom[30517] = 12'h  0;
rom[30518] = 12'h  0;
rom[30519] = 12'h  0;
rom[30520] = 12'h  0;
rom[30521] = 12'h  0;
rom[30522] = 12'h  0;
rom[30523] = 12'h  0;
rom[30524] = 12'h  0;
rom[30525] = 12'h  0;
rom[30526] = 12'h  0;
rom[30527] = 12'h100;
rom[30528] = 12'h100;
rom[30529] = 12'h200;
rom[30530] = 12'h200;
rom[30531] = 12'h200;
rom[30532] = 12'h200;
rom[30533] = 12'h300;
rom[30534] = 12'h300;
rom[30535] = 12'h400;
rom[30536] = 12'h400;
rom[30537] = 12'h400;
rom[30538] = 12'h510;
rom[30539] = 12'h510;
rom[30540] = 12'h510;
rom[30541] = 12'h510;
rom[30542] = 12'h510;
rom[30543] = 12'h510;
rom[30544] = 12'h510;
rom[30545] = 12'h610;
rom[30546] = 12'h610;
rom[30547] = 12'h610;
rom[30548] = 12'h610;
rom[30549] = 12'h610;
rom[30550] = 12'h610;
rom[30551] = 12'h610;
rom[30552] = 12'h510;
rom[30553] = 12'h510;
rom[30554] = 12'h510;
rom[30555] = 12'h510;
rom[30556] = 12'h400;
rom[30557] = 12'h400;
rom[30558] = 12'h400;
rom[30559] = 12'h300;
rom[30560] = 12'h300;
rom[30561] = 12'h300;
rom[30562] = 12'h200;
rom[30563] = 12'h200;
rom[30564] = 12'h200;
rom[30565] = 12'h200;
rom[30566] = 12'h200;
rom[30567] = 12'h100;
rom[30568] = 12'h100;
rom[30569] = 12'h100;
rom[30570] = 12'h100;
rom[30571] = 12'h  0;
rom[30572] = 12'h  0;
rom[30573] = 12'h  0;
rom[30574] = 12'h  0;
rom[30575] = 12'h  0;
rom[30576] = 12'h  0;
rom[30577] = 12'h  0;
rom[30578] = 12'h  0;
rom[30579] = 12'h  0;
rom[30580] = 12'h100;
rom[30581] = 12'h100;
rom[30582] = 12'h111;
rom[30583] = 12'h111;
rom[30584] = 12'h100;
rom[30585] = 12'h  0;
rom[30586] = 12'h  0;
rom[30587] = 12'h  0;
rom[30588] = 12'h  0;
rom[30589] = 12'h  0;
rom[30590] = 12'h  0;
rom[30591] = 12'h  0;
rom[30592] = 12'h  0;
rom[30593] = 12'h  0;
rom[30594] = 12'h  0;
rom[30595] = 12'h  0;
rom[30596] = 12'h111;
rom[30597] = 12'h111;
rom[30598] = 12'h111;
rom[30599] = 12'h222;
rom[30600] = 12'h222;
rom[30601] = 12'h222;
rom[30602] = 12'h333;
rom[30603] = 12'h333;
rom[30604] = 12'h444;
rom[30605] = 12'h555;
rom[30606] = 12'h666;
rom[30607] = 12'h777;
rom[30608] = 12'h888;
rom[30609] = 12'h888;
rom[30610] = 12'h777;
rom[30611] = 12'h777;
rom[30612] = 12'h666;
rom[30613] = 12'h666;
rom[30614] = 12'h666;
rom[30615] = 12'h666;
rom[30616] = 12'h666;
rom[30617] = 12'h666;
rom[30618] = 12'h666;
rom[30619] = 12'h666;
rom[30620] = 12'h666;
rom[30621] = 12'h666;
rom[30622] = 12'h666;
rom[30623] = 12'h666;
rom[30624] = 12'h666;
rom[30625] = 12'h666;
rom[30626] = 12'h666;
rom[30627] = 12'h666;
rom[30628] = 12'h666;
rom[30629] = 12'h666;
rom[30630] = 12'h777;
rom[30631] = 12'h777;
rom[30632] = 12'h666;
rom[30633] = 12'h666;
rom[30634] = 12'h666;
rom[30635] = 12'h666;
rom[30636] = 12'h666;
rom[30637] = 12'h555;
rom[30638] = 12'h444;
rom[30639] = 12'h333;
rom[30640] = 12'h333;
rom[30641] = 12'h333;
rom[30642] = 12'h222;
rom[30643] = 12'h222;
rom[30644] = 12'h222;
rom[30645] = 12'h222;
rom[30646] = 12'h222;
rom[30647] = 12'h111;
rom[30648] = 12'h111;
rom[30649] = 12'h111;
rom[30650] = 12'h111;
rom[30651] = 12'h  0;
rom[30652] = 12'h  0;
rom[30653] = 12'h  0;
rom[30654] = 12'h111;
rom[30655] = 12'h111;
rom[30656] = 12'h  0;
rom[30657] = 12'h  0;
rom[30658] = 12'h  0;
rom[30659] = 12'h  0;
rom[30660] = 12'h  0;
rom[30661] = 12'h  0;
rom[30662] = 12'h  0;
rom[30663] = 12'h  0;
rom[30664] = 12'h  0;
rom[30665] = 12'h  0;
rom[30666] = 12'h  0;
rom[30667] = 12'h  0;
rom[30668] = 12'h  0;
rom[30669] = 12'h  0;
rom[30670] = 12'h  0;
rom[30671] = 12'h  0;
rom[30672] = 12'h  0;
rom[30673] = 12'h  0;
rom[30674] = 12'h  0;
rom[30675] = 12'h  0;
rom[30676] = 12'h  0;
rom[30677] = 12'h  0;
rom[30678] = 12'h  0;
rom[30679] = 12'h  0;
rom[30680] = 12'h  0;
rom[30681] = 12'h  0;
rom[30682] = 12'h  0;
rom[30683] = 12'h  0;
rom[30684] = 12'h  0;
rom[30685] = 12'h  0;
rom[30686] = 12'h111;
rom[30687] = 12'h111;
rom[30688] = 12'h111;
rom[30689] = 12'h222;
rom[30690] = 12'h222;
rom[30691] = 12'h222;
rom[30692] = 12'h222;
rom[30693] = 12'h222;
rom[30694] = 12'h333;
rom[30695] = 12'h333;
rom[30696] = 12'h333;
rom[30697] = 12'h333;
rom[30698] = 12'h333;
rom[30699] = 12'h444;
rom[30700] = 12'h444;
rom[30701] = 12'h555;
rom[30702] = 12'h666;
rom[30703] = 12'h666;
rom[30704] = 12'h766;
rom[30705] = 12'h776;
rom[30706] = 12'h877;
rom[30707] = 12'h888;
rom[30708] = 12'h999;
rom[30709] = 12'ha99;
rom[30710] = 12'haaa;
rom[30711] = 12'hbbb;
rom[30712] = 12'hdcc;
rom[30713] = 12'heed;
rom[30714] = 12'hffe;
rom[30715] = 12'hfff;
rom[30716] = 12'hfff;
rom[30717] = 12'hedd;
rom[30718] = 12'h999;
rom[30719] = 12'h555;
rom[30720] = 12'h332;
rom[30721] = 12'h221;
rom[30722] = 12'h100;
rom[30723] = 12'h  0;
rom[30724] = 12'h  0;
rom[30725] = 12'h100;
rom[30726] = 12'h  0;
rom[30727] = 12'h  0;
rom[30728] = 12'h  0;
rom[30729] = 12'h100;
rom[30730] = 12'h100;
rom[30731] = 12'h100;
rom[30732] = 12'h100;
rom[30733] = 12'h200;
rom[30734] = 12'h200;
rom[30735] = 12'h200;
rom[30736] = 12'h200;
rom[30737] = 12'h200;
rom[30738] = 12'h200;
rom[30739] = 12'h300;
rom[30740] = 12'h300;
rom[30741] = 12'h400;
rom[30742] = 12'h500;
rom[30743] = 12'h500;
rom[30744] = 12'h710;
rom[30745] = 12'h810;
rom[30746] = 12'h920;
rom[30747] = 12'ha30;
rom[30748] = 12'hc30;
rom[30749] = 12'hd40;
rom[30750] = 12'hd40;
rom[30751] = 12'hd40;
rom[30752] = 12'hd50;
rom[30753] = 12'hd50;
rom[30754] = 12'hc50;
rom[30755] = 12'hb50;
rom[30756] = 12'hb60;
rom[30757] = 12'hc71;
rom[30758] = 12'hb72;
rom[30759] = 12'hb72;
rom[30760] = 12'h950;
rom[30761] = 12'h850;
rom[30762] = 12'h840;
rom[30763] = 12'h840;
rom[30764] = 12'h740;
rom[30765] = 12'h740;
rom[30766] = 12'h640;
rom[30767] = 12'h640;
rom[30768] = 12'h641;
rom[30769] = 12'h642;
rom[30770] = 12'h642;
rom[30771] = 12'h642;
rom[30772] = 12'h542;
rom[30773] = 12'h542;
rom[30774] = 12'h543;
rom[30775] = 12'h544;
rom[30776] = 12'h554;
rom[30777] = 12'h555;
rom[30778] = 12'h666;
rom[30779] = 12'h766;
rom[30780] = 12'h777;
rom[30781] = 12'h777;
rom[30782] = 12'h777;
rom[30783] = 12'h888;
rom[30784] = 12'h888;
rom[30785] = 12'h888;
rom[30786] = 12'h999;
rom[30787] = 12'h999;
rom[30788] = 12'h999;
rom[30789] = 12'h999;
rom[30790] = 12'h999;
rom[30791] = 12'h999;
rom[30792] = 12'h999;
rom[30793] = 12'h999;
rom[30794] = 12'h999;
rom[30795] = 12'haaa;
rom[30796] = 12'haaa;
rom[30797] = 12'haaa;
rom[30798] = 12'haaa;
rom[30799] = 12'haaa;
rom[30800] = 12'h777;
rom[30801] = 12'h777;
rom[30802] = 12'h666;
rom[30803] = 12'h666;
rom[30804] = 12'h666;
rom[30805] = 12'h666;
rom[30806] = 12'h666;
rom[30807] = 12'h666;
rom[30808] = 12'h666;
rom[30809] = 12'h666;
rom[30810] = 12'h666;
rom[30811] = 12'h666;
rom[30812] = 12'h666;
rom[30813] = 12'h666;
rom[30814] = 12'h666;
rom[30815] = 12'h666;
rom[30816] = 12'h666;
rom[30817] = 12'h666;
rom[30818] = 12'h666;
rom[30819] = 12'h666;
rom[30820] = 12'h666;
rom[30821] = 12'h666;
rom[30822] = 12'h666;
rom[30823] = 12'h666;
rom[30824] = 12'h777;
rom[30825] = 12'h777;
rom[30826] = 12'h777;
rom[30827] = 12'h777;
rom[30828] = 12'h777;
rom[30829] = 12'h777;
rom[30830] = 12'h888;
rom[30831] = 12'h888;
rom[30832] = 12'h888;
rom[30833] = 12'h888;
rom[30834] = 12'h888;
rom[30835] = 12'h888;
rom[30836] = 12'h888;
rom[30837] = 12'h888;
rom[30838] = 12'h999;
rom[30839] = 12'h999;
rom[30840] = 12'h999;
rom[30841] = 12'h888;
rom[30842] = 12'h888;
rom[30843] = 12'h888;
rom[30844] = 12'h777;
rom[30845] = 12'h777;
rom[30846] = 12'h777;
rom[30847] = 12'h666;
rom[30848] = 12'h666;
rom[30849] = 12'h666;
rom[30850] = 12'h666;
rom[30851] = 12'h666;
rom[30852] = 12'h666;
rom[30853] = 12'h666;
rom[30854] = 12'h666;
rom[30855] = 12'h666;
rom[30856] = 12'h666;
rom[30857] = 12'h666;
rom[30858] = 12'h777;
rom[30859] = 12'h777;
rom[30860] = 12'h777;
rom[30861] = 12'h888;
rom[30862] = 12'h888;
rom[30863] = 12'h888;
rom[30864] = 12'h999;
rom[30865] = 12'h888;
rom[30866] = 12'h888;
rom[30867] = 12'h777;
rom[30868] = 12'h777;
rom[30869] = 12'h666;
rom[30870] = 12'h666;
rom[30871] = 12'h666;
rom[30872] = 12'h555;
rom[30873] = 12'h555;
rom[30874] = 12'h555;
rom[30875] = 12'h444;
rom[30876] = 12'h444;
rom[30877] = 12'h444;
rom[30878] = 12'h444;
rom[30879] = 12'h444;
rom[30880] = 12'h333;
rom[30881] = 12'h333;
rom[30882] = 12'h333;
rom[30883] = 12'h333;
rom[30884] = 12'h333;
rom[30885] = 12'h333;
rom[30886] = 12'h222;
rom[30887] = 12'h222;
rom[30888] = 12'h222;
rom[30889] = 12'h222;
rom[30890] = 12'h222;
rom[30891] = 12'h222;
rom[30892] = 12'h111;
rom[30893] = 12'h111;
rom[30894] = 12'h111;
rom[30895] = 12'h  0;
rom[30896] = 12'h  0;
rom[30897] = 12'h  0;
rom[30898] = 12'h  0;
rom[30899] = 12'h  0;
rom[30900] = 12'h  0;
rom[30901] = 12'h  0;
rom[30902] = 12'h  0;
rom[30903] = 12'h  0;
rom[30904] = 12'h  0;
rom[30905] = 12'h  0;
rom[30906] = 12'h  0;
rom[30907] = 12'h  0;
rom[30908] = 12'h  0;
rom[30909] = 12'h  0;
rom[30910] = 12'h  0;
rom[30911] = 12'h  0;
rom[30912] = 12'h  0;
rom[30913] = 12'h  0;
rom[30914] = 12'h  0;
rom[30915] = 12'h  0;
rom[30916] = 12'h  0;
rom[30917] = 12'h  0;
rom[30918] = 12'h  0;
rom[30919] = 12'h  0;
rom[30920] = 12'h  0;
rom[30921] = 12'h  0;
rom[30922] = 12'h  0;
rom[30923] = 12'h  0;
rom[30924] = 12'h  0;
rom[30925] = 12'h  0;
rom[30926] = 12'h  0;
rom[30927] = 12'h100;
rom[30928] = 12'h100;
rom[30929] = 12'h200;
rom[30930] = 12'h200;
rom[30931] = 12'h200;
rom[30932] = 12'h200;
rom[30933] = 12'h300;
rom[30934] = 12'h300;
rom[30935] = 12'h300;
rom[30936] = 12'h400;
rom[30937] = 12'h400;
rom[30938] = 12'h400;
rom[30939] = 12'h400;
rom[30940] = 12'h410;
rom[30941] = 12'h410;
rom[30942] = 12'h410;
rom[30943] = 12'h410;
rom[30944] = 12'h410;
rom[30945] = 12'h410;
rom[30946] = 12'h510;
rom[30947] = 12'h510;
rom[30948] = 12'h510;
rom[30949] = 12'h510;
rom[30950] = 12'h510;
rom[30951] = 12'h510;
rom[30952] = 12'h410;
rom[30953] = 12'h400;
rom[30954] = 12'h400;
rom[30955] = 12'h300;
rom[30956] = 12'h300;
rom[30957] = 12'h300;
rom[30958] = 12'h300;
rom[30959] = 12'h200;
rom[30960] = 12'h200;
rom[30961] = 12'h200;
rom[30962] = 12'h200;
rom[30963] = 12'h200;
rom[30964] = 12'h100;
rom[30965] = 12'h100;
rom[30966] = 12'h100;
rom[30967] = 12'h100;
rom[30968] = 12'h100;
rom[30969] = 12'h  0;
rom[30970] = 12'h  0;
rom[30971] = 12'h  0;
rom[30972] = 12'h  0;
rom[30973] = 12'h  0;
rom[30974] = 12'h  0;
rom[30975] = 12'h  0;
rom[30976] = 12'h  0;
rom[30977] = 12'h  0;
rom[30978] = 12'h  0;
rom[30979] = 12'h  0;
rom[30980] = 12'h  0;
rom[30981] = 12'h  0;
rom[30982] = 12'h100;
rom[30983] = 12'h  0;
rom[30984] = 12'h  0;
rom[30985] = 12'h  0;
rom[30986] = 12'h  0;
rom[30987] = 12'h  0;
rom[30988] = 12'h  0;
rom[30989] = 12'h  0;
rom[30990] = 12'h  0;
rom[30991] = 12'h  0;
rom[30992] = 12'h  0;
rom[30993] = 12'h  0;
rom[30994] = 12'h  0;
rom[30995] = 12'h  0;
rom[30996] = 12'h111;
rom[30997] = 12'h111;
rom[30998] = 12'h111;
rom[30999] = 12'h111;
rom[31000] = 12'h222;
rom[31001] = 12'h222;
rom[31002] = 12'h333;
rom[31003] = 12'h444;
rom[31004] = 12'h444;
rom[31005] = 12'h555;
rom[31006] = 12'h666;
rom[31007] = 12'h666;
rom[31008] = 12'h777;
rom[31009] = 12'h777;
rom[31010] = 12'h777;
rom[31011] = 12'h777;
rom[31012] = 12'h666;
rom[31013] = 12'h666;
rom[31014] = 12'h666;
rom[31015] = 12'h666;
rom[31016] = 12'h666;
rom[31017] = 12'h666;
rom[31018] = 12'h666;
rom[31019] = 12'h666;
rom[31020] = 12'h666;
rom[31021] = 12'h666;
rom[31022] = 12'h666;
rom[31023] = 12'h666;
rom[31024] = 12'h666;
rom[31025] = 12'h666;
rom[31026] = 12'h666;
rom[31027] = 12'h666;
rom[31028] = 12'h666;
rom[31029] = 12'h666;
rom[31030] = 12'h666;
rom[31031] = 12'h777;
rom[31032] = 12'h666;
rom[31033] = 12'h666;
rom[31034] = 12'h666;
rom[31035] = 12'h666;
rom[31036] = 12'h555;
rom[31037] = 12'h555;
rom[31038] = 12'h444;
rom[31039] = 12'h333;
rom[31040] = 12'h333;
rom[31041] = 12'h333;
rom[31042] = 12'h222;
rom[31043] = 12'h222;
rom[31044] = 12'h222;
rom[31045] = 12'h222;
rom[31046] = 12'h111;
rom[31047] = 12'h111;
rom[31048] = 12'h111;
rom[31049] = 12'h111;
rom[31050] = 12'h111;
rom[31051] = 12'h  0;
rom[31052] = 12'h  0;
rom[31053] = 12'h  0;
rom[31054] = 12'h111;
rom[31055] = 12'h111;
rom[31056] = 12'h  0;
rom[31057] = 12'h  0;
rom[31058] = 12'h  0;
rom[31059] = 12'h  0;
rom[31060] = 12'h  0;
rom[31061] = 12'h  0;
rom[31062] = 12'h  0;
rom[31063] = 12'h  0;
rom[31064] = 12'h  0;
rom[31065] = 12'h  0;
rom[31066] = 12'h  0;
rom[31067] = 12'h  0;
rom[31068] = 12'h  0;
rom[31069] = 12'h  0;
rom[31070] = 12'h  0;
rom[31071] = 12'h  0;
rom[31072] = 12'h  0;
rom[31073] = 12'h  0;
rom[31074] = 12'h  0;
rom[31075] = 12'h  0;
rom[31076] = 12'h  0;
rom[31077] = 12'h  0;
rom[31078] = 12'h  0;
rom[31079] = 12'h  0;
rom[31080] = 12'h  0;
rom[31081] = 12'h  0;
rom[31082] = 12'h  0;
rom[31083] = 12'h  0;
rom[31084] = 12'h  0;
rom[31085] = 12'h  0;
rom[31086] = 12'h111;
rom[31087] = 12'h111;
rom[31088] = 12'h111;
rom[31089] = 12'h222;
rom[31090] = 12'h222;
rom[31091] = 12'h222;
rom[31092] = 12'h222;
rom[31093] = 12'h222;
rom[31094] = 12'h333;
rom[31095] = 12'h333;
rom[31096] = 12'h333;
rom[31097] = 12'h333;
rom[31098] = 12'h444;
rom[31099] = 12'h444;
rom[31100] = 12'h555;
rom[31101] = 12'h666;
rom[31102] = 12'h666;
rom[31103] = 12'h776;
rom[31104] = 12'h777;
rom[31105] = 12'h777;
rom[31106] = 12'h888;
rom[31107] = 12'h999;
rom[31108] = 12'ha99;
rom[31109] = 12'haaa;
rom[31110] = 12'hbbb;
rom[31111] = 12'hdcc;
rom[31112] = 12'heed;
rom[31113] = 12'hfff;
rom[31114] = 12'hfff;
rom[31115] = 12'hfff;
rom[31116] = 12'hdcc;
rom[31117] = 12'h988;
rom[31118] = 12'h444;
rom[31119] = 12'h111;
rom[31120] = 12'h111;
rom[31121] = 12'h 10;
rom[31122] = 12'h  0;
rom[31123] = 12'h  0;
rom[31124] = 12'h  0;
rom[31125] = 12'h  0;
rom[31126] = 12'h  0;
rom[31127] = 12'h  0;
rom[31128] = 12'h  0;
rom[31129] = 12'h  0;
rom[31130] = 12'h  0;
rom[31131] = 12'h100;
rom[31132] = 12'h100;
rom[31133] = 12'h100;
rom[31134] = 12'h100;
rom[31135] = 12'h100;
rom[31136] = 12'h200;
rom[31137] = 12'h200;
rom[31138] = 12'h200;
rom[31139] = 12'h200;
rom[31140] = 12'h300;
rom[31141] = 12'h300;
rom[31142] = 12'h400;
rom[31143] = 12'h500;
rom[31144] = 12'h610;
rom[31145] = 12'h710;
rom[31146] = 12'h920;
rom[31147] = 12'ha30;
rom[31148] = 12'hc40;
rom[31149] = 12'hd40;
rom[31150] = 12'hd50;
rom[31151] = 12'he50;
rom[31152] = 12'hd50;
rom[31153] = 12'hd50;
rom[31154] = 12'hc50;
rom[31155] = 12'hc60;
rom[31156] = 12'hc70;
rom[31157] = 12'hc82;
rom[31158] = 12'hc82;
rom[31159] = 12'hb71;
rom[31160] = 12'h950;
rom[31161] = 12'h850;
rom[31162] = 12'h840;
rom[31163] = 12'h840;
rom[31164] = 12'h740;
rom[31165] = 12'h740;
rom[31166] = 12'h640;
rom[31167] = 12'h641;
rom[31168] = 12'h641;
rom[31169] = 12'h641;
rom[31170] = 12'h642;
rom[31171] = 12'h542;
rom[31172] = 12'h542;
rom[31173] = 12'h542;
rom[31174] = 12'h543;
rom[31175] = 12'h543;
rom[31176] = 12'h544;
rom[31177] = 12'h555;
rom[31178] = 12'h665;
rom[31179] = 12'h666;
rom[31180] = 12'h666;
rom[31181] = 12'h777;
rom[31182] = 12'h777;
rom[31183] = 12'h777;
rom[31184] = 12'h888;
rom[31185] = 12'h888;
rom[31186] = 12'h999;
rom[31187] = 12'h999;
rom[31188] = 12'h999;
rom[31189] = 12'h999;
rom[31190] = 12'h999;
rom[31191] = 12'h999;
rom[31192] = 12'h999;
rom[31193] = 12'h999;
rom[31194] = 12'h999;
rom[31195] = 12'haaa;
rom[31196] = 12'haaa;
rom[31197] = 12'haaa;
rom[31198] = 12'haaa;
rom[31199] = 12'hbbb;
rom[31200] = 12'h777;
rom[31201] = 12'h777;
rom[31202] = 12'h777;
rom[31203] = 12'h666;
rom[31204] = 12'h666;
rom[31205] = 12'h666;
rom[31206] = 12'h777;
rom[31207] = 12'h777;
rom[31208] = 12'h666;
rom[31209] = 12'h666;
rom[31210] = 12'h666;
rom[31211] = 12'h666;
rom[31212] = 12'h666;
rom[31213] = 12'h666;
rom[31214] = 12'h666;
rom[31215] = 12'h666;
rom[31216] = 12'h777;
rom[31217] = 12'h777;
rom[31218] = 12'h777;
rom[31219] = 12'h777;
rom[31220] = 12'h777;
rom[31221] = 12'h777;
rom[31222] = 12'h777;
rom[31223] = 12'h777;
rom[31224] = 12'h777;
rom[31225] = 12'h777;
rom[31226] = 12'h888;
rom[31227] = 12'h888;
rom[31228] = 12'h888;
rom[31229] = 12'h888;
rom[31230] = 12'h888;
rom[31231] = 12'h888;
rom[31232] = 12'h888;
rom[31233] = 12'h888;
rom[31234] = 12'h888;
rom[31235] = 12'h888;
rom[31236] = 12'h888;
rom[31237] = 12'h888;
rom[31238] = 12'h999;
rom[31239] = 12'h999;
rom[31240] = 12'h999;
rom[31241] = 12'h888;
rom[31242] = 12'h888;
rom[31243] = 12'h888;
rom[31244] = 12'h888;
rom[31245] = 12'h777;
rom[31246] = 12'h777;
rom[31247] = 12'h777;
rom[31248] = 12'h666;
rom[31249] = 12'h666;
rom[31250] = 12'h666;
rom[31251] = 12'h666;
rom[31252] = 12'h666;
rom[31253] = 12'h666;
rom[31254] = 12'h666;
rom[31255] = 12'h666;
rom[31256] = 12'h666;
rom[31257] = 12'h666;
rom[31258] = 12'h666;
rom[31259] = 12'h777;
rom[31260] = 12'h777;
rom[31261] = 12'h888;
rom[31262] = 12'h888;
rom[31263] = 12'h999;
rom[31264] = 12'h999;
rom[31265] = 12'h999;
rom[31266] = 12'h888;
rom[31267] = 12'h888;
rom[31268] = 12'h777;
rom[31269] = 12'h777;
rom[31270] = 12'h666;
rom[31271] = 12'h666;
rom[31272] = 12'h666;
rom[31273] = 12'h555;
rom[31274] = 12'h555;
rom[31275] = 12'h555;
rom[31276] = 12'h444;
rom[31277] = 12'h444;
rom[31278] = 12'h444;
rom[31279] = 12'h444;
rom[31280] = 12'h333;
rom[31281] = 12'h333;
rom[31282] = 12'h333;
rom[31283] = 12'h333;
rom[31284] = 12'h333;
rom[31285] = 12'h333;
rom[31286] = 12'h222;
rom[31287] = 12'h222;
rom[31288] = 12'h222;
rom[31289] = 12'h222;
rom[31290] = 12'h222;
rom[31291] = 12'h222;
rom[31292] = 12'h222;
rom[31293] = 12'h111;
rom[31294] = 12'h111;
rom[31295] = 12'h  0;
rom[31296] = 12'h  0;
rom[31297] = 12'h  0;
rom[31298] = 12'h  0;
rom[31299] = 12'h  0;
rom[31300] = 12'h  0;
rom[31301] = 12'h  0;
rom[31302] = 12'h  0;
rom[31303] = 12'h  0;
rom[31304] = 12'h  0;
rom[31305] = 12'h  0;
rom[31306] = 12'h  0;
rom[31307] = 12'h  0;
rom[31308] = 12'h  0;
rom[31309] = 12'h  0;
rom[31310] = 12'h  0;
rom[31311] = 12'h  0;
rom[31312] = 12'h  0;
rom[31313] = 12'h  0;
rom[31314] = 12'h  0;
rom[31315] = 12'h  0;
rom[31316] = 12'h  0;
rom[31317] = 12'h  0;
rom[31318] = 12'h  0;
rom[31319] = 12'h  0;
rom[31320] = 12'h  0;
rom[31321] = 12'h  0;
rom[31322] = 12'h  0;
rom[31323] = 12'h  0;
rom[31324] = 12'h  0;
rom[31325] = 12'h  0;
rom[31326] = 12'h  0;
rom[31327] = 12'h  0;
rom[31328] = 12'h100;
rom[31329] = 12'h200;
rom[31330] = 12'h200;
rom[31331] = 12'h200;
rom[31332] = 12'h200;
rom[31333] = 12'h200;
rom[31334] = 12'h300;
rom[31335] = 12'h300;
rom[31336] = 12'h300;
rom[31337] = 12'h300;
rom[31338] = 12'h300;
rom[31339] = 12'h300;
rom[31340] = 12'h300;
rom[31341] = 12'h300;
rom[31342] = 12'h300;
rom[31343] = 12'h300;
rom[31344] = 12'h310;
rom[31345] = 12'h310;
rom[31346] = 12'h300;
rom[31347] = 12'h300;
rom[31348] = 12'h300;
rom[31349] = 12'h300;
rom[31350] = 12'h300;
rom[31351] = 12'h300;
rom[31352] = 12'h300;
rom[31353] = 12'h300;
rom[31354] = 12'h300;
rom[31355] = 12'h200;
rom[31356] = 12'h200;
rom[31357] = 12'h200;
rom[31358] = 12'h200;
rom[31359] = 12'h200;
rom[31360] = 12'h100;
rom[31361] = 12'h100;
rom[31362] = 12'h100;
rom[31363] = 12'h100;
rom[31364] = 12'h100;
rom[31365] = 12'h100;
rom[31366] = 12'h100;
rom[31367] = 12'h100;
rom[31368] = 12'h  0;
rom[31369] = 12'h  0;
rom[31370] = 12'h  0;
rom[31371] = 12'h  0;
rom[31372] = 12'h  0;
rom[31373] = 12'h  0;
rom[31374] = 12'h  0;
rom[31375] = 12'h  0;
rom[31376] = 12'h  0;
rom[31377] = 12'h  0;
rom[31378] = 12'h  0;
rom[31379] = 12'h  0;
rom[31380] = 12'h  0;
rom[31381] = 12'h  0;
rom[31382] = 12'h  0;
rom[31383] = 12'h  0;
rom[31384] = 12'h  0;
rom[31385] = 12'h  0;
rom[31386] = 12'h  0;
rom[31387] = 12'h  0;
rom[31388] = 12'h  0;
rom[31389] = 12'h  0;
rom[31390] = 12'h  0;
rom[31391] = 12'h  0;
rom[31392] = 12'h  0;
rom[31393] = 12'h  0;
rom[31394] = 12'h  0;
rom[31395] = 12'h  0;
rom[31396] = 12'h  0;
rom[31397] = 12'h111;
rom[31398] = 12'h111;
rom[31399] = 12'h111;
rom[31400] = 12'h111;
rom[31401] = 12'h222;
rom[31402] = 12'h333;
rom[31403] = 12'h333;
rom[31404] = 12'h444;
rom[31405] = 12'h555;
rom[31406] = 12'h666;
rom[31407] = 12'h666;
rom[31408] = 12'h777;
rom[31409] = 12'h777;
rom[31410] = 12'h777;
rom[31411] = 12'h666;
rom[31412] = 12'h666;
rom[31413] = 12'h666;
rom[31414] = 12'h666;
rom[31415] = 12'h666;
rom[31416] = 12'h666;
rom[31417] = 12'h666;
rom[31418] = 12'h666;
rom[31419] = 12'h666;
rom[31420] = 12'h666;
rom[31421] = 12'h666;
rom[31422] = 12'h666;
rom[31423] = 12'h666;
rom[31424] = 12'h666;
rom[31425] = 12'h666;
rom[31426] = 12'h666;
rom[31427] = 12'h666;
rom[31428] = 12'h666;
rom[31429] = 12'h666;
rom[31430] = 12'h666;
rom[31431] = 12'h666;
rom[31432] = 12'h666;
rom[31433] = 12'h666;
rom[31434] = 12'h666;
rom[31435] = 12'h666;
rom[31436] = 12'h555;
rom[31437] = 12'h555;
rom[31438] = 12'h444;
rom[31439] = 12'h333;
rom[31440] = 12'h333;
rom[31441] = 12'h333;
rom[31442] = 12'h222;
rom[31443] = 12'h222;
rom[31444] = 12'h222;
rom[31445] = 12'h222;
rom[31446] = 12'h111;
rom[31447] = 12'h111;
rom[31448] = 12'h111;
rom[31449] = 12'h111;
rom[31450] = 12'h111;
rom[31451] = 12'h  0;
rom[31452] = 12'h  0;
rom[31453] = 12'h  0;
rom[31454] = 12'h111;
rom[31455] = 12'h111;
rom[31456] = 12'h  0;
rom[31457] = 12'h  0;
rom[31458] = 12'h  0;
rom[31459] = 12'h  0;
rom[31460] = 12'h  0;
rom[31461] = 12'h  0;
rom[31462] = 12'h  0;
rom[31463] = 12'h  0;
rom[31464] = 12'h  0;
rom[31465] = 12'h  0;
rom[31466] = 12'h  0;
rom[31467] = 12'h  0;
rom[31468] = 12'h  0;
rom[31469] = 12'h  0;
rom[31470] = 12'h  0;
rom[31471] = 12'h  0;
rom[31472] = 12'h  0;
rom[31473] = 12'h  0;
rom[31474] = 12'h  0;
rom[31475] = 12'h  0;
rom[31476] = 12'h  0;
rom[31477] = 12'h  0;
rom[31478] = 12'h  0;
rom[31479] = 12'h  0;
rom[31480] = 12'h  0;
rom[31481] = 12'h  0;
rom[31482] = 12'h  0;
rom[31483] = 12'h  0;
rom[31484] = 12'h  0;
rom[31485] = 12'h  0;
rom[31486] = 12'h111;
rom[31487] = 12'h111;
rom[31488] = 12'h222;
rom[31489] = 12'h222;
rom[31490] = 12'h222;
rom[31491] = 12'h222;
rom[31492] = 12'h222;
rom[31493] = 12'h333;
rom[31494] = 12'h333;
rom[31495] = 12'h333;
rom[31496] = 12'h333;
rom[31497] = 12'h444;
rom[31498] = 12'h444;
rom[31499] = 12'h555;
rom[31500] = 12'h555;
rom[31501] = 12'h666;
rom[31502] = 12'h777;
rom[31503] = 12'h777;
rom[31504] = 12'h877;
rom[31505] = 12'h888;
rom[31506] = 12'h998;
rom[31507] = 12'haa9;
rom[31508] = 12'haaa;
rom[31509] = 12'hbbb;
rom[31510] = 12'hddc;
rom[31511] = 12'heee;
rom[31512] = 12'hffe;
rom[31513] = 12'hfff;
rom[31514] = 12'heee;
rom[31515] = 12'hbbb;
rom[31516] = 12'h777;
rom[31517] = 12'h433;
rom[31518] = 12'h111;
rom[31519] = 12'h  0;
rom[31520] = 12'h  0;
rom[31521] = 12'h  0;
rom[31522] = 12'h  0;
rom[31523] = 12'h  0;
rom[31524] = 12'h  0;
rom[31525] = 12'h  0;
rom[31526] = 12'h  0;
rom[31527] = 12'h  0;
rom[31528] = 12'h  0;
rom[31529] = 12'h  0;
rom[31530] = 12'h  0;
rom[31531] = 12'h  0;
rom[31532] = 12'h100;
rom[31533] = 12'h100;
rom[31534] = 12'h100;
rom[31535] = 12'h100;
rom[31536] = 12'h100;
rom[31537] = 12'h200;
rom[31538] = 12'h200;
rom[31539] = 12'h200;
rom[31540] = 12'h300;
rom[31541] = 12'h300;
rom[31542] = 12'h400;
rom[31543] = 12'h400;
rom[31544] = 12'h610;
rom[31545] = 12'h710;
rom[31546] = 12'h820;
rom[31547] = 12'ha30;
rom[31548] = 12'hc40;
rom[31549] = 12'hd40;
rom[31550] = 12'hd51;
rom[31551] = 12'he50;
rom[31552] = 12'hd50;
rom[31553] = 12'hd60;
rom[31554] = 12'hc60;
rom[31555] = 12'hc60;
rom[31556] = 12'hc71;
rom[31557] = 12'hd82;
rom[31558] = 12'hc82;
rom[31559] = 12'ha71;
rom[31560] = 12'h950;
rom[31561] = 12'h850;
rom[31562] = 12'h840;
rom[31563] = 12'h840;
rom[31564] = 12'h740;
rom[31565] = 12'h740;
rom[31566] = 12'h630;
rom[31567] = 12'h641;
rom[31568] = 12'h641;
rom[31569] = 12'h541;
rom[31570] = 12'h541;
rom[31571] = 12'h541;
rom[31572] = 12'h542;
rom[31573] = 12'h442;
rom[31574] = 12'h543;
rom[31575] = 12'h543;
rom[31576] = 12'h444;
rom[31577] = 12'h554;
rom[31578] = 12'h655;
rom[31579] = 12'h666;
rom[31580] = 12'h666;
rom[31581] = 12'h766;
rom[31582] = 12'h777;
rom[31583] = 12'h777;
rom[31584] = 12'h888;
rom[31585] = 12'h888;
rom[31586] = 12'h888;
rom[31587] = 12'h999;
rom[31588] = 12'h999;
rom[31589] = 12'h999;
rom[31590] = 12'h999;
rom[31591] = 12'h999;
rom[31592] = 12'h999;
rom[31593] = 12'h999;
rom[31594] = 12'haaa;
rom[31595] = 12'haaa;
rom[31596] = 12'haaa;
rom[31597] = 12'haaa;
rom[31598] = 12'hbbb;
rom[31599] = 12'hbbb;
rom[31600] = 12'h777;
rom[31601] = 12'h777;
rom[31602] = 12'h777;
rom[31603] = 12'h777;
rom[31604] = 12'h777;
rom[31605] = 12'h777;
rom[31606] = 12'h777;
rom[31607] = 12'h777;
rom[31608] = 12'h777;
rom[31609] = 12'h777;
rom[31610] = 12'h777;
rom[31611] = 12'h777;
rom[31612] = 12'h777;
rom[31613] = 12'h777;
rom[31614] = 12'h777;
rom[31615] = 12'h777;
rom[31616] = 12'h777;
rom[31617] = 12'h777;
rom[31618] = 12'h777;
rom[31619] = 12'h777;
rom[31620] = 12'h888;
rom[31621] = 12'h888;
rom[31622] = 12'h888;
rom[31623] = 12'h888;
rom[31624] = 12'h777;
rom[31625] = 12'h888;
rom[31626] = 12'h888;
rom[31627] = 12'h888;
rom[31628] = 12'h888;
rom[31629] = 12'h888;
rom[31630] = 12'h888;
rom[31631] = 12'h888;
rom[31632] = 12'h888;
rom[31633] = 12'h888;
rom[31634] = 12'h888;
rom[31635] = 12'h888;
rom[31636] = 12'h888;
rom[31637] = 12'h999;
rom[31638] = 12'h999;
rom[31639] = 12'h999;
rom[31640] = 12'h999;
rom[31641] = 12'h999;
rom[31642] = 12'h888;
rom[31643] = 12'h888;
rom[31644] = 12'h888;
rom[31645] = 12'h777;
rom[31646] = 12'h777;
rom[31647] = 12'h777;
rom[31648] = 12'h666;
rom[31649] = 12'h666;
rom[31650] = 12'h666;
rom[31651] = 12'h666;
rom[31652] = 12'h666;
rom[31653] = 12'h666;
rom[31654] = 12'h666;
rom[31655] = 12'h666;
rom[31656] = 12'h666;
rom[31657] = 12'h666;
rom[31658] = 12'h666;
rom[31659] = 12'h777;
rom[31660] = 12'h777;
rom[31661] = 12'h888;
rom[31662] = 12'h888;
rom[31663] = 12'h999;
rom[31664] = 12'h999;
rom[31665] = 12'h999;
rom[31666] = 12'h999;
rom[31667] = 12'h888;
rom[31668] = 12'h888;
rom[31669] = 12'h777;
rom[31670] = 12'h777;
rom[31671] = 12'h666;
rom[31672] = 12'h666;
rom[31673] = 12'h555;
rom[31674] = 12'h555;
rom[31675] = 12'h555;
rom[31676] = 12'h444;
rom[31677] = 12'h444;
rom[31678] = 12'h444;
rom[31679] = 12'h444;
rom[31680] = 12'h333;
rom[31681] = 12'h333;
rom[31682] = 12'h333;
rom[31683] = 12'h333;
rom[31684] = 12'h333;
rom[31685] = 12'h333;
rom[31686] = 12'h222;
rom[31687] = 12'h222;
rom[31688] = 12'h222;
rom[31689] = 12'h222;
rom[31690] = 12'h222;
rom[31691] = 12'h222;
rom[31692] = 12'h222;
rom[31693] = 12'h111;
rom[31694] = 12'h111;
rom[31695] = 12'h  0;
rom[31696] = 12'h  0;
rom[31697] = 12'h  0;
rom[31698] = 12'h  0;
rom[31699] = 12'h  0;
rom[31700] = 12'h  0;
rom[31701] = 12'h  0;
rom[31702] = 12'h  0;
rom[31703] = 12'h  0;
rom[31704] = 12'h  0;
rom[31705] = 12'h  0;
rom[31706] = 12'h  0;
rom[31707] = 12'h  0;
rom[31708] = 12'h  0;
rom[31709] = 12'h  0;
rom[31710] = 12'h  0;
rom[31711] = 12'h  0;
rom[31712] = 12'h  0;
rom[31713] = 12'h  0;
rom[31714] = 12'h  0;
rom[31715] = 12'h  0;
rom[31716] = 12'h  0;
rom[31717] = 12'h  0;
rom[31718] = 12'h  0;
rom[31719] = 12'h  0;
rom[31720] = 12'h  0;
rom[31721] = 12'h  0;
rom[31722] = 12'h  0;
rom[31723] = 12'h  0;
rom[31724] = 12'h  0;
rom[31725] = 12'h  0;
rom[31726] = 12'h  0;
rom[31727] = 12'h  0;
rom[31728] = 12'h100;
rom[31729] = 12'h100;
rom[31730] = 12'h100;
rom[31731] = 12'h200;
rom[31732] = 12'h200;
rom[31733] = 12'h200;
rom[31734] = 12'h200;
rom[31735] = 12'h200;
rom[31736] = 12'h200;
rom[31737] = 12'h200;
rom[31738] = 12'h200;
rom[31739] = 12'h200;
rom[31740] = 12'h200;
rom[31741] = 12'h200;
rom[31742] = 12'h200;
rom[31743] = 12'h200;
rom[31744] = 12'h300;
rom[31745] = 12'h300;
rom[31746] = 12'h300;
rom[31747] = 12'h300;
rom[31748] = 12'h300;
rom[31749] = 12'h300;
rom[31750] = 12'h200;
rom[31751] = 12'h200;
rom[31752] = 12'h200;
rom[31753] = 12'h200;
rom[31754] = 12'h200;
rom[31755] = 12'h200;
rom[31756] = 12'h200;
rom[31757] = 12'h100;
rom[31758] = 12'h100;
rom[31759] = 12'h100;
rom[31760] = 12'h100;
rom[31761] = 12'h100;
rom[31762] = 12'h100;
rom[31763] = 12'h100;
rom[31764] = 12'h100;
rom[31765] = 12'h  0;
rom[31766] = 12'h  0;
rom[31767] = 12'h  0;
rom[31768] = 12'h  0;
rom[31769] = 12'h  0;
rom[31770] = 12'h  0;
rom[31771] = 12'h  0;
rom[31772] = 12'h  0;
rom[31773] = 12'h  0;
rom[31774] = 12'h  0;
rom[31775] = 12'h  0;
rom[31776] = 12'h  0;
rom[31777] = 12'h  0;
rom[31778] = 12'h  0;
rom[31779] = 12'h  0;
rom[31780] = 12'h  0;
rom[31781] = 12'h  0;
rom[31782] = 12'h  0;
rom[31783] = 12'h  0;
rom[31784] = 12'h  0;
rom[31785] = 12'h  0;
rom[31786] = 12'h  0;
rom[31787] = 12'h  0;
rom[31788] = 12'h  0;
rom[31789] = 12'h  0;
rom[31790] = 12'h  0;
rom[31791] = 12'h  0;
rom[31792] = 12'h  0;
rom[31793] = 12'h  0;
rom[31794] = 12'h  0;
rom[31795] = 12'h  0;
rom[31796] = 12'h  0;
rom[31797] = 12'h111;
rom[31798] = 12'h111;
rom[31799] = 12'h111;
rom[31800] = 12'h111;
rom[31801] = 12'h222;
rom[31802] = 12'h222;
rom[31803] = 12'h333;
rom[31804] = 12'h444;
rom[31805] = 12'h555;
rom[31806] = 12'h666;
rom[31807] = 12'h666;
rom[31808] = 12'h777;
rom[31809] = 12'h777;
rom[31810] = 12'h777;
rom[31811] = 12'h666;
rom[31812] = 12'h666;
rom[31813] = 12'h666;
rom[31814] = 12'h666;
rom[31815] = 12'h666;
rom[31816] = 12'h666;
rom[31817] = 12'h666;
rom[31818] = 12'h666;
rom[31819] = 12'h666;
rom[31820] = 12'h666;
rom[31821] = 12'h666;
rom[31822] = 12'h666;
rom[31823] = 12'h666;
rom[31824] = 12'h666;
rom[31825] = 12'h666;
rom[31826] = 12'h666;
rom[31827] = 12'h666;
rom[31828] = 12'h666;
rom[31829] = 12'h666;
rom[31830] = 12'h666;
rom[31831] = 12'h666;
rom[31832] = 12'h666;
rom[31833] = 12'h666;
rom[31834] = 12'h666;
rom[31835] = 12'h555;
rom[31836] = 12'h555;
rom[31837] = 12'h555;
rom[31838] = 12'h444;
rom[31839] = 12'h333;
rom[31840] = 12'h333;
rom[31841] = 12'h333;
rom[31842] = 12'h222;
rom[31843] = 12'h222;
rom[31844] = 12'h222;
rom[31845] = 12'h222;
rom[31846] = 12'h111;
rom[31847] = 12'h111;
rom[31848] = 12'h111;
rom[31849] = 12'h111;
rom[31850] = 12'h111;
rom[31851] = 12'h  0;
rom[31852] = 12'h  0;
rom[31853] = 12'h  0;
rom[31854] = 12'h111;
rom[31855] = 12'h111;
rom[31856] = 12'h  0;
rom[31857] = 12'h  0;
rom[31858] = 12'h  0;
rom[31859] = 12'h  0;
rom[31860] = 12'h  0;
rom[31861] = 12'h  0;
rom[31862] = 12'h  0;
rom[31863] = 12'h  0;
rom[31864] = 12'h  0;
rom[31865] = 12'h  0;
rom[31866] = 12'h  0;
rom[31867] = 12'h  0;
rom[31868] = 12'h  0;
rom[31869] = 12'h  0;
rom[31870] = 12'h  0;
rom[31871] = 12'h  0;
rom[31872] = 12'h  0;
rom[31873] = 12'h  0;
rom[31874] = 12'h  0;
rom[31875] = 12'h  0;
rom[31876] = 12'h  0;
rom[31877] = 12'h  0;
rom[31878] = 12'h  0;
rom[31879] = 12'h  0;
rom[31880] = 12'h  0;
rom[31881] = 12'h  0;
rom[31882] = 12'h  0;
rom[31883] = 12'h  0;
rom[31884] = 12'h  0;
rom[31885] = 12'h111;
rom[31886] = 12'h111;
rom[31887] = 12'h111;
rom[31888] = 12'h222;
rom[31889] = 12'h222;
rom[31890] = 12'h333;
rom[31891] = 12'h333;
rom[31892] = 12'h333;
rom[31893] = 12'h333;
rom[31894] = 12'h333;
rom[31895] = 12'h333;
rom[31896] = 12'h333;
rom[31897] = 12'h444;
rom[31898] = 12'h555;
rom[31899] = 12'h555;
rom[31900] = 12'h655;
rom[31901] = 12'h766;
rom[31902] = 12'h777;
rom[31903] = 12'h877;
rom[31904] = 12'h888;
rom[31905] = 12'h988;
rom[31906] = 12'h999;
rom[31907] = 12'haaa;
rom[31908] = 12'hbbb;
rom[31909] = 12'hccc;
rom[31910] = 12'heed;
rom[31911] = 12'hfff;
rom[31912] = 12'hfff;
rom[31913] = 12'hedd;
rom[31914] = 12'haaa;
rom[31915] = 12'h766;
rom[31916] = 12'h333;
rom[31917] = 12'h110;
rom[31918] = 12'h100;
rom[31919] = 12'h111;
rom[31920] = 12'h  0;
rom[31921] = 12'h  0;
rom[31922] = 12'h  0;
rom[31923] = 12'h  0;
rom[31924] = 12'h  0;
rom[31925] = 12'h  0;
rom[31926] = 12'h  0;
rom[31927] = 12'h  0;
rom[31928] = 12'h  0;
rom[31929] = 12'h  0;
rom[31930] = 12'h  0;
rom[31931] = 12'h  0;
rom[31932] = 12'h  0;
rom[31933] = 12'h  0;
rom[31934] = 12'h  0;
rom[31935] = 12'h100;
rom[31936] = 12'h100;
rom[31937] = 12'h100;
rom[31938] = 12'h100;
rom[31939] = 12'h200;
rom[31940] = 12'h200;
rom[31941] = 12'h300;
rom[31942] = 12'h400;
rom[31943] = 12'h400;
rom[31944] = 12'h600;
rom[31945] = 12'h710;
rom[31946] = 12'h810;
rom[31947] = 12'ha20;
rom[31948] = 12'hb40;
rom[31949] = 12'hc40;
rom[31950] = 12'hd50;
rom[31951] = 12'hd50;
rom[31952] = 12'hd50;
rom[31953] = 12'hd60;
rom[31954] = 12'hd60;
rom[31955] = 12'hc60;
rom[31956] = 12'hd81;
rom[31957] = 12'hd92;
rom[31958] = 12'hc82;
rom[31959] = 12'ha71;
rom[31960] = 12'h950;
rom[31961] = 12'h850;
rom[31962] = 12'h840;
rom[31963] = 12'h740;
rom[31964] = 12'h740;
rom[31965] = 12'h640;
rom[31966] = 12'h630;
rom[31967] = 12'h641;
rom[31968] = 12'h531;
rom[31969] = 12'h531;
rom[31970] = 12'h531;
rom[31971] = 12'h531;
rom[31972] = 12'h432;
rom[31973] = 12'h432;
rom[31974] = 12'h443;
rom[31975] = 12'h443;
rom[31976] = 12'h443;
rom[31977] = 12'h544;
rom[31978] = 12'h555;
rom[31979] = 12'h666;
rom[31980] = 12'h666;
rom[31981] = 12'h766;
rom[31982] = 12'h777;
rom[31983] = 12'h777;
rom[31984] = 12'h877;
rom[31985] = 12'h888;
rom[31986] = 12'h888;
rom[31987] = 12'h999;
rom[31988] = 12'h999;
rom[31989] = 12'h999;
rom[31990] = 12'h999;
rom[31991] = 12'h999;
rom[31992] = 12'h999;
rom[31993] = 12'h999;
rom[31994] = 12'haaa;
rom[31995] = 12'haaa;
rom[31996] = 12'haaa;
rom[31997] = 12'haaa;
rom[31998] = 12'hbbb;
rom[31999] = 12'hbbb;
rom[32000] = 12'h888;
rom[32001] = 12'h888;
rom[32002] = 12'h888;
rom[32003] = 12'h888;
rom[32004] = 12'h888;
rom[32005] = 12'h888;
rom[32006] = 12'h888;
rom[32007] = 12'h888;
rom[32008] = 12'h888;
rom[32009] = 12'h888;
rom[32010] = 12'h888;
rom[32011] = 12'h888;
rom[32012] = 12'h888;
rom[32013] = 12'h888;
rom[32014] = 12'h888;
rom[32015] = 12'h888;
rom[32016] = 12'h888;
rom[32017] = 12'h888;
rom[32018] = 12'h888;
rom[32019] = 12'h888;
rom[32020] = 12'h888;
rom[32021] = 12'h888;
rom[32022] = 12'h777;
rom[32023] = 12'h777;
rom[32024] = 12'h777;
rom[32025] = 12'h777;
rom[32026] = 12'h888;
rom[32027] = 12'h888;
rom[32028] = 12'h888;
rom[32029] = 12'h888;
rom[32030] = 12'h888;
rom[32031] = 12'h888;
rom[32032] = 12'h888;
rom[32033] = 12'h888;
rom[32034] = 12'h999;
rom[32035] = 12'h999;
rom[32036] = 12'h999;
rom[32037] = 12'h999;
rom[32038] = 12'h999;
rom[32039] = 12'h999;
rom[32040] = 12'h999;
rom[32041] = 12'h999;
rom[32042] = 12'h888;
rom[32043] = 12'h888;
rom[32044] = 12'h888;
rom[32045] = 12'h888;
rom[32046] = 12'h777;
rom[32047] = 12'h777;
rom[32048] = 12'h666;
rom[32049] = 12'h666;
rom[32050] = 12'h666;
rom[32051] = 12'h666;
rom[32052] = 12'h666;
rom[32053] = 12'h666;
rom[32054] = 12'h666;
rom[32055] = 12'h666;
rom[32056] = 12'h666;
rom[32057] = 12'h666;
rom[32058] = 12'h666;
rom[32059] = 12'h666;
rom[32060] = 12'h777;
rom[32061] = 12'h777;
rom[32062] = 12'h888;
rom[32063] = 12'h888;
rom[32064] = 12'h888;
rom[32065] = 12'h999;
rom[32066] = 12'h999;
rom[32067] = 12'h999;
rom[32068] = 12'h888;
rom[32069] = 12'h888;
rom[32070] = 12'h777;
rom[32071] = 12'h666;
rom[32072] = 12'h666;
rom[32073] = 12'h666;
rom[32074] = 12'h555;
rom[32075] = 12'h555;
rom[32076] = 12'h444;
rom[32077] = 12'h444;
rom[32078] = 12'h444;
rom[32079] = 12'h444;
rom[32080] = 12'h333;
rom[32081] = 12'h333;
rom[32082] = 12'h333;
rom[32083] = 12'h333;
rom[32084] = 12'h333;
rom[32085] = 12'h333;
rom[32086] = 12'h222;
rom[32087] = 12'h222;
rom[32088] = 12'h222;
rom[32089] = 12'h222;
rom[32090] = 12'h222;
rom[32091] = 12'h222;
rom[32092] = 12'h222;
rom[32093] = 12'h111;
rom[32094] = 12'h111;
rom[32095] = 12'h111;
rom[32096] = 12'h  0;
rom[32097] = 12'h  0;
rom[32098] = 12'h  0;
rom[32099] = 12'h  0;
rom[32100] = 12'h  0;
rom[32101] = 12'h  0;
rom[32102] = 12'h  0;
rom[32103] = 12'h  0;
rom[32104] = 12'h  0;
rom[32105] = 12'h  0;
rom[32106] = 12'h  0;
rom[32107] = 12'h  0;
rom[32108] = 12'h  0;
rom[32109] = 12'h  0;
rom[32110] = 12'h  0;
rom[32111] = 12'h  0;
rom[32112] = 12'h  0;
rom[32113] = 12'h  0;
rom[32114] = 12'h  0;
rom[32115] = 12'h  0;
rom[32116] = 12'h  0;
rom[32117] = 12'h  0;
rom[32118] = 12'h  0;
rom[32119] = 12'h  0;
rom[32120] = 12'h  0;
rom[32121] = 12'h  0;
rom[32122] = 12'h  0;
rom[32123] = 12'h  0;
rom[32124] = 12'h  0;
rom[32125] = 12'h  0;
rom[32126] = 12'h  0;
rom[32127] = 12'h  0;
rom[32128] = 12'h  0;
rom[32129] = 12'h100;
rom[32130] = 12'h100;
rom[32131] = 12'h100;
rom[32132] = 12'h100;
rom[32133] = 12'h100;
rom[32134] = 12'h100;
rom[32135] = 12'h100;
rom[32136] = 12'h100;
rom[32137] = 12'h100;
rom[32138] = 12'h100;
rom[32139] = 12'h200;
rom[32140] = 12'h200;
rom[32141] = 12'h200;
rom[32142] = 12'h200;
rom[32143] = 12'h200;
rom[32144] = 12'h200;
rom[32145] = 12'h200;
rom[32146] = 12'h200;
rom[32147] = 12'h200;
rom[32148] = 12'h200;
rom[32149] = 12'h200;
rom[32150] = 12'h200;
rom[32151] = 12'h200;
rom[32152] = 12'h200;
rom[32153] = 12'h100;
rom[32154] = 12'h100;
rom[32155] = 12'h100;
rom[32156] = 12'h100;
rom[32157] = 12'h100;
rom[32158] = 12'h100;
rom[32159] = 12'h100;
rom[32160] = 12'h  0;
rom[32161] = 12'h  0;
rom[32162] = 12'h  0;
rom[32163] = 12'h  0;
rom[32164] = 12'h  0;
rom[32165] = 12'h  0;
rom[32166] = 12'h  0;
rom[32167] = 12'h  0;
rom[32168] = 12'h  0;
rom[32169] = 12'h  0;
rom[32170] = 12'h  0;
rom[32171] = 12'h  0;
rom[32172] = 12'h  0;
rom[32173] = 12'h  0;
rom[32174] = 12'h  0;
rom[32175] = 12'h  0;
rom[32176] = 12'h  0;
rom[32177] = 12'h  0;
rom[32178] = 12'h  0;
rom[32179] = 12'h  0;
rom[32180] = 12'h  0;
rom[32181] = 12'h  0;
rom[32182] = 12'h  0;
rom[32183] = 12'h  0;
rom[32184] = 12'h  0;
rom[32185] = 12'h  0;
rom[32186] = 12'h  0;
rom[32187] = 12'h  0;
rom[32188] = 12'h  0;
rom[32189] = 12'h  0;
rom[32190] = 12'h  0;
rom[32191] = 12'h  0;
rom[32192] = 12'h  0;
rom[32193] = 12'h  0;
rom[32194] = 12'h  0;
rom[32195] = 12'h  0;
rom[32196] = 12'h  0;
rom[32197] = 12'h111;
rom[32198] = 12'h111;
rom[32199] = 12'h111;
rom[32200] = 12'h222;
rom[32201] = 12'h222;
rom[32202] = 12'h333;
rom[32203] = 12'h333;
rom[32204] = 12'h444;
rom[32205] = 12'h555;
rom[32206] = 12'h555;
rom[32207] = 12'h555;
rom[32208] = 12'h777;
rom[32209] = 12'h777;
rom[32210] = 12'h666;
rom[32211] = 12'h666;
rom[32212] = 12'h666;
rom[32213] = 12'h666;
rom[32214] = 12'h666;
rom[32215] = 12'h555;
rom[32216] = 12'h555;
rom[32217] = 12'h555;
rom[32218] = 12'h555;
rom[32219] = 12'h666;
rom[32220] = 12'h666;
rom[32221] = 12'h666;
rom[32222] = 12'h666;
rom[32223] = 12'h666;
rom[32224] = 12'h666;
rom[32225] = 12'h666;
rom[32226] = 12'h666;
rom[32227] = 12'h666;
rom[32228] = 12'h555;
rom[32229] = 12'h666;
rom[32230] = 12'h666;
rom[32231] = 12'h777;
rom[32232] = 12'h666;
rom[32233] = 12'h666;
rom[32234] = 12'h666;
rom[32235] = 12'h555;
rom[32236] = 12'h555;
rom[32237] = 12'h444;
rom[32238] = 12'h444;
rom[32239] = 12'h333;
rom[32240] = 12'h333;
rom[32241] = 12'h333;
rom[32242] = 12'h222;
rom[32243] = 12'h222;
rom[32244] = 12'h222;
rom[32245] = 12'h222;
rom[32246] = 12'h111;
rom[32247] = 12'h111;
rom[32248] = 12'h  0;
rom[32249] = 12'h  0;
rom[32250] = 12'h  0;
rom[32251] = 12'h111;
rom[32252] = 12'h111;
rom[32253] = 12'h111;
rom[32254] = 12'h  0;
rom[32255] = 12'h  0;
rom[32256] = 12'h  0;
rom[32257] = 12'h  0;
rom[32258] = 12'h  0;
rom[32259] = 12'h  0;
rom[32260] = 12'h  0;
rom[32261] = 12'h  0;
rom[32262] = 12'h  0;
rom[32263] = 12'h  0;
rom[32264] = 12'h  0;
rom[32265] = 12'h  0;
rom[32266] = 12'h  0;
rom[32267] = 12'h  0;
rom[32268] = 12'h  0;
rom[32269] = 12'h  0;
rom[32270] = 12'h  0;
rom[32271] = 12'h  0;
rom[32272] = 12'h  0;
rom[32273] = 12'h  0;
rom[32274] = 12'h  0;
rom[32275] = 12'h  0;
rom[32276] = 12'h  0;
rom[32277] = 12'h  0;
rom[32278] = 12'h  0;
rom[32279] = 12'h  0;
rom[32280] = 12'h  0;
rom[32281] = 12'h  0;
rom[32282] = 12'h  0;
rom[32283] = 12'h  0;
rom[32284] = 12'h  0;
rom[32285] = 12'h111;
rom[32286] = 12'h111;
rom[32287] = 12'h111;
rom[32288] = 12'h222;
rom[32289] = 12'h222;
rom[32290] = 12'h333;
rom[32291] = 12'h333;
rom[32292] = 12'h333;
rom[32293] = 12'h333;
rom[32294] = 12'h333;
rom[32295] = 12'h333;
rom[32296] = 12'h444;
rom[32297] = 12'h444;
rom[32298] = 12'h555;
rom[32299] = 12'h655;
rom[32300] = 12'h766;
rom[32301] = 12'h867;
rom[32302] = 12'h877;
rom[32303] = 12'h888;
rom[32304] = 12'h988;
rom[32305] = 12'h999;
rom[32306] = 12'haaa;
rom[32307] = 12'hbbb;
rom[32308] = 12'hddc;
rom[32309] = 12'hded;
rom[32310] = 12'heee;
rom[32311] = 12'hffe;
rom[32312] = 12'heed;
rom[32313] = 12'haa9;
rom[32314] = 12'h554;
rom[32315] = 12'h222;
rom[32316] = 12'h110;
rom[32317] = 12'h100;
rom[32318] = 12'h100;
rom[32319] = 12'h100;
rom[32320] = 12'h  0;
rom[32321] = 12'h  0;
rom[32322] = 12'h  0;
rom[32323] = 12'h  0;
rom[32324] = 12'h  0;
rom[32325] = 12'h  0;
rom[32326] = 12'h  0;
rom[32327] = 12'h  0;
rom[32328] = 12'h  0;
rom[32329] = 12'h  0;
rom[32330] = 12'h  0;
rom[32331] = 12'h  0;
rom[32332] = 12'h  0;
rom[32333] = 12'h  0;
rom[32334] = 12'h  0;
rom[32335] = 12'h100;
rom[32336] = 12'h100;
rom[32337] = 12'h100;
rom[32338] = 12'h100;
rom[32339] = 12'h200;
rom[32340] = 12'h300;
rom[32341] = 12'h300;
rom[32342] = 12'h400;
rom[32343] = 12'h500;
rom[32344] = 12'h600;
rom[32345] = 12'h710;
rom[32346] = 12'h810;
rom[32347] = 12'ha30;
rom[32348] = 12'hc40;
rom[32349] = 12'hd50;
rom[32350] = 12'hd50;
rom[32351] = 12'he50;
rom[32352] = 12'he60;
rom[32353] = 12'hd60;
rom[32354] = 12'hd60;
rom[32355] = 12'he81;
rom[32356] = 12'he92;
rom[32357] = 12'he93;
rom[32358] = 12'hc81;
rom[32359] = 12'ha71;
rom[32360] = 12'h950;
rom[32361] = 12'h850;
rom[32362] = 12'h850;
rom[32363] = 12'h740;
rom[32364] = 12'h740;
rom[32365] = 12'h641;
rom[32366] = 12'h541;
rom[32367] = 12'h531;
rom[32368] = 12'h531;
rom[32369] = 12'h531;
rom[32370] = 12'h431;
rom[32371] = 12'h431;
rom[32372] = 12'h431;
rom[32373] = 12'h432;
rom[32374] = 12'h432;
rom[32375] = 12'h433;
rom[32376] = 12'h433;
rom[32377] = 12'h444;
rom[32378] = 12'h545;
rom[32379] = 12'h655;
rom[32380] = 12'h656;
rom[32381] = 12'h766;
rom[32382] = 12'h777;
rom[32383] = 12'h877;
rom[32384] = 12'h777;
rom[32385] = 12'h777;
rom[32386] = 12'h888;
rom[32387] = 12'h888;
rom[32388] = 12'h999;
rom[32389] = 12'h999;
rom[32390] = 12'h999;
rom[32391] = 12'h999;
rom[32392] = 12'h999;
rom[32393] = 12'h999;
rom[32394] = 12'haaa;
rom[32395] = 12'haaa;
rom[32396] = 12'haaa;
rom[32397] = 12'haaa;
rom[32398] = 12'hbbb;
rom[32399] = 12'hbbb;
rom[32400] = 12'h999;
rom[32401] = 12'h999;
rom[32402] = 12'h999;
rom[32403] = 12'h999;
rom[32404] = 12'h888;
rom[32405] = 12'h888;
rom[32406] = 12'h888;
rom[32407] = 12'h888;
rom[32408] = 12'h888;
rom[32409] = 12'h888;
rom[32410] = 12'h888;
rom[32411] = 12'h888;
rom[32412] = 12'h888;
rom[32413] = 12'h888;
rom[32414] = 12'h888;
rom[32415] = 12'h888;
rom[32416] = 12'h888;
rom[32417] = 12'h888;
rom[32418] = 12'h888;
rom[32419] = 12'h888;
rom[32420] = 12'h888;
rom[32421] = 12'h888;
rom[32422] = 12'h888;
rom[32423] = 12'h777;
rom[32424] = 12'h777;
rom[32425] = 12'h777;
rom[32426] = 12'h888;
rom[32427] = 12'h888;
rom[32428] = 12'h888;
rom[32429] = 12'h888;
rom[32430] = 12'h888;
rom[32431] = 12'h999;
rom[32432] = 12'h888;
rom[32433] = 12'h888;
rom[32434] = 12'h999;
rom[32435] = 12'h999;
rom[32436] = 12'h999;
rom[32437] = 12'h999;
rom[32438] = 12'h999;
rom[32439] = 12'h999;
rom[32440] = 12'h999;
rom[32441] = 12'h999;
rom[32442] = 12'h999;
rom[32443] = 12'h888;
rom[32444] = 12'h888;
rom[32445] = 12'h888;
rom[32446] = 12'h777;
rom[32447] = 12'h777;
rom[32448] = 12'h777;
rom[32449] = 12'h666;
rom[32450] = 12'h666;
rom[32451] = 12'h666;
rom[32452] = 12'h666;
rom[32453] = 12'h777;
rom[32454] = 12'h666;
rom[32455] = 12'h666;
rom[32456] = 12'h666;
rom[32457] = 12'h666;
rom[32458] = 12'h666;
rom[32459] = 12'h666;
rom[32460] = 12'h666;
rom[32461] = 12'h777;
rom[32462] = 12'h777;
rom[32463] = 12'h777;
rom[32464] = 12'h888;
rom[32465] = 12'h999;
rom[32466] = 12'h999;
rom[32467] = 12'h999;
rom[32468] = 12'h999;
rom[32469] = 12'h888;
rom[32470] = 12'h777;
rom[32471] = 12'h777;
rom[32472] = 12'h666;
rom[32473] = 12'h666;
rom[32474] = 12'h555;
rom[32475] = 12'h555;
rom[32476] = 12'h555;
rom[32477] = 12'h444;
rom[32478] = 12'h444;
rom[32479] = 12'h444;
rom[32480] = 12'h333;
rom[32481] = 12'h333;
rom[32482] = 12'h333;
rom[32483] = 12'h333;
rom[32484] = 12'h333;
rom[32485] = 12'h333;
rom[32486] = 12'h333;
rom[32487] = 12'h222;
rom[32488] = 12'h222;
rom[32489] = 12'h222;
rom[32490] = 12'h222;
rom[32491] = 12'h222;
rom[32492] = 12'h222;
rom[32493] = 12'h111;
rom[32494] = 12'h111;
rom[32495] = 12'h111;
rom[32496] = 12'h  0;
rom[32497] = 12'h  0;
rom[32498] = 12'h  0;
rom[32499] = 12'h  0;
rom[32500] = 12'h  0;
rom[32501] = 12'h  0;
rom[32502] = 12'h  0;
rom[32503] = 12'h  0;
rom[32504] = 12'h  0;
rom[32505] = 12'h  0;
rom[32506] = 12'h  0;
rom[32507] = 12'h  0;
rom[32508] = 12'h  0;
rom[32509] = 12'h  0;
rom[32510] = 12'h  0;
rom[32511] = 12'h  0;
rom[32512] = 12'h  0;
rom[32513] = 12'h  0;
rom[32514] = 12'h  0;
rom[32515] = 12'h  0;
rom[32516] = 12'h  0;
rom[32517] = 12'h  0;
rom[32518] = 12'h  0;
rom[32519] = 12'h  0;
rom[32520] = 12'h  0;
rom[32521] = 12'h  0;
rom[32522] = 12'h  0;
rom[32523] = 12'h  0;
rom[32524] = 12'h  0;
rom[32525] = 12'h  0;
rom[32526] = 12'h  0;
rom[32527] = 12'h  0;
rom[32528] = 12'h  0;
rom[32529] = 12'h  0;
rom[32530] = 12'h  0;
rom[32531] = 12'h  0;
rom[32532] = 12'h  0;
rom[32533] = 12'h  0;
rom[32534] = 12'h  0;
rom[32535] = 12'h100;
rom[32536] = 12'h100;
rom[32537] = 12'h100;
rom[32538] = 12'h100;
rom[32539] = 12'h100;
rom[32540] = 12'h100;
rom[32541] = 12'h100;
rom[32542] = 12'h100;
rom[32543] = 12'h200;
rom[32544] = 12'h200;
rom[32545] = 12'h200;
rom[32546] = 12'h200;
rom[32547] = 12'h200;
rom[32548] = 12'h200;
rom[32549] = 12'h200;
rom[32550] = 12'h200;
rom[32551] = 12'h200;
rom[32552] = 12'h100;
rom[32553] = 12'h100;
rom[32554] = 12'h100;
rom[32555] = 12'h100;
rom[32556] = 12'h100;
rom[32557] = 12'h100;
rom[32558] = 12'h100;
rom[32559] = 12'h100;
rom[32560] = 12'h  0;
rom[32561] = 12'h  0;
rom[32562] = 12'h  0;
rom[32563] = 12'h  0;
rom[32564] = 12'h  0;
rom[32565] = 12'h  0;
rom[32566] = 12'h  0;
rom[32567] = 12'h  0;
rom[32568] = 12'h  0;
rom[32569] = 12'h  0;
rom[32570] = 12'h  0;
rom[32571] = 12'h  0;
rom[32572] = 12'h  0;
rom[32573] = 12'h  0;
rom[32574] = 12'h  0;
rom[32575] = 12'h  0;
rom[32576] = 12'h  0;
rom[32577] = 12'h  0;
rom[32578] = 12'h  0;
rom[32579] = 12'h  0;
rom[32580] = 12'h  0;
rom[32581] = 12'h  0;
rom[32582] = 12'h  0;
rom[32583] = 12'h  0;
rom[32584] = 12'h  0;
rom[32585] = 12'h  0;
rom[32586] = 12'h  0;
rom[32587] = 12'h  0;
rom[32588] = 12'h  0;
rom[32589] = 12'h  0;
rom[32590] = 12'h  0;
rom[32591] = 12'h  0;
rom[32592] = 12'h  0;
rom[32593] = 12'h  0;
rom[32594] = 12'h  0;
rom[32595] = 12'h  0;
rom[32596] = 12'h  0;
rom[32597] = 12'h111;
rom[32598] = 12'h111;
rom[32599] = 12'h111;
rom[32600] = 12'h222;
rom[32601] = 12'h222;
rom[32602] = 12'h333;
rom[32603] = 12'h444;
rom[32604] = 12'h444;
rom[32605] = 12'h555;
rom[32606] = 12'h555;
rom[32607] = 12'h555;
rom[32608] = 12'h666;
rom[32609] = 12'h777;
rom[32610] = 12'h666;
rom[32611] = 12'h666;
rom[32612] = 12'h666;
rom[32613] = 12'h666;
rom[32614] = 12'h666;
rom[32615] = 12'h555;
rom[32616] = 12'h555;
rom[32617] = 12'h555;
rom[32618] = 12'h555;
rom[32619] = 12'h555;
rom[32620] = 12'h555;
rom[32621] = 12'h555;
rom[32622] = 12'h555;
rom[32623] = 12'h555;
rom[32624] = 12'h666;
rom[32625] = 12'h666;
rom[32626] = 12'h666;
rom[32627] = 12'h555;
rom[32628] = 12'h555;
rom[32629] = 12'h666;
rom[32630] = 12'h666;
rom[32631] = 12'h666;
rom[32632] = 12'h666;
rom[32633] = 12'h666;
rom[32634] = 12'h666;
rom[32635] = 12'h555;
rom[32636] = 12'h555;
rom[32637] = 12'h444;
rom[32638] = 12'h444;
rom[32639] = 12'h333;
rom[32640] = 12'h333;
rom[32641] = 12'h333;
rom[32642] = 12'h222;
rom[32643] = 12'h222;
rom[32644] = 12'h222;
rom[32645] = 12'h222;
rom[32646] = 12'h111;
rom[32647] = 12'h111;
rom[32648] = 12'h111;
rom[32649] = 12'h111;
rom[32650] = 12'h111;
rom[32651] = 12'h111;
rom[32652] = 12'h111;
rom[32653] = 12'h111;
rom[32654] = 12'h  0;
rom[32655] = 12'h  0;
rom[32656] = 12'h  0;
rom[32657] = 12'h  0;
rom[32658] = 12'h  0;
rom[32659] = 12'h  0;
rom[32660] = 12'h  0;
rom[32661] = 12'h  0;
rom[32662] = 12'h  0;
rom[32663] = 12'h  0;
rom[32664] = 12'h  0;
rom[32665] = 12'h  0;
rom[32666] = 12'h  0;
rom[32667] = 12'h  0;
rom[32668] = 12'h  0;
rom[32669] = 12'h  0;
rom[32670] = 12'h  0;
rom[32671] = 12'h  0;
rom[32672] = 12'h  0;
rom[32673] = 12'h  0;
rom[32674] = 12'h  0;
rom[32675] = 12'h  0;
rom[32676] = 12'h  0;
rom[32677] = 12'h  0;
rom[32678] = 12'h  0;
rom[32679] = 12'h  0;
rom[32680] = 12'h  0;
rom[32681] = 12'h  0;
rom[32682] = 12'h  0;
rom[32683] = 12'h  0;
rom[32684] = 12'h  0;
rom[32685] = 12'h111;
rom[32686] = 12'h111;
rom[32687] = 12'h222;
rom[32688] = 12'h222;
rom[32689] = 12'h322;
rom[32690] = 12'h333;
rom[32691] = 12'h333;
rom[32692] = 12'h333;
rom[32693] = 12'h333;
rom[32694] = 12'h333;
rom[32695] = 12'h333;
rom[32696] = 12'h444;
rom[32697] = 12'h544;
rom[32698] = 12'h655;
rom[32699] = 12'h666;
rom[32700] = 12'h767;
rom[32701] = 12'h877;
rom[32702] = 12'h978;
rom[32703] = 12'h988;
rom[32704] = 12'h999;
rom[32705] = 12'haaa;
rom[32706] = 12'hcbb;
rom[32707] = 12'hccc;
rom[32708] = 12'hedd;
rom[32709] = 12'hffe;
rom[32710] = 12'hffe;
rom[32711] = 12'heed;
rom[32712] = 12'h998;
rom[32713] = 12'h665;
rom[32714] = 12'h222;
rom[32715] = 12'h110;
rom[32716] = 12'h100;
rom[32717] = 12'h100;
rom[32718] = 12'h  0;
rom[32719] = 12'h  0;
rom[32720] = 12'h  0;
rom[32721] = 12'h  0;
rom[32722] = 12'h  0;
rom[32723] = 12'h  0;
rom[32724] = 12'h  0;
rom[32725] = 12'h  0;
rom[32726] = 12'h  0;
rom[32727] = 12'h  0;
rom[32728] = 12'h  0;
rom[32729] = 12'h  0;
rom[32730] = 12'h  0;
rom[32731] = 12'h  0;
rom[32732] = 12'h  0;
rom[32733] = 12'h  0;
rom[32734] = 12'h  0;
rom[32735] = 12'h  0;
rom[32736] = 12'h100;
rom[32737] = 12'h100;
rom[32738] = 12'h100;
rom[32739] = 12'h200;
rom[32740] = 12'h200;
rom[32741] = 12'h300;
rom[32742] = 12'h400;
rom[32743] = 12'h500;
rom[32744] = 12'h600;
rom[32745] = 12'h700;
rom[32746] = 12'h810;
rom[32747] = 12'ha20;
rom[32748] = 12'hc40;
rom[32749] = 12'hd50;
rom[32750] = 12'hd50;
rom[32751] = 12'he50;
rom[32752] = 12'he60;
rom[32753] = 12'hd60;
rom[32754] = 12'hd60;
rom[32755] = 12'he81;
rom[32756] = 12'hf93;
rom[32757] = 12'he93;
rom[32758] = 12'hc81;
rom[32759] = 12'ha60;
rom[32760] = 12'h950;
rom[32761] = 12'h850;
rom[32762] = 12'h850;
rom[32763] = 12'h740;
rom[32764] = 12'h640;
rom[32765] = 12'h530;
rom[32766] = 12'h530;
rom[32767] = 12'h531;
rom[32768] = 12'h431;
rom[32769] = 12'h421;
rom[32770] = 12'h421;
rom[32771] = 12'h421;
rom[32772] = 12'h421;
rom[32773] = 12'h322;
rom[32774] = 12'h322;
rom[32775] = 12'h332;
rom[32776] = 12'h433;
rom[32777] = 12'h433;
rom[32778] = 12'h444;
rom[32779] = 12'h555;
rom[32780] = 12'h656;
rom[32781] = 12'h766;
rom[32782] = 12'h767;
rom[32783] = 12'h777;
rom[32784] = 12'h777;
rom[32785] = 12'h777;
rom[32786] = 12'h888;
rom[32787] = 12'h888;
rom[32788] = 12'h999;
rom[32789] = 12'h999;
rom[32790] = 12'h999;
rom[32791] = 12'h999;
rom[32792] = 12'h999;
rom[32793] = 12'h999;
rom[32794] = 12'haaa;
rom[32795] = 12'haaa;
rom[32796] = 12'haaa;
rom[32797] = 12'haaa;
rom[32798] = 12'hbbb;
rom[32799] = 12'hbbb;
rom[32800] = 12'h999;
rom[32801] = 12'h999;
rom[32802] = 12'h999;
rom[32803] = 12'h999;
rom[32804] = 12'h999;
rom[32805] = 12'h999;
rom[32806] = 12'h888;
rom[32807] = 12'h888;
rom[32808] = 12'h888;
rom[32809] = 12'h888;
rom[32810] = 12'h888;
rom[32811] = 12'h888;
rom[32812] = 12'h888;
rom[32813] = 12'h888;
rom[32814] = 12'h888;
rom[32815] = 12'h888;
rom[32816] = 12'h888;
rom[32817] = 12'h888;
rom[32818] = 12'h888;
rom[32819] = 12'h888;
rom[32820] = 12'h888;
rom[32821] = 12'h888;
rom[32822] = 12'h888;
rom[32823] = 12'h888;
rom[32824] = 12'h888;
rom[32825] = 12'h888;
rom[32826] = 12'h888;
rom[32827] = 12'h888;
rom[32828] = 12'h888;
rom[32829] = 12'h888;
rom[32830] = 12'h888;
rom[32831] = 12'h888;
rom[32832] = 12'h888;
rom[32833] = 12'h888;
rom[32834] = 12'h999;
rom[32835] = 12'h999;
rom[32836] = 12'h999;
rom[32837] = 12'h999;
rom[32838] = 12'h999;
rom[32839] = 12'h999;
rom[32840] = 12'h999;
rom[32841] = 12'h999;
rom[32842] = 12'h999;
rom[32843] = 12'h999;
rom[32844] = 12'h888;
rom[32845] = 12'h888;
rom[32846] = 12'h888;
rom[32847] = 12'h777;
rom[32848] = 12'h777;
rom[32849] = 12'h777;
rom[32850] = 12'h666;
rom[32851] = 12'h666;
rom[32852] = 12'h777;
rom[32853] = 12'h777;
rom[32854] = 12'h777;
rom[32855] = 12'h666;
rom[32856] = 12'h666;
rom[32857] = 12'h666;
rom[32858] = 12'h666;
rom[32859] = 12'h666;
rom[32860] = 12'h666;
rom[32861] = 12'h666;
rom[32862] = 12'h666;
rom[32863] = 12'h777;
rom[32864] = 12'h888;
rom[32865] = 12'h888;
rom[32866] = 12'h999;
rom[32867] = 12'h999;
rom[32868] = 12'h999;
rom[32869] = 12'h999;
rom[32870] = 12'h888;
rom[32871] = 12'h888;
rom[32872] = 12'h777;
rom[32873] = 12'h777;
rom[32874] = 12'h666;
rom[32875] = 12'h555;
rom[32876] = 12'h555;
rom[32877] = 12'h555;
rom[32878] = 12'h444;
rom[32879] = 12'h444;
rom[32880] = 12'h444;
rom[32881] = 12'h444;
rom[32882] = 12'h333;
rom[32883] = 12'h333;
rom[32884] = 12'h333;
rom[32885] = 12'h333;
rom[32886] = 12'h333;
rom[32887] = 12'h222;
rom[32888] = 12'h222;
rom[32889] = 12'h222;
rom[32890] = 12'h222;
rom[32891] = 12'h222;
rom[32892] = 12'h222;
rom[32893] = 12'h222;
rom[32894] = 12'h111;
rom[32895] = 12'h111;
rom[32896] = 12'h  0;
rom[32897] = 12'h  0;
rom[32898] = 12'h  0;
rom[32899] = 12'h  0;
rom[32900] = 12'h  0;
rom[32901] = 12'h  0;
rom[32902] = 12'h  0;
rom[32903] = 12'h  0;
rom[32904] = 12'h  0;
rom[32905] = 12'h  0;
rom[32906] = 12'h  0;
rom[32907] = 12'h  0;
rom[32908] = 12'h  0;
rom[32909] = 12'h  0;
rom[32910] = 12'h  0;
rom[32911] = 12'h  0;
rom[32912] = 12'h  0;
rom[32913] = 12'h  0;
rom[32914] = 12'h  0;
rom[32915] = 12'h  0;
rom[32916] = 12'h  0;
rom[32917] = 12'h  0;
rom[32918] = 12'h  0;
rom[32919] = 12'h  0;
rom[32920] = 12'h  0;
rom[32921] = 12'h  0;
rom[32922] = 12'h  0;
rom[32923] = 12'h  0;
rom[32924] = 12'h  0;
rom[32925] = 12'h  0;
rom[32926] = 12'h  0;
rom[32927] = 12'h  0;
rom[32928] = 12'h  0;
rom[32929] = 12'h  0;
rom[32930] = 12'h  0;
rom[32931] = 12'h  0;
rom[32932] = 12'h  0;
rom[32933] = 12'h  0;
rom[32934] = 12'h  0;
rom[32935] = 12'h  0;
rom[32936] = 12'h100;
rom[32937] = 12'h100;
rom[32938] = 12'h100;
rom[32939] = 12'h100;
rom[32940] = 12'h100;
rom[32941] = 12'h100;
rom[32942] = 12'h100;
rom[32943] = 12'h100;
rom[32944] = 12'h200;
rom[32945] = 12'h200;
rom[32946] = 12'h200;
rom[32947] = 12'h200;
rom[32948] = 12'h200;
rom[32949] = 12'h200;
rom[32950] = 12'h100;
rom[32951] = 12'h100;
rom[32952] = 12'h100;
rom[32953] = 12'h100;
rom[32954] = 12'h100;
rom[32955] = 12'h100;
rom[32956] = 12'h100;
rom[32957] = 12'h100;
rom[32958] = 12'h100;
rom[32959] = 12'h  0;
rom[32960] = 12'h  0;
rom[32961] = 12'h  0;
rom[32962] = 12'h  0;
rom[32963] = 12'h  0;
rom[32964] = 12'h  0;
rom[32965] = 12'h  0;
rom[32966] = 12'h  0;
rom[32967] = 12'h  0;
rom[32968] = 12'h  0;
rom[32969] = 12'h  0;
rom[32970] = 12'h  0;
rom[32971] = 12'h  0;
rom[32972] = 12'h  0;
rom[32973] = 12'h  0;
rom[32974] = 12'h  0;
rom[32975] = 12'h  0;
rom[32976] = 12'h  0;
rom[32977] = 12'h  0;
rom[32978] = 12'h  0;
rom[32979] = 12'h  0;
rom[32980] = 12'h  0;
rom[32981] = 12'h  0;
rom[32982] = 12'h  0;
rom[32983] = 12'h  0;
rom[32984] = 12'h  0;
rom[32985] = 12'h  0;
rom[32986] = 12'h  0;
rom[32987] = 12'h  0;
rom[32988] = 12'h  0;
rom[32989] = 12'h  0;
rom[32990] = 12'h  0;
rom[32991] = 12'h  0;
rom[32992] = 12'h  0;
rom[32993] = 12'h  0;
rom[32994] = 12'h  0;
rom[32995] = 12'h  0;
rom[32996] = 12'h  0;
rom[32997] = 12'h  0;
rom[32998] = 12'h111;
rom[32999] = 12'h111;
rom[33000] = 12'h222;
rom[33001] = 12'h222;
rom[33002] = 12'h333;
rom[33003] = 12'h444;
rom[33004] = 12'h444;
rom[33005] = 12'h555;
rom[33006] = 12'h555;
rom[33007] = 12'h555;
rom[33008] = 12'h666;
rom[33009] = 12'h666;
rom[33010] = 12'h666;
rom[33011] = 12'h666;
rom[33012] = 12'h666;
rom[33013] = 12'h666;
rom[33014] = 12'h666;
rom[33015] = 12'h555;
rom[33016] = 12'h555;
rom[33017] = 12'h555;
rom[33018] = 12'h555;
rom[33019] = 12'h555;
rom[33020] = 12'h555;
rom[33021] = 12'h555;
rom[33022] = 12'h555;
rom[33023] = 12'h555;
rom[33024] = 12'h555;
rom[33025] = 12'h555;
rom[33026] = 12'h555;
rom[33027] = 12'h555;
rom[33028] = 12'h555;
rom[33029] = 12'h555;
rom[33030] = 12'h666;
rom[33031] = 12'h666;
rom[33032] = 12'h666;
rom[33033] = 12'h666;
rom[33034] = 12'h555;
rom[33035] = 12'h555;
rom[33036] = 12'h555;
rom[33037] = 12'h444;
rom[33038] = 12'h333;
rom[33039] = 12'h333;
rom[33040] = 12'h333;
rom[33041] = 12'h333;
rom[33042] = 12'h222;
rom[33043] = 12'h222;
rom[33044] = 12'h222;
rom[33045] = 12'h111;
rom[33046] = 12'h111;
rom[33047] = 12'h111;
rom[33048] = 12'h111;
rom[33049] = 12'h111;
rom[33050] = 12'h111;
rom[33051] = 12'h111;
rom[33052] = 12'h111;
rom[33053] = 12'h111;
rom[33054] = 12'h  0;
rom[33055] = 12'h  0;
rom[33056] = 12'h  0;
rom[33057] = 12'h  0;
rom[33058] = 12'h  0;
rom[33059] = 12'h  0;
rom[33060] = 12'h  0;
rom[33061] = 12'h  0;
rom[33062] = 12'h  0;
rom[33063] = 12'h  0;
rom[33064] = 12'h  0;
rom[33065] = 12'h  0;
rom[33066] = 12'h  0;
rom[33067] = 12'h  0;
rom[33068] = 12'h  0;
rom[33069] = 12'h  0;
rom[33070] = 12'h  0;
rom[33071] = 12'h  0;
rom[33072] = 12'h  0;
rom[33073] = 12'h  0;
rom[33074] = 12'h  0;
rom[33075] = 12'h  0;
rom[33076] = 12'h  0;
rom[33077] = 12'h  0;
rom[33078] = 12'h  0;
rom[33079] = 12'h  0;
rom[33080] = 12'h  0;
rom[33081] = 12'h  0;
rom[33082] = 12'h  0;
rom[33083] = 12'h  0;
rom[33084] = 12'h  0;
rom[33085] = 12'h111;
rom[33086] = 12'h111;
rom[33087] = 12'h222;
rom[33088] = 12'h333;
rom[33089] = 12'h333;
rom[33090] = 12'h333;
rom[33091] = 12'h333;
rom[33092] = 12'h333;
rom[33093] = 12'h333;
rom[33094] = 12'h333;
rom[33095] = 12'h444;
rom[33096] = 12'h444;
rom[33097] = 12'h555;
rom[33098] = 12'h656;
rom[33099] = 12'h766;
rom[33100] = 12'h877;
rom[33101] = 12'h878;
rom[33102] = 12'h988;
rom[33103] = 12'ha99;
rom[33104] = 12'haaa;
rom[33105] = 12'hcbb;
rom[33106] = 12'hdcc;
rom[33107] = 12'hddd;
rom[33108] = 12'hffe;
rom[33109] = 12'hfff;
rom[33110] = 12'heed;
rom[33111] = 12'hbba;
rom[33112] = 12'h443;
rom[33113] = 12'h221;
rom[33114] = 12'h  0;
rom[33115] = 12'h  0;
rom[33116] = 12'h100;
rom[33117] = 12'h100;
rom[33118] = 12'h100;
rom[33119] = 12'h  0;
rom[33120] = 12'h  0;
rom[33121] = 12'h  0;
rom[33122] = 12'h  0;
rom[33123] = 12'h  0;
rom[33124] = 12'h  0;
rom[33125] = 12'h  0;
rom[33126] = 12'h  0;
rom[33127] = 12'h  0;
rom[33128] = 12'h  0;
rom[33129] = 12'h  0;
rom[33130] = 12'h  0;
rom[33131] = 12'h  0;
rom[33132] = 12'h  0;
rom[33133] = 12'h  0;
rom[33134] = 12'h  0;
rom[33135] = 12'h  0;
rom[33136] = 12'h100;
rom[33137] = 12'h100;
rom[33138] = 12'h100;
rom[33139] = 12'h200;
rom[33140] = 12'h200;
rom[33141] = 12'h300;
rom[33142] = 12'h300;
rom[33143] = 12'h400;
rom[33144] = 12'h500;
rom[33145] = 12'h700;
rom[33146] = 12'h810;
rom[33147] = 12'ha20;
rom[33148] = 12'hb40;
rom[33149] = 12'hd50;
rom[33150] = 12'he50;
rom[33151] = 12'he60;
rom[33152] = 12'he60;
rom[33153] = 12'he60;
rom[33154] = 12'he70;
rom[33155] = 12'hf92;
rom[33156] = 12'hfa3;
rom[33157] = 12'he93;
rom[33158] = 12'hb71;
rom[33159] = 12'h960;
rom[33160] = 12'h950;
rom[33161] = 12'h850;
rom[33162] = 12'h840;
rom[33163] = 12'h740;
rom[33164] = 12'h630;
rom[33165] = 12'h530;
rom[33166] = 12'h430;
rom[33167] = 12'h430;
rom[33168] = 12'h420;
rom[33169] = 12'h420;
rom[33170] = 12'h320;
rom[33171] = 12'h320;
rom[33172] = 12'h321;
rom[33173] = 12'h321;
rom[33174] = 12'h322;
rom[33175] = 12'h322;
rom[33176] = 12'h322;
rom[33177] = 12'h333;
rom[33178] = 12'h433;
rom[33179] = 12'h544;
rom[33180] = 12'h555;
rom[33181] = 12'h666;
rom[33182] = 12'h767;
rom[33183] = 12'h767;
rom[33184] = 12'h777;
rom[33185] = 12'h777;
rom[33186] = 12'h888;
rom[33187] = 12'h888;
rom[33188] = 12'h999;
rom[33189] = 12'h999;
rom[33190] = 12'h999;
rom[33191] = 12'h999;
rom[33192] = 12'h999;
rom[33193] = 12'h999;
rom[33194] = 12'haaa;
rom[33195] = 12'haaa;
rom[33196] = 12'haaa;
rom[33197] = 12'haaa;
rom[33198] = 12'hbbb;
rom[33199] = 12'hbbb;
rom[33200] = 12'h999;
rom[33201] = 12'h999;
rom[33202] = 12'h999;
rom[33203] = 12'h999;
rom[33204] = 12'h999;
rom[33205] = 12'h888;
rom[33206] = 12'h888;
rom[33207] = 12'h888;
rom[33208] = 12'h888;
rom[33209] = 12'h888;
rom[33210] = 12'h888;
rom[33211] = 12'h888;
rom[33212] = 12'h777;
rom[33213] = 12'h777;
rom[33214] = 12'h888;
rom[33215] = 12'h888;
rom[33216] = 12'h888;
rom[33217] = 12'h888;
rom[33218] = 12'h888;
rom[33219] = 12'h888;
rom[33220] = 12'h888;
rom[33221] = 12'h888;
rom[33222] = 12'h888;
rom[33223] = 12'h888;
rom[33224] = 12'h888;
rom[33225] = 12'h888;
rom[33226] = 12'h888;
rom[33227] = 12'h888;
rom[33228] = 12'h888;
rom[33229] = 12'h888;
rom[33230] = 12'h888;
rom[33231] = 12'h888;
rom[33232] = 12'h888;
rom[33233] = 12'h888;
rom[33234] = 12'h999;
rom[33235] = 12'h999;
rom[33236] = 12'h999;
rom[33237] = 12'h999;
rom[33238] = 12'h999;
rom[33239] = 12'h999;
rom[33240] = 12'h999;
rom[33241] = 12'h999;
rom[33242] = 12'h999;
rom[33243] = 12'h999;
rom[33244] = 12'h999;
rom[33245] = 12'h888;
rom[33246] = 12'h888;
rom[33247] = 12'h888;
rom[33248] = 12'h777;
rom[33249] = 12'h777;
rom[33250] = 12'h777;
rom[33251] = 12'h777;
rom[33252] = 12'h777;
rom[33253] = 12'h777;
rom[33254] = 12'h777;
rom[33255] = 12'h777;
rom[33256] = 12'h777;
rom[33257] = 12'h666;
rom[33258] = 12'h666;
rom[33259] = 12'h666;
rom[33260] = 12'h666;
rom[33261] = 12'h666;
rom[33262] = 12'h666;
rom[33263] = 12'h666;
rom[33264] = 12'h777;
rom[33265] = 12'h888;
rom[33266] = 12'h888;
rom[33267] = 12'h999;
rom[33268] = 12'h999;
rom[33269] = 12'h999;
rom[33270] = 12'h999;
rom[33271] = 12'h888;
rom[33272] = 12'h888;
rom[33273] = 12'h777;
rom[33274] = 12'h777;
rom[33275] = 12'h666;
rom[33276] = 12'h666;
rom[33277] = 12'h555;
rom[33278] = 12'h555;
rom[33279] = 12'h444;
rom[33280] = 12'h444;
rom[33281] = 12'h444;
rom[33282] = 12'h444;
rom[33283] = 12'h333;
rom[33284] = 12'h333;
rom[33285] = 12'h333;
rom[33286] = 12'h333;
rom[33287] = 12'h222;
rom[33288] = 12'h222;
rom[33289] = 12'h222;
rom[33290] = 12'h222;
rom[33291] = 12'h222;
rom[33292] = 12'h222;
rom[33293] = 12'h222;
rom[33294] = 12'h111;
rom[33295] = 12'h111;
rom[33296] = 12'h111;
rom[33297] = 12'h  0;
rom[33298] = 12'h  0;
rom[33299] = 12'h  0;
rom[33300] = 12'h  0;
rom[33301] = 12'h  0;
rom[33302] = 12'h  0;
rom[33303] = 12'h  0;
rom[33304] = 12'h  0;
rom[33305] = 12'h  0;
rom[33306] = 12'h  0;
rom[33307] = 12'h  0;
rom[33308] = 12'h  0;
rom[33309] = 12'h  0;
rom[33310] = 12'h  0;
rom[33311] = 12'h  0;
rom[33312] = 12'h  0;
rom[33313] = 12'h  0;
rom[33314] = 12'h  0;
rom[33315] = 12'h  0;
rom[33316] = 12'h  0;
rom[33317] = 12'h  0;
rom[33318] = 12'h  0;
rom[33319] = 12'h  0;
rom[33320] = 12'h  0;
rom[33321] = 12'h  0;
rom[33322] = 12'h  0;
rom[33323] = 12'h  0;
rom[33324] = 12'h  0;
rom[33325] = 12'h  0;
rom[33326] = 12'h  0;
rom[33327] = 12'h  0;
rom[33328] = 12'h  0;
rom[33329] = 12'h  0;
rom[33330] = 12'h  0;
rom[33331] = 12'h  0;
rom[33332] = 12'h  0;
rom[33333] = 12'h  0;
rom[33334] = 12'h  0;
rom[33335] = 12'h  0;
rom[33336] = 12'h  0;
rom[33337] = 12'h100;
rom[33338] = 12'h100;
rom[33339] = 12'h100;
rom[33340] = 12'h100;
rom[33341] = 12'h100;
rom[33342] = 12'h100;
rom[33343] = 12'h100;
rom[33344] = 12'h100;
rom[33345] = 12'h100;
rom[33346] = 12'h100;
rom[33347] = 12'h100;
rom[33348] = 12'h100;
rom[33349] = 12'h100;
rom[33350] = 12'h100;
rom[33351] = 12'h100;
rom[33352] = 12'h100;
rom[33353] = 12'h100;
rom[33354] = 12'h100;
rom[33355] = 12'h100;
rom[33356] = 12'h  0;
rom[33357] = 12'h  0;
rom[33358] = 12'h  0;
rom[33359] = 12'h  0;
rom[33360] = 12'h  0;
rom[33361] = 12'h  0;
rom[33362] = 12'h  0;
rom[33363] = 12'h  0;
rom[33364] = 12'h  0;
rom[33365] = 12'h  0;
rom[33366] = 12'h  0;
rom[33367] = 12'h  0;
rom[33368] = 12'h  0;
rom[33369] = 12'h  0;
rom[33370] = 12'h  0;
rom[33371] = 12'h  0;
rom[33372] = 12'h  0;
rom[33373] = 12'h  0;
rom[33374] = 12'h  0;
rom[33375] = 12'h  0;
rom[33376] = 12'h  0;
rom[33377] = 12'h  0;
rom[33378] = 12'h  0;
rom[33379] = 12'h  0;
rom[33380] = 12'h  0;
rom[33381] = 12'h  0;
rom[33382] = 12'h  0;
rom[33383] = 12'h  0;
rom[33384] = 12'h  0;
rom[33385] = 12'h  0;
rom[33386] = 12'h  0;
rom[33387] = 12'h  0;
rom[33388] = 12'h  0;
rom[33389] = 12'h  0;
rom[33390] = 12'h  0;
rom[33391] = 12'h  0;
rom[33392] = 12'h  0;
rom[33393] = 12'h  0;
rom[33394] = 12'h  0;
rom[33395] = 12'h  0;
rom[33396] = 12'h  0;
rom[33397] = 12'h  0;
rom[33398] = 12'h111;
rom[33399] = 12'h111;
rom[33400] = 12'h222;
rom[33401] = 12'h222;
rom[33402] = 12'h333;
rom[33403] = 12'h444;
rom[33404] = 12'h444;
rom[33405] = 12'h555;
rom[33406] = 12'h555;
rom[33407] = 12'h555;
rom[33408] = 12'h666;
rom[33409] = 12'h666;
rom[33410] = 12'h666;
rom[33411] = 12'h666;
rom[33412] = 12'h555;
rom[33413] = 12'h666;
rom[33414] = 12'h555;
rom[33415] = 12'h555;
rom[33416] = 12'h555;
rom[33417] = 12'h555;
rom[33418] = 12'h555;
rom[33419] = 12'h555;
rom[33420] = 12'h555;
rom[33421] = 12'h555;
rom[33422] = 12'h555;
rom[33423] = 12'h555;
rom[33424] = 12'h555;
rom[33425] = 12'h555;
rom[33426] = 12'h555;
rom[33427] = 12'h555;
rom[33428] = 12'h555;
rom[33429] = 12'h555;
rom[33430] = 12'h666;
rom[33431] = 12'h666;
rom[33432] = 12'h666;
rom[33433] = 12'h666;
rom[33434] = 12'h555;
rom[33435] = 12'h555;
rom[33436] = 12'h444;
rom[33437] = 12'h444;
rom[33438] = 12'h333;
rom[33439] = 12'h333;
rom[33440] = 12'h333;
rom[33441] = 12'h333;
rom[33442] = 12'h222;
rom[33443] = 12'h222;
rom[33444] = 12'h222;
rom[33445] = 12'h111;
rom[33446] = 12'h111;
rom[33447] = 12'h111;
rom[33448] = 12'h111;
rom[33449] = 12'h111;
rom[33450] = 12'h111;
rom[33451] = 12'h111;
rom[33452] = 12'h111;
rom[33453] = 12'h  0;
rom[33454] = 12'h  0;
rom[33455] = 12'h  0;
rom[33456] = 12'h  0;
rom[33457] = 12'h  0;
rom[33458] = 12'h  0;
rom[33459] = 12'h  0;
rom[33460] = 12'h  0;
rom[33461] = 12'h  0;
rom[33462] = 12'h  0;
rom[33463] = 12'h  0;
rom[33464] = 12'h  0;
rom[33465] = 12'h  0;
rom[33466] = 12'h  0;
rom[33467] = 12'h  0;
rom[33468] = 12'h  0;
rom[33469] = 12'h  0;
rom[33470] = 12'h  0;
rom[33471] = 12'h  0;
rom[33472] = 12'h  0;
rom[33473] = 12'h  0;
rom[33474] = 12'h  0;
rom[33475] = 12'h  0;
rom[33476] = 12'h  0;
rom[33477] = 12'h  0;
rom[33478] = 12'h  0;
rom[33479] = 12'h  0;
rom[33480] = 12'h  0;
rom[33481] = 12'h  0;
rom[33482] = 12'h  0;
rom[33483] = 12'h  0;
rom[33484] = 12'h111;
rom[33485] = 12'h111;
rom[33486] = 12'h222;
rom[33487] = 12'h222;
rom[33488] = 12'h333;
rom[33489] = 12'h333;
rom[33490] = 12'h333;
rom[33491] = 12'h333;
rom[33492] = 12'h333;
rom[33493] = 12'h333;
rom[33494] = 12'h344;
rom[33495] = 12'h444;
rom[33496] = 12'h444;
rom[33497] = 12'h555;
rom[33498] = 12'h666;
rom[33499] = 12'h777;
rom[33500] = 12'h878;
rom[33501] = 12'h988;
rom[33502] = 12'ha99;
rom[33503] = 12'hbaa;
rom[33504] = 12'hcbb;
rom[33505] = 12'hccc;
rom[33506] = 12'hddd;
rom[33507] = 12'hfee;
rom[33508] = 12'hfff;
rom[33509] = 12'hffe;
rom[33510] = 12'hbba;
rom[33511] = 12'h665;
rom[33512] = 12'h221;
rom[33513] = 12'h110;
rom[33514] = 12'h  0;
rom[33515] = 12'h100;
rom[33516] = 12'h110;
rom[33517] = 12'h100;
rom[33518] = 12'h100;
rom[33519] = 12'h  0;
rom[33520] = 12'h  0;
rom[33521] = 12'h  0;
rom[33522] = 12'h  0;
rom[33523] = 12'h  0;
rom[33524] = 12'h  0;
rom[33525] = 12'h  0;
rom[33526] = 12'h  0;
rom[33527] = 12'h  0;
rom[33528] = 12'h  0;
rom[33529] = 12'h  0;
rom[33530] = 12'h  0;
rom[33531] = 12'h  0;
rom[33532] = 12'h  0;
rom[33533] = 12'h  0;
rom[33534] = 12'h  0;
rom[33535] = 12'h  0;
rom[33536] = 12'h  0;
rom[33537] = 12'h100;
rom[33538] = 12'h100;
rom[33539] = 12'h100;
rom[33540] = 12'h200;
rom[33541] = 12'h200;
rom[33542] = 12'h300;
rom[33543] = 12'h400;
rom[33544] = 12'h500;
rom[33545] = 12'h600;
rom[33546] = 12'h810;
rom[33547] = 12'ha20;
rom[33548] = 12'hc40;
rom[33549] = 12'hd50;
rom[33550] = 12'he51;
rom[33551] = 12'hf60;
rom[33552] = 12'he60;
rom[33553] = 12'he70;
rom[33554] = 12'he81;
rom[33555] = 12'hfa3;
rom[33556] = 12'hfa3;
rom[33557] = 12'hd93;
rom[33558] = 12'hb71;
rom[33559] = 12'h950;
rom[33560] = 12'h850;
rom[33561] = 12'h850;
rom[33562] = 12'h740;
rom[33563] = 12'h630;
rom[33564] = 12'h530;
rom[33565] = 12'h530;
rom[33566] = 12'h420;
rom[33567] = 12'h420;
rom[33568] = 12'h320;
rom[33569] = 12'h320;
rom[33570] = 12'h320;
rom[33571] = 12'h310;
rom[33572] = 12'h311;
rom[33573] = 12'h321;
rom[33574] = 12'h321;
rom[33575] = 12'h322;
rom[33576] = 12'h222;
rom[33577] = 12'h222;
rom[33578] = 12'h333;
rom[33579] = 12'h444;
rom[33580] = 12'h555;
rom[33581] = 12'h656;
rom[33582] = 12'h666;
rom[33583] = 12'h666;
rom[33584] = 12'h777;
rom[33585] = 12'h777;
rom[33586] = 12'h888;
rom[33587] = 12'h888;
rom[33588] = 12'h888;
rom[33589] = 12'h999;
rom[33590] = 12'h999;
rom[33591] = 12'h999;
rom[33592] = 12'h999;
rom[33593] = 12'h999;
rom[33594] = 12'haaa;
rom[33595] = 12'haaa;
rom[33596] = 12'haaa;
rom[33597] = 12'haaa;
rom[33598] = 12'hbbb;
rom[33599] = 12'hbbb;
rom[33600] = 12'haaa;
rom[33601] = 12'h999;
rom[33602] = 12'h999;
rom[33603] = 12'h999;
rom[33604] = 12'h999;
rom[33605] = 12'h999;
rom[33606] = 12'h999;
rom[33607] = 12'h999;
rom[33608] = 12'h888;
rom[33609] = 12'h888;
rom[33610] = 12'h888;
rom[33611] = 12'h888;
rom[33612] = 12'h888;
rom[33613] = 12'h888;
rom[33614] = 12'h888;
rom[33615] = 12'h888;
rom[33616] = 12'h888;
rom[33617] = 12'h888;
rom[33618] = 12'h888;
rom[33619] = 12'h888;
rom[33620] = 12'h888;
rom[33621] = 12'h888;
rom[33622] = 12'h888;
rom[33623] = 12'h888;
rom[33624] = 12'h888;
rom[33625] = 12'h888;
rom[33626] = 12'h888;
rom[33627] = 12'h999;
rom[33628] = 12'h999;
rom[33629] = 12'h999;
rom[33630] = 12'h999;
rom[33631] = 12'h999;
rom[33632] = 12'h888;
rom[33633] = 12'h888;
rom[33634] = 12'h999;
rom[33635] = 12'h999;
rom[33636] = 12'h999;
rom[33637] = 12'h999;
rom[33638] = 12'h999;
rom[33639] = 12'h999;
rom[33640] = 12'h999;
rom[33641] = 12'h999;
rom[33642] = 12'h999;
rom[33643] = 12'h999;
rom[33644] = 12'h999;
rom[33645] = 12'h888;
rom[33646] = 12'h888;
rom[33647] = 12'h888;
rom[33648] = 12'h777;
rom[33649] = 12'h777;
rom[33650] = 12'h777;
rom[33651] = 12'h777;
rom[33652] = 12'h777;
rom[33653] = 12'h777;
rom[33654] = 12'h777;
rom[33655] = 12'h777;
rom[33656] = 12'h777;
rom[33657] = 12'h777;
rom[33658] = 12'h666;
rom[33659] = 12'h666;
rom[33660] = 12'h666;
rom[33661] = 12'h666;
rom[33662] = 12'h666;
rom[33663] = 12'h666;
rom[33664] = 12'h666;
rom[33665] = 12'h777;
rom[33666] = 12'h888;
rom[33667] = 12'h999;
rom[33668] = 12'h999;
rom[33669] = 12'h999;
rom[33670] = 12'h999;
rom[33671] = 12'h999;
rom[33672] = 12'h888;
rom[33673] = 12'h888;
rom[33674] = 12'h777;
rom[33675] = 12'h777;
rom[33676] = 12'h666;
rom[33677] = 12'h666;
rom[33678] = 12'h555;
rom[33679] = 12'h555;
rom[33680] = 12'h444;
rom[33681] = 12'h444;
rom[33682] = 12'h444;
rom[33683] = 12'h333;
rom[33684] = 12'h333;
rom[33685] = 12'h333;
rom[33686] = 12'h333;
rom[33687] = 12'h222;
rom[33688] = 12'h222;
rom[33689] = 12'h222;
rom[33690] = 12'h222;
rom[33691] = 12'h222;
rom[33692] = 12'h222;
rom[33693] = 12'h222;
rom[33694] = 12'h111;
rom[33695] = 12'h111;
rom[33696] = 12'h111;
rom[33697] = 12'h  0;
rom[33698] = 12'h  0;
rom[33699] = 12'h  0;
rom[33700] = 12'h  0;
rom[33701] = 12'h  0;
rom[33702] = 12'h  0;
rom[33703] = 12'h  0;
rom[33704] = 12'h  0;
rom[33705] = 12'h  0;
rom[33706] = 12'h  0;
rom[33707] = 12'h  0;
rom[33708] = 12'h  0;
rom[33709] = 12'h  0;
rom[33710] = 12'h  0;
rom[33711] = 12'h  0;
rom[33712] = 12'h  0;
rom[33713] = 12'h  0;
rom[33714] = 12'h  0;
rom[33715] = 12'h  0;
rom[33716] = 12'h  0;
rom[33717] = 12'h  0;
rom[33718] = 12'h  0;
rom[33719] = 12'h  0;
rom[33720] = 12'h  0;
rom[33721] = 12'h  0;
rom[33722] = 12'h  0;
rom[33723] = 12'h  0;
rom[33724] = 12'h  0;
rom[33725] = 12'h  0;
rom[33726] = 12'h  0;
rom[33727] = 12'h  0;
rom[33728] = 12'h  0;
rom[33729] = 12'h  0;
rom[33730] = 12'h  0;
rom[33731] = 12'h  0;
rom[33732] = 12'h  0;
rom[33733] = 12'h  0;
rom[33734] = 12'h  0;
rom[33735] = 12'h  0;
rom[33736] = 12'h  0;
rom[33737] = 12'h  0;
rom[33738] = 12'h  0;
rom[33739] = 12'h  0;
rom[33740] = 12'h100;
rom[33741] = 12'h100;
rom[33742] = 12'h100;
rom[33743] = 12'h100;
rom[33744] = 12'h100;
rom[33745] = 12'h100;
rom[33746] = 12'h100;
rom[33747] = 12'h100;
rom[33748] = 12'h100;
rom[33749] = 12'h100;
rom[33750] = 12'h100;
rom[33751] = 12'h100;
rom[33752] = 12'h100;
rom[33753] = 12'h100;
rom[33754] = 12'h  0;
rom[33755] = 12'h  0;
rom[33756] = 12'h  0;
rom[33757] = 12'h  0;
rom[33758] = 12'h  0;
rom[33759] = 12'h  0;
rom[33760] = 12'h  0;
rom[33761] = 12'h  0;
rom[33762] = 12'h  0;
rom[33763] = 12'h  0;
rom[33764] = 12'h  0;
rom[33765] = 12'h  0;
rom[33766] = 12'h  0;
rom[33767] = 12'h  0;
rom[33768] = 12'h  0;
rom[33769] = 12'h  0;
rom[33770] = 12'h  0;
rom[33771] = 12'h  0;
rom[33772] = 12'h  0;
rom[33773] = 12'h  0;
rom[33774] = 12'h  0;
rom[33775] = 12'h  0;
rom[33776] = 12'h  0;
rom[33777] = 12'h  0;
rom[33778] = 12'h  0;
rom[33779] = 12'h  0;
rom[33780] = 12'h  0;
rom[33781] = 12'h  0;
rom[33782] = 12'h  0;
rom[33783] = 12'h  0;
rom[33784] = 12'h  0;
rom[33785] = 12'h  0;
rom[33786] = 12'h  0;
rom[33787] = 12'h  0;
rom[33788] = 12'h  0;
rom[33789] = 12'h  0;
rom[33790] = 12'h  0;
rom[33791] = 12'h  0;
rom[33792] = 12'h  0;
rom[33793] = 12'h  0;
rom[33794] = 12'h  0;
rom[33795] = 12'h  0;
rom[33796] = 12'h  0;
rom[33797] = 12'h  0;
rom[33798] = 12'h111;
rom[33799] = 12'h111;
rom[33800] = 12'h222;
rom[33801] = 12'h333;
rom[33802] = 12'h333;
rom[33803] = 12'h444;
rom[33804] = 12'h555;
rom[33805] = 12'h555;
rom[33806] = 12'h555;
rom[33807] = 12'h555;
rom[33808] = 12'h666;
rom[33809] = 12'h666;
rom[33810] = 12'h666;
rom[33811] = 12'h555;
rom[33812] = 12'h555;
rom[33813] = 12'h555;
rom[33814] = 12'h555;
rom[33815] = 12'h555;
rom[33816] = 12'h555;
rom[33817] = 12'h555;
rom[33818] = 12'h555;
rom[33819] = 12'h555;
rom[33820] = 12'h555;
rom[33821] = 12'h555;
rom[33822] = 12'h555;
rom[33823] = 12'h555;
rom[33824] = 12'h555;
rom[33825] = 12'h555;
rom[33826] = 12'h555;
rom[33827] = 12'h555;
rom[33828] = 12'h555;
rom[33829] = 12'h555;
rom[33830] = 12'h666;
rom[33831] = 12'h666;
rom[33832] = 12'h666;
rom[33833] = 12'h666;
rom[33834] = 12'h555;
rom[33835] = 12'h555;
rom[33836] = 12'h444;
rom[33837] = 12'h444;
rom[33838] = 12'h333;
rom[33839] = 12'h333;
rom[33840] = 12'h333;
rom[33841] = 12'h333;
rom[33842] = 12'h222;
rom[33843] = 12'h222;
rom[33844] = 12'h222;
rom[33845] = 12'h111;
rom[33846] = 12'h111;
rom[33847] = 12'h111;
rom[33848] = 12'h111;
rom[33849] = 12'h111;
rom[33850] = 12'h111;
rom[33851] = 12'h111;
rom[33852] = 12'h111;
rom[33853] = 12'h  0;
rom[33854] = 12'h  0;
rom[33855] = 12'h  0;
rom[33856] = 12'h  0;
rom[33857] = 12'h  0;
rom[33858] = 12'h  0;
rom[33859] = 12'h  0;
rom[33860] = 12'h  0;
rom[33861] = 12'h  0;
rom[33862] = 12'h  0;
rom[33863] = 12'h  0;
rom[33864] = 12'h  0;
rom[33865] = 12'h  0;
rom[33866] = 12'h  0;
rom[33867] = 12'h  0;
rom[33868] = 12'h  0;
rom[33869] = 12'h  0;
rom[33870] = 12'h  0;
rom[33871] = 12'h  0;
rom[33872] = 12'h  0;
rom[33873] = 12'h  0;
rom[33874] = 12'h  0;
rom[33875] = 12'h  0;
rom[33876] = 12'h  0;
rom[33877] = 12'h  0;
rom[33878] = 12'h  0;
rom[33879] = 12'h  0;
rom[33880] = 12'h  0;
rom[33881] = 12'h  0;
rom[33882] = 12'h  0;
rom[33883] = 12'h  0;
rom[33884] = 12'h111;
rom[33885] = 12'h111;
rom[33886] = 12'h222;
rom[33887] = 12'h222;
rom[33888] = 12'h333;
rom[33889] = 12'h333;
rom[33890] = 12'h333;
rom[33891] = 12'h333;
rom[33892] = 12'h333;
rom[33893] = 12'h333;
rom[33894] = 12'h444;
rom[33895] = 12'h444;
rom[33896] = 12'h555;
rom[33897] = 12'h566;
rom[33898] = 12'h777;
rom[33899] = 12'h877;
rom[33900] = 12'h888;
rom[33901] = 12'h999;
rom[33902] = 12'haaa;
rom[33903] = 12'hbbb;
rom[33904] = 12'hccb;
rom[33905] = 12'hddc;
rom[33906] = 12'hfee;
rom[33907] = 12'hfff;
rom[33908] = 12'hffe;
rom[33909] = 12'hcba;
rom[33910] = 12'h765;
rom[33911] = 12'h322;
rom[33912] = 12'h110;
rom[33913] = 12'h110;
rom[33914] = 12'h100;
rom[33915] = 12'h100;
rom[33916] = 12'h  0;
rom[33917] = 12'h  0;
rom[33918] = 12'h  0;
rom[33919] = 12'h  0;
rom[33920] = 12'h  0;
rom[33921] = 12'h  0;
rom[33922] = 12'h  0;
rom[33923] = 12'h  0;
rom[33924] = 12'h  0;
rom[33925] = 12'h  0;
rom[33926] = 12'h  0;
rom[33927] = 12'h  0;
rom[33928] = 12'h  0;
rom[33929] = 12'h  0;
rom[33930] = 12'h  0;
rom[33931] = 12'h  0;
rom[33932] = 12'h  0;
rom[33933] = 12'h  0;
rom[33934] = 12'h  0;
rom[33935] = 12'h  0;
rom[33936] = 12'h  0;
rom[33937] = 12'h100;
rom[33938] = 12'h100;
rom[33939] = 12'h100;
rom[33940] = 12'h200;
rom[33941] = 12'h200;
rom[33942] = 12'h300;
rom[33943] = 12'h400;
rom[33944] = 12'h500;
rom[33945] = 12'h600;
rom[33946] = 12'h810;
rom[33947] = 12'ha20;
rom[33948] = 12'hc40;
rom[33949] = 12'he51;
rom[33950] = 12'hf51;
rom[33951] = 12'hf60;
rom[33952] = 12'he60;
rom[33953] = 12'he70;
rom[33954] = 12'hf81;
rom[33955] = 12'hfa3;
rom[33956] = 12'hfb4;
rom[33957] = 12'hd92;
rom[33958] = 12'ha70;
rom[33959] = 12'h950;
rom[33960] = 12'h850;
rom[33961] = 12'h840;
rom[33962] = 12'h740;
rom[33963] = 12'h630;
rom[33964] = 12'h530;
rom[33965] = 12'h420;
rom[33966] = 12'h420;
rom[33967] = 12'h320;
rom[33968] = 12'h310;
rom[33969] = 12'h310;
rom[33970] = 12'h310;
rom[33971] = 12'h210;
rom[33972] = 12'h210;
rom[33973] = 12'h211;
rom[33974] = 12'h211;
rom[33975] = 12'h222;
rom[33976] = 12'h222;
rom[33977] = 12'h222;
rom[33978] = 12'h323;
rom[33979] = 12'h434;
rom[33980] = 12'h545;
rom[33981] = 12'h656;
rom[33982] = 12'h666;
rom[33983] = 12'h667;
rom[33984] = 12'h777;
rom[33985] = 12'h777;
rom[33986] = 12'h777;
rom[33987] = 12'h888;
rom[33988] = 12'h888;
rom[33989] = 12'h999;
rom[33990] = 12'h999;
rom[33991] = 12'h999;
rom[33992] = 12'h999;
rom[33993] = 12'haaa;
rom[33994] = 12'haaa;
rom[33995] = 12'haaa;
rom[33996] = 12'haaa;
rom[33997] = 12'haaa;
rom[33998] = 12'hbbb;
rom[33999] = 12'hbbb;
rom[34000] = 12'haaa;
rom[34001] = 12'haaa;
rom[34002] = 12'h999;
rom[34003] = 12'h999;
rom[34004] = 12'h999;
rom[34005] = 12'h999;
rom[34006] = 12'h999;
rom[34007] = 12'h999;
rom[34008] = 12'h999;
rom[34009] = 12'h999;
rom[34010] = 12'h999;
rom[34011] = 12'h888;
rom[34012] = 12'h888;
rom[34013] = 12'h999;
rom[34014] = 12'h999;
rom[34015] = 12'h999;
rom[34016] = 12'h888;
rom[34017] = 12'h888;
rom[34018] = 12'h888;
rom[34019] = 12'h888;
rom[34020] = 12'h888;
rom[34021] = 12'h888;
rom[34022] = 12'h888;
rom[34023] = 12'h888;
rom[34024] = 12'h888;
rom[34025] = 12'h888;
rom[34026] = 12'h888;
rom[34027] = 12'h888;
rom[34028] = 12'h999;
rom[34029] = 12'h999;
rom[34030] = 12'h999;
rom[34031] = 12'h999;
rom[34032] = 12'h999;
rom[34033] = 12'h999;
rom[34034] = 12'h999;
rom[34035] = 12'h999;
rom[34036] = 12'h999;
rom[34037] = 12'h999;
rom[34038] = 12'h999;
rom[34039] = 12'h999;
rom[34040] = 12'h999;
rom[34041] = 12'h999;
rom[34042] = 12'h999;
rom[34043] = 12'h999;
rom[34044] = 12'h999;
rom[34045] = 12'h999;
rom[34046] = 12'h888;
rom[34047] = 12'h888;
rom[34048] = 12'h888;
rom[34049] = 12'h777;
rom[34050] = 12'h777;
rom[34051] = 12'h777;
rom[34052] = 12'h777;
rom[34053] = 12'h777;
rom[34054] = 12'h777;
rom[34055] = 12'h777;
rom[34056] = 12'h777;
rom[34057] = 12'h777;
rom[34058] = 12'h666;
rom[34059] = 12'h666;
rom[34060] = 12'h666;
rom[34061] = 12'h666;
rom[34062] = 12'h666;
rom[34063] = 12'h666;
rom[34064] = 12'h666;
rom[34065] = 12'h777;
rom[34066] = 12'h777;
rom[34067] = 12'h888;
rom[34068] = 12'h999;
rom[34069] = 12'h999;
rom[34070] = 12'haaa;
rom[34071] = 12'haaa;
rom[34072] = 12'h999;
rom[34073] = 12'h888;
rom[34074] = 12'h777;
rom[34075] = 12'h777;
rom[34076] = 12'h777;
rom[34077] = 12'h666;
rom[34078] = 12'h555;
rom[34079] = 12'h555;
rom[34080] = 12'h555;
rom[34081] = 12'h444;
rom[34082] = 12'h444;
rom[34083] = 12'h444;
rom[34084] = 12'h333;
rom[34085] = 12'h333;
rom[34086] = 12'h333;
rom[34087] = 12'h333;
rom[34088] = 12'h222;
rom[34089] = 12'h222;
rom[34090] = 12'h222;
rom[34091] = 12'h222;
rom[34092] = 12'h222;
rom[34093] = 12'h222;
rom[34094] = 12'h111;
rom[34095] = 12'h111;
rom[34096] = 12'h111;
rom[34097] = 12'h111;
rom[34098] = 12'h  0;
rom[34099] = 12'h  0;
rom[34100] = 12'h  0;
rom[34101] = 12'h  0;
rom[34102] = 12'h  0;
rom[34103] = 12'h  0;
rom[34104] = 12'h  0;
rom[34105] = 12'h  0;
rom[34106] = 12'h  0;
rom[34107] = 12'h  0;
rom[34108] = 12'h  0;
rom[34109] = 12'h  0;
rom[34110] = 12'h  0;
rom[34111] = 12'h  0;
rom[34112] = 12'h  0;
rom[34113] = 12'h  0;
rom[34114] = 12'h  0;
rom[34115] = 12'h  0;
rom[34116] = 12'h  0;
rom[34117] = 12'h  0;
rom[34118] = 12'h  0;
rom[34119] = 12'h  0;
rom[34120] = 12'h  0;
rom[34121] = 12'h  0;
rom[34122] = 12'h  0;
rom[34123] = 12'h  0;
rom[34124] = 12'h  0;
rom[34125] = 12'h  0;
rom[34126] = 12'h  0;
rom[34127] = 12'h  0;
rom[34128] = 12'h  0;
rom[34129] = 12'h  0;
rom[34130] = 12'h  0;
rom[34131] = 12'h  0;
rom[34132] = 12'h  0;
rom[34133] = 12'h  0;
rom[34134] = 12'h  0;
rom[34135] = 12'h  0;
rom[34136] = 12'h  0;
rom[34137] = 12'h  0;
rom[34138] = 12'h  0;
rom[34139] = 12'h  0;
rom[34140] = 12'h  0;
rom[34141] = 12'h  0;
rom[34142] = 12'h  0;
rom[34143] = 12'h100;
rom[34144] = 12'h100;
rom[34145] = 12'h100;
rom[34146] = 12'h100;
rom[34147] = 12'h100;
rom[34148] = 12'h100;
rom[34149] = 12'h100;
rom[34150] = 12'h  0;
rom[34151] = 12'h  0;
rom[34152] = 12'h  0;
rom[34153] = 12'h  0;
rom[34154] = 12'h  0;
rom[34155] = 12'h  0;
rom[34156] = 12'h  0;
rom[34157] = 12'h  0;
rom[34158] = 12'h  0;
rom[34159] = 12'h  0;
rom[34160] = 12'h  0;
rom[34161] = 12'h  0;
rom[34162] = 12'h  0;
rom[34163] = 12'h  0;
rom[34164] = 12'h  0;
rom[34165] = 12'h  0;
rom[34166] = 12'h  0;
rom[34167] = 12'h  0;
rom[34168] = 12'h  0;
rom[34169] = 12'h  0;
rom[34170] = 12'h  0;
rom[34171] = 12'h  0;
rom[34172] = 12'h  0;
rom[34173] = 12'h  0;
rom[34174] = 12'h  0;
rom[34175] = 12'h  0;
rom[34176] = 12'h  0;
rom[34177] = 12'h  0;
rom[34178] = 12'h  0;
rom[34179] = 12'h  0;
rom[34180] = 12'h  0;
rom[34181] = 12'h  0;
rom[34182] = 12'h  0;
rom[34183] = 12'h  0;
rom[34184] = 12'h  0;
rom[34185] = 12'h  0;
rom[34186] = 12'h  0;
rom[34187] = 12'h  0;
rom[34188] = 12'h  0;
rom[34189] = 12'h  0;
rom[34190] = 12'h  0;
rom[34191] = 12'h  0;
rom[34192] = 12'h  0;
rom[34193] = 12'h  0;
rom[34194] = 12'h  0;
rom[34195] = 12'h  0;
rom[34196] = 12'h  0;
rom[34197] = 12'h  0;
rom[34198] = 12'h111;
rom[34199] = 12'h111;
rom[34200] = 12'h222;
rom[34201] = 12'h333;
rom[34202] = 12'h444;
rom[34203] = 12'h444;
rom[34204] = 12'h555;
rom[34205] = 12'h555;
rom[34206] = 12'h555;
rom[34207] = 12'h555;
rom[34208] = 12'h666;
rom[34209] = 12'h666;
rom[34210] = 12'h666;
rom[34211] = 12'h555;
rom[34212] = 12'h555;
rom[34213] = 12'h555;
rom[34214] = 12'h555;
rom[34215] = 12'h555;
rom[34216] = 12'h555;
rom[34217] = 12'h555;
rom[34218] = 12'h555;
rom[34219] = 12'h555;
rom[34220] = 12'h555;
rom[34221] = 12'h555;
rom[34222] = 12'h555;
rom[34223] = 12'h555;
rom[34224] = 12'h555;
rom[34225] = 12'h444;
rom[34226] = 12'h444;
rom[34227] = 12'h444;
rom[34228] = 12'h555;
rom[34229] = 12'h555;
rom[34230] = 12'h555;
rom[34231] = 12'h666;
rom[34232] = 12'h666;
rom[34233] = 12'h555;
rom[34234] = 12'h555;
rom[34235] = 12'h444;
rom[34236] = 12'h444;
rom[34237] = 12'h444;
rom[34238] = 12'h333;
rom[34239] = 12'h333;
rom[34240] = 12'h333;
rom[34241] = 12'h333;
rom[34242] = 12'h222;
rom[34243] = 12'h222;
rom[34244] = 12'h222;
rom[34245] = 12'h111;
rom[34246] = 12'h111;
rom[34247] = 12'h111;
rom[34248] = 12'h111;
rom[34249] = 12'h111;
rom[34250] = 12'h111;
rom[34251] = 12'h111;
rom[34252] = 12'h111;
rom[34253] = 12'h  0;
rom[34254] = 12'h  0;
rom[34255] = 12'h  0;
rom[34256] = 12'h  0;
rom[34257] = 12'h  0;
rom[34258] = 12'h  0;
rom[34259] = 12'h  0;
rom[34260] = 12'h  0;
rom[34261] = 12'h  0;
rom[34262] = 12'h  0;
rom[34263] = 12'h  0;
rom[34264] = 12'h  0;
rom[34265] = 12'h  0;
rom[34266] = 12'h  0;
rom[34267] = 12'h  0;
rom[34268] = 12'h  0;
rom[34269] = 12'h  0;
rom[34270] = 12'h  0;
rom[34271] = 12'h  0;
rom[34272] = 12'h  0;
rom[34273] = 12'h  0;
rom[34274] = 12'h  0;
rom[34275] = 12'h  0;
rom[34276] = 12'h  0;
rom[34277] = 12'h  0;
rom[34278] = 12'h  0;
rom[34279] = 12'h  0;
rom[34280] = 12'h  0;
rom[34281] = 12'h  0;
rom[34282] = 12'h  0;
rom[34283] = 12'h  0;
rom[34284] = 12'h111;
rom[34285] = 12'h111;
rom[34286] = 12'h222;
rom[34287] = 12'h322;
rom[34288] = 12'h333;
rom[34289] = 12'h333;
rom[34290] = 12'h333;
rom[34291] = 12'h333;
rom[34292] = 12'h333;
rom[34293] = 12'h333;
rom[34294] = 12'h444;
rom[34295] = 12'h455;
rom[34296] = 12'h555;
rom[34297] = 12'h666;
rom[34298] = 12'h777;
rom[34299] = 12'h888;
rom[34300] = 12'h999;
rom[34301] = 12'haa9;
rom[34302] = 12'hbbb;
rom[34303] = 12'hccb;
rom[34304] = 12'hdcc;
rom[34305] = 12'hfee;
rom[34306] = 12'hfff;
rom[34307] = 12'hffe;
rom[34308] = 12'hcba;
rom[34309] = 12'h766;
rom[34310] = 12'h432;
rom[34311] = 12'h221;
rom[34312] = 12'h110;
rom[34313] = 12'h110;
rom[34314] = 12'h110;
rom[34315] = 12'h  0;
rom[34316] = 12'h  0;
rom[34317] = 12'h  0;
rom[34318] = 12'h  0;
rom[34319] = 12'h  0;
rom[34320] = 12'h  0;
rom[34321] = 12'h  0;
rom[34322] = 12'h  0;
rom[34323] = 12'h  0;
rom[34324] = 12'h  0;
rom[34325] = 12'h  0;
rom[34326] = 12'h  0;
rom[34327] = 12'h  0;
rom[34328] = 12'h  0;
rom[34329] = 12'h  0;
rom[34330] = 12'h  0;
rom[34331] = 12'h  0;
rom[34332] = 12'h  0;
rom[34333] = 12'h  0;
rom[34334] = 12'h  0;
rom[34335] = 12'h  0;
rom[34336] = 12'h  0;
rom[34337] = 12'h100;
rom[34338] = 12'h100;
rom[34339] = 12'h100;
rom[34340] = 12'h200;
rom[34341] = 12'h200;
rom[34342] = 12'h300;
rom[34343] = 12'h300;
rom[34344] = 12'h500;
rom[34345] = 12'h610;
rom[34346] = 12'h820;
rom[34347] = 12'ha30;
rom[34348] = 12'hc40;
rom[34349] = 12'he51;
rom[34350] = 12'hf51;
rom[34351] = 12'hf60;
rom[34352] = 12'he60;
rom[34353] = 12'he70;
rom[34354] = 12'hf92;
rom[34355] = 12'hfb4;
rom[34356] = 12'hfa4;
rom[34357] = 12'hc82;
rom[34358] = 12'ha60;
rom[34359] = 12'h950;
rom[34360] = 12'h850;
rom[34361] = 12'h740;
rom[34362] = 12'h630;
rom[34363] = 12'h630;
rom[34364] = 12'h520;
rom[34365] = 12'h420;
rom[34366] = 12'h320;
rom[34367] = 12'h310;
rom[34368] = 12'h310;
rom[34369] = 12'h210;
rom[34370] = 12'h210;
rom[34371] = 12'h210;
rom[34372] = 12'h210;
rom[34373] = 12'h211;
rom[34374] = 12'h211;
rom[34375] = 12'h211;
rom[34376] = 12'h222;
rom[34377] = 12'h223;
rom[34378] = 12'h323;
rom[34379] = 12'h334;
rom[34380] = 12'h445;
rom[34381] = 12'h556;
rom[34382] = 12'h666;
rom[34383] = 12'h667;
rom[34384] = 12'h777;
rom[34385] = 12'h777;
rom[34386] = 12'h777;
rom[34387] = 12'h888;
rom[34388] = 12'h888;
rom[34389] = 12'h999;
rom[34390] = 12'h999;
rom[34391] = 12'h999;
rom[34392] = 12'h999;
rom[34393] = 12'haaa;
rom[34394] = 12'haaa;
rom[34395] = 12'haaa;
rom[34396] = 12'haaa;
rom[34397] = 12'haaa;
rom[34398] = 12'haaa;
rom[34399] = 12'hbbb;
rom[34400] = 12'h999;
rom[34401] = 12'h999;
rom[34402] = 12'h999;
rom[34403] = 12'h999;
rom[34404] = 12'h999;
rom[34405] = 12'h999;
rom[34406] = 12'h999;
rom[34407] = 12'h999;
rom[34408] = 12'h999;
rom[34409] = 12'h999;
rom[34410] = 12'h999;
rom[34411] = 12'h999;
rom[34412] = 12'h999;
rom[34413] = 12'h999;
rom[34414] = 12'h999;
rom[34415] = 12'h999;
rom[34416] = 12'h999;
rom[34417] = 12'h999;
rom[34418] = 12'h999;
rom[34419] = 12'h999;
rom[34420] = 12'h999;
rom[34421] = 12'h999;
rom[34422] = 12'h888;
rom[34423] = 12'h888;
rom[34424] = 12'h888;
rom[34425] = 12'h888;
rom[34426] = 12'h999;
rom[34427] = 12'h999;
rom[34428] = 12'h999;
rom[34429] = 12'h999;
rom[34430] = 12'h999;
rom[34431] = 12'h999;
rom[34432] = 12'h999;
rom[34433] = 12'h999;
rom[34434] = 12'h999;
rom[34435] = 12'h999;
rom[34436] = 12'h999;
rom[34437] = 12'h999;
rom[34438] = 12'h999;
rom[34439] = 12'h999;
rom[34440] = 12'haaa;
rom[34441] = 12'haaa;
rom[34442] = 12'h999;
rom[34443] = 12'h999;
rom[34444] = 12'h999;
rom[34445] = 12'h999;
rom[34446] = 12'h999;
rom[34447] = 12'h888;
rom[34448] = 12'h888;
rom[34449] = 12'h888;
rom[34450] = 12'h777;
rom[34451] = 12'h777;
rom[34452] = 12'h777;
rom[34453] = 12'h777;
rom[34454] = 12'h777;
rom[34455] = 12'h777;
rom[34456] = 12'h777;
rom[34457] = 12'h777;
rom[34458] = 12'h666;
rom[34459] = 12'h666;
rom[34460] = 12'h666;
rom[34461] = 12'h666;
rom[34462] = 12'h666;
rom[34463] = 12'h666;
rom[34464] = 12'h777;
rom[34465] = 12'h777;
rom[34466] = 12'h777;
rom[34467] = 12'h777;
rom[34468] = 12'h888;
rom[34469] = 12'h999;
rom[34470] = 12'h999;
rom[34471] = 12'haaa;
rom[34472] = 12'h999;
rom[34473] = 12'h999;
rom[34474] = 12'h888;
rom[34475] = 12'h888;
rom[34476] = 12'h777;
rom[34477] = 12'h777;
rom[34478] = 12'h666;
rom[34479] = 12'h555;
rom[34480] = 12'h555;
rom[34481] = 12'h555;
rom[34482] = 12'h555;
rom[34483] = 12'h444;
rom[34484] = 12'h444;
rom[34485] = 12'h444;
rom[34486] = 12'h333;
rom[34487] = 12'h333;
rom[34488] = 12'h333;
rom[34489] = 12'h333;
rom[34490] = 12'h222;
rom[34491] = 12'h222;
rom[34492] = 12'h222;
rom[34493] = 12'h222;
rom[34494] = 12'h222;
rom[34495] = 12'h111;
rom[34496] = 12'h111;
rom[34497] = 12'h111;
rom[34498] = 12'h  0;
rom[34499] = 12'h  0;
rom[34500] = 12'h  0;
rom[34501] = 12'h  0;
rom[34502] = 12'h  0;
rom[34503] = 12'h  0;
rom[34504] = 12'h  0;
rom[34505] = 12'h  0;
rom[34506] = 12'h  0;
rom[34507] = 12'h  0;
rom[34508] = 12'h  0;
rom[34509] = 12'h  0;
rom[34510] = 12'h  0;
rom[34511] = 12'h  0;
rom[34512] = 12'h  0;
rom[34513] = 12'h  0;
rom[34514] = 12'h  0;
rom[34515] = 12'h  0;
rom[34516] = 12'h  0;
rom[34517] = 12'h  0;
rom[34518] = 12'h  0;
rom[34519] = 12'h  0;
rom[34520] = 12'h  0;
rom[34521] = 12'h  0;
rom[34522] = 12'h  0;
rom[34523] = 12'h  0;
rom[34524] = 12'h  0;
rom[34525] = 12'h  0;
rom[34526] = 12'h  0;
rom[34527] = 12'h  0;
rom[34528] = 12'h  0;
rom[34529] = 12'h  0;
rom[34530] = 12'h  0;
rom[34531] = 12'h  0;
rom[34532] = 12'h  0;
rom[34533] = 12'h  0;
rom[34534] = 12'h  0;
rom[34535] = 12'h  0;
rom[34536] = 12'h  0;
rom[34537] = 12'h  0;
rom[34538] = 12'h  0;
rom[34539] = 12'h  0;
rom[34540] = 12'h  0;
rom[34541] = 12'h  0;
rom[34542] = 12'h  0;
rom[34543] = 12'h  0;
rom[34544] = 12'h  0;
rom[34545] = 12'h  0;
rom[34546] = 12'h  0;
rom[34547] = 12'h  0;
rom[34548] = 12'h  0;
rom[34549] = 12'h  0;
rom[34550] = 12'h  0;
rom[34551] = 12'h  0;
rom[34552] = 12'h  0;
rom[34553] = 12'h  0;
rom[34554] = 12'h  0;
rom[34555] = 12'h  0;
rom[34556] = 12'h  0;
rom[34557] = 12'h  0;
rom[34558] = 12'h  0;
rom[34559] = 12'h  0;
rom[34560] = 12'h  0;
rom[34561] = 12'h  0;
rom[34562] = 12'h  0;
rom[34563] = 12'h  0;
rom[34564] = 12'h  0;
rom[34565] = 12'h  0;
rom[34566] = 12'h  0;
rom[34567] = 12'h  0;
rom[34568] = 12'h  0;
rom[34569] = 12'h  0;
rom[34570] = 12'h  0;
rom[34571] = 12'h  0;
rom[34572] = 12'h  0;
rom[34573] = 12'h  0;
rom[34574] = 12'h  0;
rom[34575] = 12'h  0;
rom[34576] = 12'h  0;
rom[34577] = 12'h  0;
rom[34578] = 12'h  0;
rom[34579] = 12'h  0;
rom[34580] = 12'h  0;
rom[34581] = 12'h  0;
rom[34582] = 12'h  0;
rom[34583] = 12'h  0;
rom[34584] = 12'h  0;
rom[34585] = 12'h  0;
rom[34586] = 12'h  0;
rom[34587] = 12'h  0;
rom[34588] = 12'h  0;
rom[34589] = 12'h  0;
rom[34590] = 12'h  0;
rom[34591] = 12'h  0;
rom[34592] = 12'h  0;
rom[34593] = 12'h  0;
rom[34594] = 12'h  0;
rom[34595] = 12'h  0;
rom[34596] = 12'h  0;
rom[34597] = 12'h  0;
rom[34598] = 12'h111;
rom[34599] = 12'h111;
rom[34600] = 12'h222;
rom[34601] = 12'h333;
rom[34602] = 12'h444;
rom[34603] = 12'h444;
rom[34604] = 12'h555;
rom[34605] = 12'h555;
rom[34606] = 12'h555;
rom[34607] = 12'h555;
rom[34608] = 12'h666;
rom[34609] = 12'h666;
rom[34610] = 12'h666;
rom[34611] = 12'h555;
rom[34612] = 12'h555;
rom[34613] = 12'h555;
rom[34614] = 12'h555;
rom[34615] = 12'h555;
rom[34616] = 12'h555;
rom[34617] = 12'h555;
rom[34618] = 12'h555;
rom[34619] = 12'h555;
rom[34620] = 12'h555;
rom[34621] = 12'h555;
rom[34622] = 12'h555;
rom[34623] = 12'h444;
rom[34624] = 12'h555;
rom[34625] = 12'h444;
rom[34626] = 12'h444;
rom[34627] = 12'h444;
rom[34628] = 12'h555;
rom[34629] = 12'h555;
rom[34630] = 12'h555;
rom[34631] = 12'h666;
rom[34632] = 12'h666;
rom[34633] = 12'h555;
rom[34634] = 12'h555;
rom[34635] = 12'h444;
rom[34636] = 12'h444;
rom[34637] = 12'h444;
rom[34638] = 12'h333;
rom[34639] = 12'h333;
rom[34640] = 12'h333;
rom[34641] = 12'h333;
rom[34642] = 12'h222;
rom[34643] = 12'h222;
rom[34644] = 12'h222;
rom[34645] = 12'h111;
rom[34646] = 12'h111;
rom[34647] = 12'h111;
rom[34648] = 12'h111;
rom[34649] = 12'h111;
rom[34650] = 12'h111;
rom[34651] = 12'h111;
rom[34652] = 12'h111;
rom[34653] = 12'h  0;
rom[34654] = 12'h  0;
rom[34655] = 12'h  0;
rom[34656] = 12'h  0;
rom[34657] = 12'h  0;
rom[34658] = 12'h  0;
rom[34659] = 12'h  0;
rom[34660] = 12'h  0;
rom[34661] = 12'h  0;
rom[34662] = 12'h  0;
rom[34663] = 12'h  0;
rom[34664] = 12'h  0;
rom[34665] = 12'h  0;
rom[34666] = 12'h  0;
rom[34667] = 12'h  0;
rom[34668] = 12'h  0;
rom[34669] = 12'h  0;
rom[34670] = 12'h  0;
rom[34671] = 12'h  0;
rom[34672] = 12'h  0;
rom[34673] = 12'h  0;
rom[34674] = 12'h  0;
rom[34675] = 12'h  0;
rom[34676] = 12'h  0;
rom[34677] = 12'h  0;
rom[34678] = 12'h  0;
rom[34679] = 12'h  0;
rom[34680] = 12'h  0;
rom[34681] = 12'h  0;
rom[34682] = 12'h  0;
rom[34683] = 12'h111;
rom[34684] = 12'h111;
rom[34685] = 12'h222;
rom[34686] = 12'h222;
rom[34687] = 12'h333;
rom[34688] = 12'h433;
rom[34689] = 12'h333;
rom[34690] = 12'h333;
rom[34691] = 12'h333;
rom[34692] = 12'h333;
rom[34693] = 12'h444;
rom[34694] = 12'h454;
rom[34695] = 12'h555;
rom[34696] = 12'h666;
rom[34697] = 12'h777;
rom[34698] = 12'h888;
rom[34699] = 12'h999;
rom[34700] = 12'h999;
rom[34701] = 12'haaa;
rom[34702] = 12'hbbb;
rom[34703] = 12'hdcc;
rom[34704] = 12'hedd;
rom[34705] = 12'hffe;
rom[34706] = 12'hffe;
rom[34707] = 12'hdcb;
rom[34708] = 12'h876;
rom[34709] = 12'h432;
rom[34710] = 12'h321;
rom[34711] = 12'h210;
rom[34712] = 12'h210;
rom[34713] = 12'h110;
rom[34714] = 12'h100;
rom[34715] = 12'h  0;
rom[34716] = 12'h  0;
rom[34717] = 12'h  0;
rom[34718] = 12'h  0;
rom[34719] = 12'h  0;
rom[34720] = 12'h  0;
rom[34721] = 12'h  0;
rom[34722] = 12'h  0;
rom[34723] = 12'h  0;
rom[34724] = 12'h  0;
rom[34725] = 12'h  0;
rom[34726] = 12'h  0;
rom[34727] = 12'h  0;
rom[34728] = 12'h  0;
rom[34729] = 12'h  0;
rom[34730] = 12'h  0;
rom[34731] = 12'h  0;
rom[34732] = 12'h  0;
rom[34733] = 12'h  0;
rom[34734] = 12'h  0;
rom[34735] = 12'h  0;
rom[34736] = 12'h  0;
rom[34737] = 12'h100;
rom[34738] = 12'h100;
rom[34739] = 12'h100;
rom[34740] = 12'h200;
rom[34741] = 12'h200;
rom[34742] = 12'h300;
rom[34743] = 12'h400;
rom[34744] = 12'h500;
rom[34745] = 12'h710;
rom[34746] = 12'h820;
rom[34747] = 12'hb30;
rom[34748] = 12'hd41;
rom[34749] = 12'hf51;
rom[34750] = 12'hf61;
rom[34751] = 12'hf60;
rom[34752] = 12'he70;
rom[34753] = 12'he81;
rom[34754] = 12'hfa3;
rom[34755] = 12'hfb4;
rom[34756] = 12'hea3;
rom[34757] = 12'hb71;
rom[34758] = 12'h950;
rom[34759] = 12'h950;
rom[34760] = 12'h840;
rom[34761] = 12'h730;
rom[34762] = 12'h630;
rom[34763] = 12'h520;
rom[34764] = 12'h520;
rom[34765] = 12'h420;
rom[34766] = 12'h320;
rom[34767] = 12'h310;
rom[34768] = 12'h310;
rom[34769] = 12'h210;
rom[34770] = 12'h210;
rom[34771] = 12'h210;
rom[34772] = 12'h210;
rom[34773] = 12'h211;
rom[34774] = 12'h211;
rom[34775] = 12'h211;
rom[34776] = 12'h223;
rom[34777] = 12'h323;
rom[34778] = 12'h333;
rom[34779] = 12'h334;
rom[34780] = 12'h445;
rom[34781] = 12'h555;
rom[34782] = 12'h666;
rom[34783] = 12'h667;
rom[34784] = 12'h777;
rom[34785] = 12'h777;
rom[34786] = 12'h777;
rom[34787] = 12'h888;
rom[34788] = 12'h888;
rom[34789] = 12'h999;
rom[34790] = 12'h999;
rom[34791] = 12'h999;
rom[34792] = 12'haaa;
rom[34793] = 12'haaa;
rom[34794] = 12'haaa;
rom[34795] = 12'haaa;
rom[34796] = 12'haaa;
rom[34797] = 12'haaa;
rom[34798] = 12'haaa;
rom[34799] = 12'hbbb;
rom[34800] = 12'h888;
rom[34801] = 12'h888;
rom[34802] = 12'h888;
rom[34803] = 12'h888;
rom[34804] = 12'h888;
rom[34805] = 12'h888;
rom[34806] = 12'h888;
rom[34807] = 12'h888;
rom[34808] = 12'h888;
rom[34809] = 12'h999;
rom[34810] = 12'h999;
rom[34811] = 12'h999;
rom[34812] = 12'h999;
rom[34813] = 12'h999;
rom[34814] = 12'h999;
rom[34815] = 12'h999;
rom[34816] = 12'h999;
rom[34817] = 12'h999;
rom[34818] = 12'h999;
rom[34819] = 12'h999;
rom[34820] = 12'h999;
rom[34821] = 12'h999;
rom[34822] = 12'h999;
rom[34823] = 12'h999;
rom[34824] = 12'h999;
rom[34825] = 12'h999;
rom[34826] = 12'h999;
rom[34827] = 12'h999;
rom[34828] = 12'h999;
rom[34829] = 12'h999;
rom[34830] = 12'h999;
rom[34831] = 12'h999;
rom[34832] = 12'h999;
rom[34833] = 12'h999;
rom[34834] = 12'h999;
rom[34835] = 12'h999;
rom[34836] = 12'h999;
rom[34837] = 12'h999;
rom[34838] = 12'h999;
rom[34839] = 12'h999;
rom[34840] = 12'haaa;
rom[34841] = 12'haaa;
rom[34842] = 12'h999;
rom[34843] = 12'h999;
rom[34844] = 12'h999;
rom[34845] = 12'h999;
rom[34846] = 12'h999;
rom[34847] = 12'h999;
rom[34848] = 12'h888;
rom[34849] = 12'h888;
rom[34850] = 12'h888;
rom[34851] = 12'h777;
rom[34852] = 12'h777;
rom[34853] = 12'h777;
rom[34854] = 12'h777;
rom[34855] = 12'h777;
rom[34856] = 12'h777;
rom[34857] = 12'h777;
rom[34858] = 12'h777;
rom[34859] = 12'h777;
rom[34860] = 12'h777;
rom[34861] = 12'h666;
rom[34862] = 12'h666;
rom[34863] = 12'h666;
rom[34864] = 12'h777;
rom[34865] = 12'h777;
rom[34866] = 12'h666;
rom[34867] = 12'h666;
rom[34868] = 12'h777;
rom[34869] = 12'h888;
rom[34870] = 12'h999;
rom[34871] = 12'h999;
rom[34872] = 12'haaa;
rom[34873] = 12'h999;
rom[34874] = 12'h999;
rom[34875] = 12'h888;
rom[34876] = 12'h888;
rom[34877] = 12'h888;
rom[34878] = 12'h777;
rom[34879] = 12'h666;
rom[34880] = 12'h666;
rom[34881] = 12'h555;
rom[34882] = 12'h555;
rom[34883] = 12'h444;
rom[34884] = 12'h444;
rom[34885] = 12'h444;
rom[34886] = 12'h444;
rom[34887] = 12'h333;
rom[34888] = 12'h333;
rom[34889] = 12'h333;
rom[34890] = 12'h222;
rom[34891] = 12'h222;
rom[34892] = 12'h222;
rom[34893] = 12'h222;
rom[34894] = 12'h222;
rom[34895] = 12'h222;
rom[34896] = 12'h111;
rom[34897] = 12'h111;
rom[34898] = 12'h  0;
rom[34899] = 12'h  0;
rom[34900] = 12'h  0;
rom[34901] = 12'h  0;
rom[34902] = 12'h  0;
rom[34903] = 12'h  0;
rom[34904] = 12'h  0;
rom[34905] = 12'h  0;
rom[34906] = 12'h  0;
rom[34907] = 12'h  0;
rom[34908] = 12'h  0;
rom[34909] = 12'h  0;
rom[34910] = 12'h  0;
rom[34911] = 12'h  0;
rom[34912] = 12'h  0;
rom[34913] = 12'h  0;
rom[34914] = 12'h  0;
rom[34915] = 12'h  0;
rom[34916] = 12'h  0;
rom[34917] = 12'h  0;
rom[34918] = 12'h  0;
rom[34919] = 12'h  0;
rom[34920] = 12'h  0;
rom[34921] = 12'h  0;
rom[34922] = 12'h  0;
rom[34923] = 12'h  0;
rom[34924] = 12'h  0;
rom[34925] = 12'h  0;
rom[34926] = 12'h  0;
rom[34927] = 12'h  0;
rom[34928] = 12'h  0;
rom[34929] = 12'h  0;
rom[34930] = 12'h  0;
rom[34931] = 12'h  0;
rom[34932] = 12'h  0;
rom[34933] = 12'h  0;
rom[34934] = 12'h  0;
rom[34935] = 12'h  0;
rom[34936] = 12'h  0;
rom[34937] = 12'h  0;
rom[34938] = 12'h  0;
rom[34939] = 12'h  0;
rom[34940] = 12'h  0;
rom[34941] = 12'h  0;
rom[34942] = 12'h  0;
rom[34943] = 12'h  0;
rom[34944] = 12'h  0;
rom[34945] = 12'h  0;
rom[34946] = 12'h  0;
rom[34947] = 12'h  0;
rom[34948] = 12'h  0;
rom[34949] = 12'h  0;
rom[34950] = 12'h  0;
rom[34951] = 12'h  0;
rom[34952] = 12'h  0;
rom[34953] = 12'h  0;
rom[34954] = 12'h  0;
rom[34955] = 12'h  0;
rom[34956] = 12'h  0;
rom[34957] = 12'h  0;
rom[34958] = 12'h  0;
rom[34959] = 12'h  0;
rom[34960] = 12'h  0;
rom[34961] = 12'h  0;
rom[34962] = 12'h  0;
rom[34963] = 12'h  0;
rom[34964] = 12'h  0;
rom[34965] = 12'h  0;
rom[34966] = 12'h  0;
rom[34967] = 12'h  0;
rom[34968] = 12'h  0;
rom[34969] = 12'h  0;
rom[34970] = 12'h  0;
rom[34971] = 12'h  0;
rom[34972] = 12'h  0;
rom[34973] = 12'h  0;
rom[34974] = 12'h  0;
rom[34975] = 12'h  0;
rom[34976] = 12'h  0;
rom[34977] = 12'h  0;
rom[34978] = 12'h  0;
rom[34979] = 12'h  0;
rom[34980] = 12'h  0;
rom[34981] = 12'h  0;
rom[34982] = 12'h  0;
rom[34983] = 12'h  0;
rom[34984] = 12'h  0;
rom[34985] = 12'h  0;
rom[34986] = 12'h  0;
rom[34987] = 12'h  0;
rom[34988] = 12'h  0;
rom[34989] = 12'h  0;
rom[34990] = 12'h  0;
rom[34991] = 12'h  0;
rom[34992] = 12'h  0;
rom[34993] = 12'h  0;
rom[34994] = 12'h  0;
rom[34995] = 12'h  0;
rom[34996] = 12'h  0;
rom[34997] = 12'h  0;
rom[34998] = 12'h111;
rom[34999] = 12'h222;
rom[35000] = 12'h222;
rom[35001] = 12'h333;
rom[35002] = 12'h444;
rom[35003] = 12'h555;
rom[35004] = 12'h555;
rom[35005] = 12'h555;
rom[35006] = 12'h555;
rom[35007] = 12'h555;
rom[35008] = 12'h666;
rom[35009] = 12'h666;
rom[35010] = 12'h666;
rom[35011] = 12'h555;
rom[35012] = 12'h555;
rom[35013] = 12'h555;
rom[35014] = 12'h555;
rom[35015] = 12'h555;
rom[35016] = 12'h555;
rom[35017] = 12'h555;
rom[35018] = 12'h555;
rom[35019] = 12'h555;
rom[35020] = 12'h555;
rom[35021] = 12'h555;
rom[35022] = 12'h444;
rom[35023] = 12'h444;
rom[35024] = 12'h555;
rom[35025] = 12'h444;
rom[35026] = 12'h444;
rom[35027] = 12'h444;
rom[35028] = 12'h555;
rom[35029] = 12'h555;
rom[35030] = 12'h555;
rom[35031] = 12'h666;
rom[35032] = 12'h555;
rom[35033] = 12'h555;
rom[35034] = 12'h555;
rom[35035] = 12'h444;
rom[35036] = 12'h444;
rom[35037] = 12'h444;
rom[35038] = 12'h333;
rom[35039] = 12'h333;
rom[35040] = 12'h333;
rom[35041] = 12'h333;
rom[35042] = 12'h222;
rom[35043] = 12'h222;
rom[35044] = 12'h222;
rom[35045] = 12'h111;
rom[35046] = 12'h111;
rom[35047] = 12'h111;
rom[35048] = 12'h111;
rom[35049] = 12'h111;
rom[35050] = 12'h111;
rom[35051] = 12'h  0;
rom[35052] = 12'h  0;
rom[35053] = 12'h  0;
rom[35054] = 12'h  0;
rom[35055] = 12'h  0;
rom[35056] = 12'h  0;
rom[35057] = 12'h  0;
rom[35058] = 12'h  0;
rom[35059] = 12'h  0;
rom[35060] = 12'h  0;
rom[35061] = 12'h  0;
rom[35062] = 12'h  0;
rom[35063] = 12'h  0;
rom[35064] = 12'h  0;
rom[35065] = 12'h  0;
rom[35066] = 12'h  0;
rom[35067] = 12'h  0;
rom[35068] = 12'h  0;
rom[35069] = 12'h  0;
rom[35070] = 12'h  0;
rom[35071] = 12'h  0;
rom[35072] = 12'h  0;
rom[35073] = 12'h  0;
rom[35074] = 12'h  0;
rom[35075] = 12'h  0;
rom[35076] = 12'h  0;
rom[35077] = 12'h  0;
rom[35078] = 12'h  0;
rom[35079] = 12'h  0;
rom[35080] = 12'h  0;
rom[35081] = 12'h  0;
rom[35082] = 12'h111;
rom[35083] = 12'h111;
rom[35084] = 12'h111;
rom[35085] = 12'h222;
rom[35086] = 12'h333;
rom[35087] = 12'h333;
rom[35088] = 12'h433;
rom[35089] = 12'h333;
rom[35090] = 12'h333;
rom[35091] = 12'h333;
rom[35092] = 12'h444;
rom[35093] = 12'h444;
rom[35094] = 12'h555;
rom[35095] = 12'h555;
rom[35096] = 12'h666;
rom[35097] = 12'h777;
rom[35098] = 12'h898;
rom[35099] = 12'h999;
rom[35100] = 12'haaa;
rom[35101] = 12'haba;
rom[35102] = 12'hccc;
rom[35103] = 12'hddc;
rom[35104] = 12'hfee;
rom[35105] = 12'hffe;
rom[35106] = 12'hedc;
rom[35107] = 12'h987;
rom[35108] = 12'h543;
rom[35109] = 12'h421;
rom[35110] = 12'h310;
rom[35111] = 12'h210;
rom[35112] = 12'h200;
rom[35113] = 12'h100;
rom[35114] = 12'h100;
rom[35115] = 12'h  0;
rom[35116] = 12'h  0;
rom[35117] = 12'h  0;
rom[35118] = 12'h  0;
rom[35119] = 12'h  0;
rom[35120] = 12'h  0;
rom[35121] = 12'h  0;
rom[35122] = 12'h  0;
rom[35123] = 12'h  0;
rom[35124] = 12'h  0;
rom[35125] = 12'h  0;
rom[35126] = 12'h  0;
rom[35127] = 12'h  0;
rom[35128] = 12'h  0;
rom[35129] = 12'h  0;
rom[35130] = 12'h  0;
rom[35131] = 12'h  0;
rom[35132] = 12'h  0;
rom[35133] = 12'h  0;
rom[35134] = 12'h  0;
rom[35135] = 12'h  0;
rom[35136] = 12'h100;
rom[35137] = 12'h100;
rom[35138] = 12'h100;
rom[35139] = 12'h100;
rom[35140] = 12'h200;
rom[35141] = 12'h200;
rom[35142] = 12'h300;
rom[35143] = 12'h400;
rom[35144] = 12'h500;
rom[35145] = 12'h710;
rom[35146] = 12'h920;
rom[35147] = 12'hb30;
rom[35148] = 12'hd51;
rom[35149] = 12'hf51;
rom[35150] = 12'hf61;
rom[35151] = 12'hf60;
rom[35152] = 12'he70;
rom[35153] = 12'he91;
rom[35154] = 12'hfa3;
rom[35155] = 12'hfb4;
rom[35156] = 12'hea3;
rom[35157] = 12'ha70;
rom[35158] = 12'h850;
rom[35159] = 12'h850;
rom[35160] = 12'h740;
rom[35161] = 12'h730;
rom[35162] = 12'h620;
rom[35163] = 12'h520;
rom[35164] = 12'h520;
rom[35165] = 12'h420;
rom[35166] = 12'h420;
rom[35167] = 12'h310;
rom[35168] = 12'h310;
rom[35169] = 12'h210;
rom[35170] = 12'h210;
rom[35171] = 12'h210;
rom[35172] = 12'h210;
rom[35173] = 12'h211;
rom[35174] = 12'h211;
rom[35175] = 12'h222;
rom[35176] = 12'h323;
rom[35177] = 12'h333;
rom[35178] = 12'h333;
rom[35179] = 12'h334;
rom[35180] = 12'h444;
rom[35181] = 12'h545;
rom[35182] = 12'h656;
rom[35183] = 12'h667;
rom[35184] = 12'h777;
rom[35185] = 12'h777;
rom[35186] = 12'h777;
rom[35187] = 12'h888;
rom[35188] = 12'h888;
rom[35189] = 12'h888;
rom[35190] = 12'h999;
rom[35191] = 12'h999;
rom[35192] = 12'haaa;
rom[35193] = 12'haaa;
rom[35194] = 12'haaa;
rom[35195] = 12'haaa;
rom[35196] = 12'haaa;
rom[35197] = 12'haaa;
rom[35198] = 12'haaa;
rom[35199] = 12'hbbb;
rom[35200] = 12'h888;
rom[35201] = 12'h888;
rom[35202] = 12'h888;
rom[35203] = 12'h888;
rom[35204] = 12'h888;
rom[35205] = 12'h888;
rom[35206] = 12'h888;
rom[35207] = 12'h888;
rom[35208] = 12'h888;
rom[35209] = 12'h888;
rom[35210] = 12'h888;
rom[35211] = 12'h888;
rom[35212] = 12'h888;
rom[35213] = 12'h999;
rom[35214] = 12'h999;
rom[35215] = 12'h999;
rom[35216] = 12'h999;
rom[35217] = 12'h999;
rom[35218] = 12'h999;
rom[35219] = 12'haaa;
rom[35220] = 12'haaa;
rom[35221] = 12'haaa;
rom[35222] = 12'haaa;
rom[35223] = 12'haaa;
rom[35224] = 12'haaa;
rom[35225] = 12'haaa;
rom[35226] = 12'haaa;
rom[35227] = 12'haaa;
rom[35228] = 12'haaa;
rom[35229] = 12'haaa;
rom[35230] = 12'h999;
rom[35231] = 12'h999;
rom[35232] = 12'h999;
rom[35233] = 12'h999;
rom[35234] = 12'h999;
rom[35235] = 12'haaa;
rom[35236] = 12'haaa;
rom[35237] = 12'haaa;
rom[35238] = 12'haaa;
rom[35239] = 12'haaa;
rom[35240] = 12'haaa;
rom[35241] = 12'haaa;
rom[35242] = 12'haaa;
rom[35243] = 12'h999;
rom[35244] = 12'h999;
rom[35245] = 12'h999;
rom[35246] = 12'h999;
rom[35247] = 12'h999;
rom[35248] = 12'h999;
rom[35249] = 12'h888;
rom[35250] = 12'h888;
rom[35251] = 12'h888;
rom[35252] = 12'h777;
rom[35253] = 12'h777;
rom[35254] = 12'h777;
rom[35255] = 12'h777;
rom[35256] = 12'h777;
rom[35257] = 12'h777;
rom[35258] = 12'h777;
rom[35259] = 12'h777;
rom[35260] = 12'h777;
rom[35261] = 12'h777;
rom[35262] = 12'h777;
rom[35263] = 12'h777;
rom[35264] = 12'h777;
rom[35265] = 12'h777;
rom[35266] = 12'h777;
rom[35267] = 12'h777;
rom[35268] = 12'h666;
rom[35269] = 12'h777;
rom[35270] = 12'h777;
rom[35271] = 12'h888;
rom[35272] = 12'haaa;
rom[35273] = 12'haaa;
rom[35274] = 12'haaa;
rom[35275] = 12'h999;
rom[35276] = 12'h999;
rom[35277] = 12'h888;
rom[35278] = 12'h777;
rom[35279] = 12'h666;
rom[35280] = 12'h666;
rom[35281] = 12'h666;
rom[35282] = 12'h555;
rom[35283] = 12'h555;
rom[35284] = 12'h444;
rom[35285] = 12'h444;
rom[35286] = 12'h444;
rom[35287] = 12'h444;
rom[35288] = 12'h333;
rom[35289] = 12'h333;
rom[35290] = 12'h333;
rom[35291] = 12'h222;
rom[35292] = 12'h222;
rom[35293] = 12'h222;
rom[35294] = 12'h222;
rom[35295] = 12'h111;
rom[35296] = 12'h111;
rom[35297] = 12'h111;
rom[35298] = 12'h111;
rom[35299] = 12'h  0;
rom[35300] = 12'h  0;
rom[35301] = 12'h  0;
rom[35302] = 12'h  0;
rom[35303] = 12'h  0;
rom[35304] = 12'h  0;
rom[35305] = 12'h  0;
rom[35306] = 12'h  0;
rom[35307] = 12'h  0;
rom[35308] = 12'h  0;
rom[35309] = 12'h  0;
rom[35310] = 12'h  0;
rom[35311] = 12'h  0;
rom[35312] = 12'h  0;
rom[35313] = 12'h  0;
rom[35314] = 12'h  0;
rom[35315] = 12'h  0;
rom[35316] = 12'h  0;
rom[35317] = 12'h  0;
rom[35318] = 12'h  0;
rom[35319] = 12'h  0;
rom[35320] = 12'h  0;
rom[35321] = 12'h  0;
rom[35322] = 12'h  0;
rom[35323] = 12'h  0;
rom[35324] = 12'h  0;
rom[35325] = 12'h  0;
rom[35326] = 12'h  0;
rom[35327] = 12'h  0;
rom[35328] = 12'h  0;
rom[35329] = 12'h  0;
rom[35330] = 12'h  0;
rom[35331] = 12'h  0;
rom[35332] = 12'h  0;
rom[35333] = 12'h  0;
rom[35334] = 12'h  0;
rom[35335] = 12'h  0;
rom[35336] = 12'h  0;
rom[35337] = 12'h  0;
rom[35338] = 12'h  0;
rom[35339] = 12'h  0;
rom[35340] = 12'h  0;
rom[35341] = 12'h  0;
rom[35342] = 12'h  0;
rom[35343] = 12'h  0;
rom[35344] = 12'h  0;
rom[35345] = 12'h  0;
rom[35346] = 12'h  0;
rom[35347] = 12'h  0;
rom[35348] = 12'h  0;
rom[35349] = 12'h  0;
rom[35350] = 12'h  0;
rom[35351] = 12'h  0;
rom[35352] = 12'h  0;
rom[35353] = 12'h  0;
rom[35354] = 12'h  0;
rom[35355] = 12'h  0;
rom[35356] = 12'h  0;
rom[35357] = 12'h  0;
rom[35358] = 12'h  0;
rom[35359] = 12'h  0;
rom[35360] = 12'h  0;
rom[35361] = 12'h  0;
rom[35362] = 12'h  0;
rom[35363] = 12'h  0;
rom[35364] = 12'h  0;
rom[35365] = 12'h  0;
rom[35366] = 12'h  0;
rom[35367] = 12'h  0;
rom[35368] = 12'h  0;
rom[35369] = 12'h  0;
rom[35370] = 12'h  0;
rom[35371] = 12'h  0;
rom[35372] = 12'h  0;
rom[35373] = 12'h  0;
rom[35374] = 12'h  0;
rom[35375] = 12'h  0;
rom[35376] = 12'h  0;
rom[35377] = 12'h  0;
rom[35378] = 12'h  0;
rom[35379] = 12'h  0;
rom[35380] = 12'h  0;
rom[35381] = 12'h  0;
rom[35382] = 12'h  0;
rom[35383] = 12'h  0;
rom[35384] = 12'h  0;
rom[35385] = 12'h  0;
rom[35386] = 12'h  0;
rom[35387] = 12'h  0;
rom[35388] = 12'h  0;
rom[35389] = 12'h  0;
rom[35390] = 12'h  0;
rom[35391] = 12'h  0;
rom[35392] = 12'h  0;
rom[35393] = 12'h  0;
rom[35394] = 12'h  0;
rom[35395] = 12'h  0;
rom[35396] = 12'h  0;
rom[35397] = 12'h111;
rom[35398] = 12'h111;
rom[35399] = 12'h222;
rom[35400] = 12'h333;
rom[35401] = 12'h444;
rom[35402] = 12'h444;
rom[35403] = 12'h444;
rom[35404] = 12'h444;
rom[35405] = 12'h444;
rom[35406] = 12'h555;
rom[35407] = 12'h555;
rom[35408] = 12'h555;
rom[35409] = 12'h555;
rom[35410] = 12'h555;
rom[35411] = 12'h555;
rom[35412] = 12'h555;
rom[35413] = 12'h555;
rom[35414] = 12'h555;
rom[35415] = 12'h555;
rom[35416] = 12'h444;
rom[35417] = 12'h444;
rom[35418] = 12'h555;
rom[35419] = 12'h555;
rom[35420] = 12'h444;
rom[35421] = 12'h444;
rom[35422] = 12'h444;
rom[35423] = 12'h444;
rom[35424] = 12'h444;
rom[35425] = 12'h444;
rom[35426] = 12'h444;
rom[35427] = 12'h444;
rom[35428] = 12'h555;
rom[35429] = 12'h555;
rom[35430] = 12'h555;
rom[35431] = 12'h666;
rom[35432] = 12'h555;
rom[35433] = 12'h555;
rom[35434] = 12'h444;
rom[35435] = 12'h444;
rom[35436] = 12'h444;
rom[35437] = 12'h333;
rom[35438] = 12'h333;
rom[35439] = 12'h333;
rom[35440] = 12'h222;
rom[35441] = 12'h222;
rom[35442] = 12'h222;
rom[35443] = 12'h222;
rom[35444] = 12'h222;
rom[35445] = 12'h222;
rom[35446] = 12'h111;
rom[35447] = 12'h111;
rom[35448] = 12'h111;
rom[35449] = 12'h111;
rom[35450] = 12'h111;
rom[35451] = 12'h  0;
rom[35452] = 12'h  0;
rom[35453] = 12'h  0;
rom[35454] = 12'h  0;
rom[35455] = 12'h  0;
rom[35456] = 12'h  0;
rom[35457] = 12'h  0;
rom[35458] = 12'h  0;
rom[35459] = 12'h  0;
rom[35460] = 12'h  0;
rom[35461] = 12'h  0;
rom[35462] = 12'h  0;
rom[35463] = 12'h  0;
rom[35464] = 12'h  0;
rom[35465] = 12'h  0;
rom[35466] = 12'h  0;
rom[35467] = 12'h  0;
rom[35468] = 12'h  0;
rom[35469] = 12'h  0;
rom[35470] = 12'h  0;
rom[35471] = 12'h  0;
rom[35472] = 12'h  0;
rom[35473] = 12'h  0;
rom[35474] = 12'h  0;
rom[35475] = 12'h  0;
rom[35476] = 12'h  0;
rom[35477] = 12'h  0;
rom[35478] = 12'h  0;
rom[35479] = 12'h  0;
rom[35480] = 12'h  0;
rom[35481] = 12'h  0;
rom[35482] = 12'h111;
rom[35483] = 12'h111;
rom[35484] = 12'h222;
rom[35485] = 12'h222;
rom[35486] = 12'h333;
rom[35487] = 12'h333;
rom[35488] = 12'h444;
rom[35489] = 12'h333;
rom[35490] = 12'h333;
rom[35491] = 12'h333;
rom[35492] = 12'h444;
rom[35493] = 12'h455;
rom[35494] = 12'h555;
rom[35495] = 12'h666;
rom[35496] = 12'h676;
rom[35497] = 12'h999;
rom[35498] = 12'h898;
rom[35499] = 12'h898;
rom[35500] = 12'hbcb;
rom[35501] = 12'hccc;
rom[35502] = 12'hccc;
rom[35503] = 12'heed;
rom[35504] = 12'hffe;
rom[35505] = 12'hfed;
rom[35506] = 12'ha97;
rom[35507] = 12'h532;
rom[35508] = 12'h421;
rom[35509] = 12'h421;
rom[35510] = 12'h310;
rom[35511] = 12'h310;
rom[35512] = 12'h200;
rom[35513] = 12'h200;
rom[35514] = 12'h100;
rom[35515] = 12'h100;
rom[35516] = 12'h  0;
rom[35517] = 12'h  0;
rom[35518] = 12'h  0;
rom[35519] = 12'h  0;
rom[35520] = 12'h  0;
rom[35521] = 12'h  0;
rom[35522] = 12'h  0;
rom[35523] = 12'h  0;
rom[35524] = 12'h  0;
rom[35525] = 12'h  0;
rom[35526] = 12'h  0;
rom[35527] = 12'h  0;
rom[35528] = 12'h  0;
rom[35529] = 12'h  0;
rom[35530] = 12'h  0;
rom[35531] = 12'h  0;
rom[35532] = 12'h  0;
rom[35533] = 12'h  0;
rom[35534] = 12'h100;
rom[35535] = 12'h100;
rom[35536] = 12'h100;
rom[35537] = 12'h100;
rom[35538] = 12'h100;
rom[35539] = 12'h200;
rom[35540] = 12'h200;
rom[35541] = 12'h300;
rom[35542] = 12'h410;
rom[35543] = 12'h510;
rom[35544] = 12'h610;
rom[35545] = 12'h810;
rom[35546] = 12'ha30;
rom[35547] = 12'hc40;
rom[35548] = 12'hd51;
rom[35549] = 12'hf51;
rom[35550] = 12'hf61;
rom[35551] = 12'hf60;
rom[35552] = 12'hf80;
rom[35553] = 12'hfa2;
rom[35554] = 12'hfb4;
rom[35555] = 12'hfb4;
rom[35556] = 12'hc82;
rom[35557] = 12'h960;
rom[35558] = 12'h850;
rom[35559] = 12'h850;
rom[35560] = 12'h730;
rom[35561] = 12'h730;
rom[35562] = 12'h630;
rom[35563] = 12'h620;
rom[35564] = 12'h520;
rom[35565] = 12'h420;
rom[35566] = 12'h420;
rom[35567] = 12'h320;
rom[35568] = 12'h310;
rom[35569] = 12'h210;
rom[35570] = 12'h210;
rom[35571] = 12'h210;
rom[35572] = 12'h210;
rom[35573] = 12'h211;
rom[35574] = 12'h221;
rom[35575] = 12'h222;
rom[35576] = 12'h323;
rom[35577] = 12'h323;
rom[35578] = 12'h333;
rom[35579] = 12'h333;
rom[35580] = 12'h444;
rom[35581] = 12'h545;
rom[35582] = 12'h556;
rom[35583] = 12'h666;
rom[35584] = 12'h767;
rom[35585] = 12'h777;
rom[35586] = 12'h777;
rom[35587] = 12'h888;
rom[35588] = 12'h888;
rom[35589] = 12'h999;
rom[35590] = 12'h999;
rom[35591] = 12'h999;
rom[35592] = 12'haaa;
rom[35593] = 12'haaa;
rom[35594] = 12'haaa;
rom[35595] = 12'haaa;
rom[35596] = 12'haaa;
rom[35597] = 12'haaa;
rom[35598] = 12'haaa;
rom[35599] = 12'haaa;
rom[35600] = 12'h888;
rom[35601] = 12'h888;
rom[35602] = 12'h888;
rom[35603] = 12'h888;
rom[35604] = 12'h888;
rom[35605] = 12'h888;
rom[35606] = 12'h888;
rom[35607] = 12'h888;
rom[35608] = 12'h777;
rom[35609] = 12'h777;
rom[35610] = 12'h777;
rom[35611] = 12'h888;
rom[35612] = 12'h888;
rom[35613] = 12'h888;
rom[35614] = 12'h888;
rom[35615] = 12'h888;
rom[35616] = 12'h999;
rom[35617] = 12'h999;
rom[35618] = 12'h999;
rom[35619] = 12'h999;
rom[35620] = 12'haaa;
rom[35621] = 12'haaa;
rom[35622] = 12'haaa;
rom[35623] = 12'haaa;
rom[35624] = 12'haaa;
rom[35625] = 12'haaa;
rom[35626] = 12'haaa;
rom[35627] = 12'haaa;
rom[35628] = 12'haaa;
rom[35629] = 12'haaa;
rom[35630] = 12'haaa;
rom[35631] = 12'haaa;
rom[35632] = 12'haaa;
rom[35633] = 12'haaa;
rom[35634] = 12'haaa;
rom[35635] = 12'haaa;
rom[35636] = 12'haaa;
rom[35637] = 12'haaa;
rom[35638] = 12'haaa;
rom[35639] = 12'haaa;
rom[35640] = 12'haaa;
rom[35641] = 12'haaa;
rom[35642] = 12'haaa;
rom[35643] = 12'haaa;
rom[35644] = 12'h999;
rom[35645] = 12'h999;
rom[35646] = 12'h999;
rom[35647] = 12'h999;
rom[35648] = 12'h999;
rom[35649] = 12'h888;
rom[35650] = 12'h888;
rom[35651] = 12'h888;
rom[35652] = 12'h888;
rom[35653] = 12'h777;
rom[35654] = 12'h777;
rom[35655] = 12'h777;
rom[35656] = 12'h777;
rom[35657] = 12'h777;
rom[35658] = 12'h777;
rom[35659] = 12'h777;
rom[35660] = 12'h777;
rom[35661] = 12'h777;
rom[35662] = 12'h777;
rom[35663] = 12'h777;
rom[35664] = 12'h777;
rom[35665] = 12'h777;
rom[35666] = 12'h777;
rom[35667] = 12'h777;
rom[35668] = 12'h777;
rom[35669] = 12'h777;
rom[35670] = 12'h777;
rom[35671] = 12'h888;
rom[35672] = 12'h888;
rom[35673] = 12'h999;
rom[35674] = 12'h999;
rom[35675] = 12'haaa;
rom[35676] = 12'h999;
rom[35677] = 12'h999;
rom[35678] = 12'h888;
rom[35679] = 12'h777;
rom[35680] = 12'h666;
rom[35681] = 12'h666;
rom[35682] = 12'h555;
rom[35683] = 12'h555;
rom[35684] = 12'h444;
rom[35685] = 12'h444;
rom[35686] = 12'h333;
rom[35687] = 12'h333;
rom[35688] = 12'h333;
rom[35689] = 12'h333;
rom[35690] = 12'h333;
rom[35691] = 12'h222;
rom[35692] = 12'h222;
rom[35693] = 12'h222;
rom[35694] = 12'h222;
rom[35695] = 12'h222;
rom[35696] = 12'h111;
rom[35697] = 12'h111;
rom[35698] = 12'h111;
rom[35699] = 12'h111;
rom[35700] = 12'h  0;
rom[35701] = 12'h  0;
rom[35702] = 12'h  0;
rom[35703] = 12'h  0;
rom[35704] = 12'h  0;
rom[35705] = 12'h  0;
rom[35706] = 12'h  0;
rom[35707] = 12'h  0;
rom[35708] = 12'h  0;
rom[35709] = 12'h  0;
rom[35710] = 12'h  0;
rom[35711] = 12'h  0;
rom[35712] = 12'h  0;
rom[35713] = 12'h  0;
rom[35714] = 12'h  0;
rom[35715] = 12'h  0;
rom[35716] = 12'h  0;
rom[35717] = 12'h  0;
rom[35718] = 12'h  0;
rom[35719] = 12'h  0;
rom[35720] = 12'h  0;
rom[35721] = 12'h  0;
rom[35722] = 12'h  0;
rom[35723] = 12'h  0;
rom[35724] = 12'h  0;
rom[35725] = 12'h  0;
rom[35726] = 12'h  0;
rom[35727] = 12'h  0;
rom[35728] = 12'h  0;
rom[35729] = 12'h  0;
rom[35730] = 12'h  0;
rom[35731] = 12'h  0;
rom[35732] = 12'h  0;
rom[35733] = 12'h  0;
rom[35734] = 12'h  0;
rom[35735] = 12'h  0;
rom[35736] = 12'h  0;
rom[35737] = 12'h  0;
rom[35738] = 12'h  0;
rom[35739] = 12'h  0;
rom[35740] = 12'h  0;
rom[35741] = 12'h  0;
rom[35742] = 12'h  0;
rom[35743] = 12'h  0;
rom[35744] = 12'h  0;
rom[35745] = 12'h  0;
rom[35746] = 12'h  0;
rom[35747] = 12'h  0;
rom[35748] = 12'h  0;
rom[35749] = 12'h  0;
rom[35750] = 12'h  0;
rom[35751] = 12'h  0;
rom[35752] = 12'h  0;
rom[35753] = 12'h  0;
rom[35754] = 12'h  0;
rom[35755] = 12'h  0;
rom[35756] = 12'h  0;
rom[35757] = 12'h  0;
rom[35758] = 12'h  0;
rom[35759] = 12'h  0;
rom[35760] = 12'h  0;
rom[35761] = 12'h  0;
rom[35762] = 12'h  0;
rom[35763] = 12'h  0;
rom[35764] = 12'h  0;
rom[35765] = 12'h  0;
rom[35766] = 12'h  0;
rom[35767] = 12'h  0;
rom[35768] = 12'h  0;
rom[35769] = 12'h  0;
rom[35770] = 12'h  0;
rom[35771] = 12'h  0;
rom[35772] = 12'h  0;
rom[35773] = 12'h  0;
rom[35774] = 12'h  0;
rom[35775] = 12'h  0;
rom[35776] = 12'h  0;
rom[35777] = 12'h  0;
rom[35778] = 12'h  0;
rom[35779] = 12'h  0;
rom[35780] = 12'h  0;
rom[35781] = 12'h  0;
rom[35782] = 12'h  0;
rom[35783] = 12'h  0;
rom[35784] = 12'h  0;
rom[35785] = 12'h  0;
rom[35786] = 12'h  0;
rom[35787] = 12'h  0;
rom[35788] = 12'h  0;
rom[35789] = 12'h  0;
rom[35790] = 12'h  0;
rom[35791] = 12'h  0;
rom[35792] = 12'h  0;
rom[35793] = 12'h  0;
rom[35794] = 12'h  0;
rom[35795] = 12'h  0;
rom[35796] = 12'h111;
rom[35797] = 12'h111;
rom[35798] = 12'h222;
rom[35799] = 12'h222;
rom[35800] = 12'h333;
rom[35801] = 12'h444;
rom[35802] = 12'h444;
rom[35803] = 12'h444;
rom[35804] = 12'h444;
rom[35805] = 12'h444;
rom[35806] = 12'h444;
rom[35807] = 12'h555;
rom[35808] = 12'h555;
rom[35809] = 12'h555;
rom[35810] = 12'h555;
rom[35811] = 12'h555;
rom[35812] = 12'h555;
rom[35813] = 12'h555;
rom[35814] = 12'h555;
rom[35815] = 12'h555;
rom[35816] = 12'h444;
rom[35817] = 12'h444;
rom[35818] = 12'h444;
rom[35819] = 12'h444;
rom[35820] = 12'h444;
rom[35821] = 12'h444;
rom[35822] = 12'h444;
rom[35823] = 12'h444;
rom[35824] = 12'h444;
rom[35825] = 12'h444;
rom[35826] = 12'h444;
rom[35827] = 12'h444;
rom[35828] = 12'h555;
rom[35829] = 12'h555;
rom[35830] = 12'h555;
rom[35831] = 12'h555;
rom[35832] = 12'h555;
rom[35833] = 12'h555;
rom[35834] = 12'h444;
rom[35835] = 12'h444;
rom[35836] = 12'h444;
rom[35837] = 12'h333;
rom[35838] = 12'h333;
rom[35839] = 12'h333;
rom[35840] = 12'h222;
rom[35841] = 12'h222;
rom[35842] = 12'h222;
rom[35843] = 12'h222;
rom[35844] = 12'h222;
rom[35845] = 12'h222;
rom[35846] = 12'h111;
rom[35847] = 12'h111;
rom[35848] = 12'h111;
rom[35849] = 12'h111;
rom[35850] = 12'h  0;
rom[35851] = 12'h  0;
rom[35852] = 12'h  0;
rom[35853] = 12'h  0;
rom[35854] = 12'h  0;
rom[35855] = 12'h  0;
rom[35856] = 12'h  0;
rom[35857] = 12'h  0;
rom[35858] = 12'h  0;
rom[35859] = 12'h  0;
rom[35860] = 12'h  0;
rom[35861] = 12'h  0;
rom[35862] = 12'h  0;
rom[35863] = 12'h  0;
rom[35864] = 12'h  0;
rom[35865] = 12'h  0;
rom[35866] = 12'h  0;
rom[35867] = 12'h  0;
rom[35868] = 12'h  0;
rom[35869] = 12'h  0;
rom[35870] = 12'h  0;
rom[35871] = 12'h  0;
rom[35872] = 12'h  0;
rom[35873] = 12'h  0;
rom[35874] = 12'h  0;
rom[35875] = 12'h  0;
rom[35876] = 12'h  0;
rom[35877] = 12'h  0;
rom[35878] = 12'h  0;
rom[35879] = 12'h  0;
rom[35880] = 12'h  0;
rom[35881] = 12'h111;
rom[35882] = 12'h111;
rom[35883] = 12'h111;
rom[35884] = 12'h222;
rom[35885] = 12'h333;
rom[35886] = 12'h333;
rom[35887] = 12'h433;
rom[35888] = 12'h434;
rom[35889] = 12'h333;
rom[35890] = 12'h333;
rom[35891] = 12'h444;
rom[35892] = 12'h444;
rom[35893] = 12'h555;
rom[35894] = 12'h566;
rom[35895] = 12'h676;
rom[35896] = 12'h777;
rom[35897] = 12'h899;
rom[35898] = 12'h999;
rom[35899] = 12'haa9;
rom[35900] = 12'hccb;
rom[35901] = 12'hccc;
rom[35902] = 12'hddc;
rom[35903] = 12'hffe;
rom[35904] = 12'hffe;
rom[35905] = 12'hdba;
rom[35906] = 12'h864;
rom[35907] = 12'h521;
rom[35908] = 12'h420;
rom[35909] = 12'h410;
rom[35910] = 12'h310;
rom[35911] = 12'h310;
rom[35912] = 12'h300;
rom[35913] = 12'h200;
rom[35914] = 12'h100;
rom[35915] = 12'h100;
rom[35916] = 12'h  0;
rom[35917] = 12'h  0;
rom[35918] = 12'h  0;
rom[35919] = 12'h  0;
rom[35920] = 12'h  0;
rom[35921] = 12'h  0;
rom[35922] = 12'h  0;
rom[35923] = 12'h  0;
rom[35924] = 12'h  0;
rom[35925] = 12'h  0;
rom[35926] = 12'h  0;
rom[35927] = 12'h  0;
rom[35928] = 12'h  0;
rom[35929] = 12'h  0;
rom[35930] = 12'h  0;
rom[35931] = 12'h  0;
rom[35932] = 12'h  0;
rom[35933] = 12'h  0;
rom[35934] = 12'h100;
rom[35935] = 12'h100;
rom[35936] = 12'h100;
rom[35937] = 12'h100;
rom[35938] = 12'h200;
rom[35939] = 12'h200;
rom[35940] = 12'h300;
rom[35941] = 12'h400;
rom[35942] = 12'h510;
rom[35943] = 12'h610;
rom[35944] = 12'h710;
rom[35945] = 12'h920;
rom[35946] = 12'hb30;
rom[35947] = 12'hc40;
rom[35948] = 12'he50;
rom[35949] = 12'hf61;
rom[35950] = 12'hf61;
rom[35951] = 12'hf60;
rom[35952] = 12'he81;
rom[35953] = 12'hfa2;
rom[35954] = 12'hfb4;
rom[35955] = 12'hea3;
rom[35956] = 12'hb71;
rom[35957] = 12'h950;
rom[35958] = 12'h840;
rom[35959] = 12'h740;
rom[35960] = 12'h730;
rom[35961] = 12'h730;
rom[35962] = 12'h630;
rom[35963] = 12'h630;
rom[35964] = 12'h520;
rom[35965] = 12'h420;
rom[35966] = 12'h420;
rom[35967] = 12'h420;
rom[35968] = 12'h320;
rom[35969] = 12'h320;
rom[35970] = 12'h310;
rom[35971] = 12'h210;
rom[35972] = 12'h210;
rom[35973] = 12'h211;
rom[35974] = 12'h221;
rom[35975] = 12'h222;
rom[35976] = 12'h322;
rom[35977] = 12'h223;
rom[35978] = 12'h333;
rom[35979] = 12'h333;
rom[35980] = 12'h444;
rom[35981] = 12'h445;
rom[35982] = 12'h556;
rom[35983] = 12'h666;
rom[35984] = 12'h767;
rom[35985] = 12'h777;
rom[35986] = 12'h777;
rom[35987] = 12'h888;
rom[35988] = 12'h888;
rom[35989] = 12'h999;
rom[35990] = 12'h999;
rom[35991] = 12'h999;
rom[35992] = 12'haaa;
rom[35993] = 12'haaa;
rom[35994] = 12'haaa;
rom[35995] = 12'haaa;
rom[35996] = 12'haaa;
rom[35997] = 12'haaa;
rom[35998] = 12'haaa;
rom[35999] = 12'haaa;
rom[36000] = 12'h888;
rom[36001] = 12'h888;
rom[36002] = 12'h888;
rom[36003] = 12'h888;
rom[36004] = 12'h888;
rom[36005] = 12'h777;
rom[36006] = 12'h777;
rom[36007] = 12'h777;
rom[36008] = 12'h777;
rom[36009] = 12'h777;
rom[36010] = 12'h777;
rom[36011] = 12'h888;
rom[36012] = 12'h888;
rom[36013] = 12'h888;
rom[36014] = 12'h888;
rom[36015] = 12'h888;
rom[36016] = 12'h888;
rom[36017] = 12'h888;
rom[36018] = 12'h999;
rom[36019] = 12'h999;
rom[36020] = 12'h999;
rom[36021] = 12'h999;
rom[36022] = 12'haaa;
rom[36023] = 12'haaa;
rom[36024] = 12'haaa;
rom[36025] = 12'haaa;
rom[36026] = 12'haaa;
rom[36027] = 12'haaa;
rom[36028] = 12'haaa;
rom[36029] = 12'haaa;
rom[36030] = 12'haaa;
rom[36031] = 12'haaa;
rom[36032] = 12'haaa;
rom[36033] = 12'haaa;
rom[36034] = 12'haaa;
rom[36035] = 12'haaa;
rom[36036] = 12'haaa;
rom[36037] = 12'haaa;
rom[36038] = 12'haaa;
rom[36039] = 12'haaa;
rom[36040] = 12'haaa;
rom[36041] = 12'haaa;
rom[36042] = 12'haaa;
rom[36043] = 12'haaa;
rom[36044] = 12'haaa;
rom[36045] = 12'haaa;
rom[36046] = 12'h999;
rom[36047] = 12'h999;
rom[36048] = 12'h999;
rom[36049] = 12'h999;
rom[36050] = 12'h999;
rom[36051] = 12'h888;
rom[36052] = 12'h888;
rom[36053] = 12'h888;
rom[36054] = 12'h888;
rom[36055] = 12'h888;
rom[36056] = 12'h888;
rom[36057] = 12'h888;
rom[36058] = 12'h777;
rom[36059] = 12'h777;
rom[36060] = 12'h777;
rom[36061] = 12'h777;
rom[36062] = 12'h777;
rom[36063] = 12'h777;
rom[36064] = 12'h777;
rom[36065] = 12'h777;
rom[36066] = 12'h888;
rom[36067] = 12'h888;
rom[36068] = 12'h777;
rom[36069] = 12'h777;
rom[36070] = 12'h777;
rom[36071] = 12'h777;
rom[36072] = 12'h777;
rom[36073] = 12'h888;
rom[36074] = 12'h888;
rom[36075] = 12'h999;
rom[36076] = 12'haaa;
rom[36077] = 12'haaa;
rom[36078] = 12'h999;
rom[36079] = 12'h888;
rom[36080] = 12'h777;
rom[36081] = 12'h666;
rom[36082] = 12'h555;
rom[36083] = 12'h555;
rom[36084] = 12'h444;
rom[36085] = 12'h444;
rom[36086] = 12'h444;
rom[36087] = 12'h333;
rom[36088] = 12'h333;
rom[36089] = 12'h333;
rom[36090] = 12'h333;
rom[36091] = 12'h222;
rom[36092] = 12'h222;
rom[36093] = 12'h222;
rom[36094] = 12'h222;
rom[36095] = 12'h222;
rom[36096] = 12'h222;
rom[36097] = 12'h222;
rom[36098] = 12'h111;
rom[36099] = 12'h111;
rom[36100] = 12'h111;
rom[36101] = 12'h  0;
rom[36102] = 12'h  0;
rom[36103] = 12'h  0;
rom[36104] = 12'h  0;
rom[36105] = 12'h  0;
rom[36106] = 12'h  0;
rom[36107] = 12'h  0;
rom[36108] = 12'h  0;
rom[36109] = 12'h  0;
rom[36110] = 12'h  0;
rom[36111] = 12'h  0;
rom[36112] = 12'h  0;
rom[36113] = 12'h  0;
rom[36114] = 12'h  0;
rom[36115] = 12'h  0;
rom[36116] = 12'h  0;
rom[36117] = 12'h  0;
rom[36118] = 12'h  0;
rom[36119] = 12'h  0;
rom[36120] = 12'h  0;
rom[36121] = 12'h  0;
rom[36122] = 12'h  0;
rom[36123] = 12'h  0;
rom[36124] = 12'h  0;
rom[36125] = 12'h  0;
rom[36126] = 12'h  0;
rom[36127] = 12'h  0;
rom[36128] = 12'h  0;
rom[36129] = 12'h  0;
rom[36130] = 12'h  0;
rom[36131] = 12'h  0;
rom[36132] = 12'h  0;
rom[36133] = 12'h  0;
rom[36134] = 12'h  0;
rom[36135] = 12'h  0;
rom[36136] = 12'h  0;
rom[36137] = 12'h  0;
rom[36138] = 12'h  0;
rom[36139] = 12'h  0;
rom[36140] = 12'h  0;
rom[36141] = 12'h  0;
rom[36142] = 12'h  0;
rom[36143] = 12'h  0;
rom[36144] = 12'h  0;
rom[36145] = 12'h  0;
rom[36146] = 12'h  0;
rom[36147] = 12'h  0;
rom[36148] = 12'h  0;
rom[36149] = 12'h  0;
rom[36150] = 12'h  0;
rom[36151] = 12'h  0;
rom[36152] = 12'h  0;
rom[36153] = 12'h  0;
rom[36154] = 12'h  0;
rom[36155] = 12'h  0;
rom[36156] = 12'h  0;
rom[36157] = 12'h  0;
rom[36158] = 12'h  0;
rom[36159] = 12'h  0;
rom[36160] = 12'h  0;
rom[36161] = 12'h  0;
rom[36162] = 12'h  0;
rom[36163] = 12'h  0;
rom[36164] = 12'h  0;
rom[36165] = 12'h  0;
rom[36166] = 12'h  0;
rom[36167] = 12'h  0;
rom[36168] = 12'h  0;
rom[36169] = 12'h  0;
rom[36170] = 12'h  0;
rom[36171] = 12'h  0;
rom[36172] = 12'h  0;
rom[36173] = 12'h  0;
rom[36174] = 12'h  0;
rom[36175] = 12'h  0;
rom[36176] = 12'h  0;
rom[36177] = 12'h  0;
rom[36178] = 12'h  0;
rom[36179] = 12'h  0;
rom[36180] = 12'h  0;
rom[36181] = 12'h  0;
rom[36182] = 12'h  0;
rom[36183] = 12'h  0;
rom[36184] = 12'h  0;
rom[36185] = 12'h  0;
rom[36186] = 12'h  0;
rom[36187] = 12'h  0;
rom[36188] = 12'h  0;
rom[36189] = 12'h  0;
rom[36190] = 12'h  0;
rom[36191] = 12'h  0;
rom[36192] = 12'h  0;
rom[36193] = 12'h  0;
rom[36194] = 12'h  0;
rom[36195] = 12'h111;
rom[36196] = 12'h111;
rom[36197] = 12'h111;
rom[36198] = 12'h222;
rom[36199] = 12'h222;
rom[36200] = 12'h333;
rom[36201] = 12'h444;
rom[36202] = 12'h444;
rom[36203] = 12'h444;
rom[36204] = 12'h444;
rom[36205] = 12'h444;
rom[36206] = 12'h444;
rom[36207] = 12'h555;
rom[36208] = 12'h555;
rom[36209] = 12'h555;
rom[36210] = 12'h555;
rom[36211] = 12'h555;
rom[36212] = 12'h555;
rom[36213] = 12'h555;
rom[36214] = 12'h555;
rom[36215] = 12'h444;
rom[36216] = 12'h444;
rom[36217] = 12'h444;
rom[36218] = 12'h444;
rom[36219] = 12'h444;
rom[36220] = 12'h444;
rom[36221] = 12'h444;
rom[36222] = 12'h444;
rom[36223] = 12'h444;
rom[36224] = 12'h444;
rom[36225] = 12'h444;
rom[36226] = 12'h444;
rom[36227] = 12'h444;
rom[36228] = 12'h555;
rom[36229] = 12'h555;
rom[36230] = 12'h555;
rom[36231] = 12'h555;
rom[36232] = 12'h555;
rom[36233] = 12'h555;
rom[36234] = 12'h444;
rom[36235] = 12'h444;
rom[36236] = 12'h333;
rom[36237] = 12'h333;
rom[36238] = 12'h333;
rom[36239] = 12'h333;
rom[36240] = 12'h222;
rom[36241] = 12'h222;
rom[36242] = 12'h222;
rom[36243] = 12'h222;
rom[36244] = 12'h222;
rom[36245] = 12'h222;
rom[36246] = 12'h111;
rom[36247] = 12'h111;
rom[36248] = 12'h111;
rom[36249] = 12'h111;
rom[36250] = 12'h  0;
rom[36251] = 12'h  0;
rom[36252] = 12'h  0;
rom[36253] = 12'h  0;
rom[36254] = 12'h  0;
rom[36255] = 12'h  0;
rom[36256] = 12'h  0;
rom[36257] = 12'h  0;
rom[36258] = 12'h  0;
rom[36259] = 12'h  0;
rom[36260] = 12'h  0;
rom[36261] = 12'h  0;
rom[36262] = 12'h  0;
rom[36263] = 12'h  0;
rom[36264] = 12'h  0;
rom[36265] = 12'h  0;
rom[36266] = 12'h  0;
rom[36267] = 12'h  0;
rom[36268] = 12'h  0;
rom[36269] = 12'h  0;
rom[36270] = 12'h  0;
rom[36271] = 12'h  0;
rom[36272] = 12'h  0;
rom[36273] = 12'h  0;
rom[36274] = 12'h  0;
rom[36275] = 12'h  0;
rom[36276] = 12'h  0;
rom[36277] = 12'h  0;
rom[36278] = 12'h  0;
rom[36279] = 12'h111;
rom[36280] = 12'h111;
rom[36281] = 12'h111;
rom[36282] = 12'h111;
rom[36283] = 12'h111;
rom[36284] = 12'h222;
rom[36285] = 12'h333;
rom[36286] = 12'h444;
rom[36287] = 12'h444;
rom[36288] = 12'h433;
rom[36289] = 12'h433;
rom[36290] = 12'h444;
rom[36291] = 12'h444;
rom[36292] = 12'h555;
rom[36293] = 12'h666;
rom[36294] = 12'h676;
rom[36295] = 12'h777;
rom[36296] = 12'h888;
rom[36297] = 12'h898;
rom[36298] = 12'haaa;
rom[36299] = 12'hbcb;
rom[36300] = 12'hccc;
rom[36301] = 12'hccc;
rom[36302] = 12'heed;
rom[36303] = 12'hfff;
rom[36304] = 12'hfec;
rom[36305] = 12'ha76;
rom[36306] = 12'h531;
rom[36307] = 12'h521;
rom[36308] = 12'h521;
rom[36309] = 12'h410;
rom[36310] = 12'h410;
rom[36311] = 12'h410;
rom[36312] = 12'h300;
rom[36313] = 12'h300;
rom[36314] = 12'h200;
rom[36315] = 12'h100;
rom[36316] = 12'h100;
rom[36317] = 12'h  0;
rom[36318] = 12'h  0;
rom[36319] = 12'h  0;
rom[36320] = 12'h  0;
rom[36321] = 12'h  0;
rom[36322] = 12'h  0;
rom[36323] = 12'h  0;
rom[36324] = 12'h  0;
rom[36325] = 12'h  0;
rom[36326] = 12'h  0;
rom[36327] = 12'h  0;
rom[36328] = 12'h  0;
rom[36329] = 12'h  0;
rom[36330] = 12'h  0;
rom[36331] = 12'h  0;
rom[36332] = 12'h  0;
rom[36333] = 12'h100;
rom[36334] = 12'h100;
rom[36335] = 12'h100;
rom[36336] = 12'h100;
rom[36337] = 12'h100;
rom[36338] = 12'h200;
rom[36339] = 12'h300;
rom[36340] = 12'h300;
rom[36341] = 12'h500;
rom[36342] = 12'h610;
rom[36343] = 12'h710;
rom[36344] = 12'h920;
rom[36345] = 12'ha30;
rom[36346] = 12'hc40;
rom[36347] = 12'hd50;
rom[36348] = 12'he51;
rom[36349] = 12'hf61;
rom[36350] = 12'hf61;
rom[36351] = 12'hf70;
rom[36352] = 12'he81;
rom[36353] = 12'hfa3;
rom[36354] = 12'hfb4;
rom[36355] = 12'hd92;
rom[36356] = 12'ha60;
rom[36357] = 12'h850;
rom[36358] = 12'h740;
rom[36359] = 12'h740;
rom[36360] = 12'h730;
rom[36361] = 12'h730;
rom[36362] = 12'h631;
rom[36363] = 12'h631;
rom[36364] = 12'h631;
rom[36365] = 12'h531;
rom[36366] = 12'h430;
rom[36367] = 12'h420;
rom[36368] = 12'h420;
rom[36369] = 12'h320;
rom[36370] = 12'h320;
rom[36371] = 12'h320;
rom[36372] = 12'h321;
rom[36373] = 12'h221;
rom[36374] = 12'h221;
rom[36375] = 12'h222;
rom[36376] = 12'h322;
rom[36377] = 12'h322;
rom[36378] = 12'h333;
rom[36379] = 12'h333;
rom[36380] = 12'h444;
rom[36381] = 12'h545;
rom[36382] = 12'h556;
rom[36383] = 12'h666;
rom[36384] = 12'h667;
rom[36385] = 12'h777;
rom[36386] = 12'h777;
rom[36387] = 12'h888;
rom[36388] = 12'h888;
rom[36389] = 12'h999;
rom[36390] = 12'h999;
rom[36391] = 12'h999;
rom[36392] = 12'haaa;
rom[36393] = 12'haaa;
rom[36394] = 12'haaa;
rom[36395] = 12'haaa;
rom[36396] = 12'haaa;
rom[36397] = 12'haaa;
rom[36398] = 12'haaa;
rom[36399] = 12'haaa;
rom[36400] = 12'h888;
rom[36401] = 12'h888;
rom[36402] = 12'h888;
rom[36403] = 12'h888;
rom[36404] = 12'h888;
rom[36405] = 12'h888;
rom[36406] = 12'h888;
rom[36407] = 12'h888;
rom[36408] = 12'h888;
rom[36409] = 12'h888;
rom[36410] = 12'h888;
rom[36411] = 12'h888;
rom[36412] = 12'h888;
rom[36413] = 12'h888;
rom[36414] = 12'h888;
rom[36415] = 12'h888;
rom[36416] = 12'h888;
rom[36417] = 12'h888;
rom[36418] = 12'h888;
rom[36419] = 12'h888;
rom[36420] = 12'h999;
rom[36421] = 12'h999;
rom[36422] = 12'h999;
rom[36423] = 12'h999;
rom[36424] = 12'h999;
rom[36425] = 12'h999;
rom[36426] = 12'haaa;
rom[36427] = 12'haaa;
rom[36428] = 12'haaa;
rom[36429] = 12'haaa;
rom[36430] = 12'haaa;
rom[36431] = 12'haaa;
rom[36432] = 12'haaa;
rom[36433] = 12'haaa;
rom[36434] = 12'haaa;
rom[36435] = 12'haaa;
rom[36436] = 12'haaa;
rom[36437] = 12'haaa;
rom[36438] = 12'haaa;
rom[36439] = 12'haaa;
rom[36440] = 12'haaa;
rom[36441] = 12'haaa;
rom[36442] = 12'haaa;
rom[36443] = 12'haaa;
rom[36444] = 12'haaa;
rom[36445] = 12'haaa;
rom[36446] = 12'haaa;
rom[36447] = 12'haaa;
rom[36448] = 12'haaa;
rom[36449] = 12'h999;
rom[36450] = 12'h999;
rom[36451] = 12'h999;
rom[36452] = 12'h999;
rom[36453] = 12'h888;
rom[36454] = 12'h888;
rom[36455] = 12'h888;
rom[36456] = 12'h888;
rom[36457] = 12'h888;
rom[36458] = 12'h888;
rom[36459] = 12'h888;
rom[36460] = 12'h888;
rom[36461] = 12'h888;
rom[36462] = 12'h888;
rom[36463] = 12'h888;
rom[36464] = 12'h777;
rom[36465] = 12'h777;
rom[36466] = 12'h888;
rom[36467] = 12'h888;
rom[36468] = 12'h777;
rom[36469] = 12'h777;
rom[36470] = 12'h777;
rom[36471] = 12'h777;
rom[36472] = 12'h777;
rom[36473] = 12'h777;
rom[36474] = 12'h888;
rom[36475] = 12'h999;
rom[36476] = 12'haaa;
rom[36477] = 12'haaa;
rom[36478] = 12'h999;
rom[36479] = 12'h999;
rom[36480] = 12'h888;
rom[36481] = 12'h777;
rom[36482] = 12'h666;
rom[36483] = 12'h555;
rom[36484] = 12'h555;
rom[36485] = 12'h555;
rom[36486] = 12'h444;
rom[36487] = 12'h444;
rom[36488] = 12'h444;
rom[36489] = 12'h333;
rom[36490] = 12'h333;
rom[36491] = 12'h333;
rom[36492] = 12'h222;
rom[36493] = 12'h222;
rom[36494] = 12'h222;
rom[36495] = 12'h222;
rom[36496] = 12'h222;
rom[36497] = 12'h222;
rom[36498] = 12'h111;
rom[36499] = 12'h111;
rom[36500] = 12'h111;
rom[36501] = 12'h111;
rom[36502] = 12'h  0;
rom[36503] = 12'h  0;
rom[36504] = 12'h  0;
rom[36505] = 12'h  0;
rom[36506] = 12'h  0;
rom[36507] = 12'h  0;
rom[36508] = 12'h  0;
rom[36509] = 12'h  0;
rom[36510] = 12'h  0;
rom[36511] = 12'h  0;
rom[36512] = 12'h  0;
rom[36513] = 12'h  0;
rom[36514] = 12'h  0;
rom[36515] = 12'h  0;
rom[36516] = 12'h  0;
rom[36517] = 12'h  0;
rom[36518] = 12'h  0;
rom[36519] = 12'h  0;
rom[36520] = 12'h  0;
rom[36521] = 12'h  0;
rom[36522] = 12'h  0;
rom[36523] = 12'h  0;
rom[36524] = 12'h  0;
rom[36525] = 12'h  0;
rom[36526] = 12'h  0;
rom[36527] = 12'h  0;
rom[36528] = 12'h  0;
rom[36529] = 12'h  0;
rom[36530] = 12'h  0;
rom[36531] = 12'h  0;
rom[36532] = 12'h  0;
rom[36533] = 12'h  0;
rom[36534] = 12'h  0;
rom[36535] = 12'h  0;
rom[36536] = 12'h  0;
rom[36537] = 12'h  0;
rom[36538] = 12'h  0;
rom[36539] = 12'h  0;
rom[36540] = 12'h  0;
rom[36541] = 12'h  0;
rom[36542] = 12'h  0;
rom[36543] = 12'h  0;
rom[36544] = 12'h  0;
rom[36545] = 12'h  0;
rom[36546] = 12'h  0;
rom[36547] = 12'h  0;
rom[36548] = 12'h  0;
rom[36549] = 12'h  0;
rom[36550] = 12'h  0;
rom[36551] = 12'h  0;
rom[36552] = 12'h  0;
rom[36553] = 12'h  0;
rom[36554] = 12'h  0;
rom[36555] = 12'h  0;
rom[36556] = 12'h  0;
rom[36557] = 12'h  0;
rom[36558] = 12'h  0;
rom[36559] = 12'h  0;
rom[36560] = 12'h  0;
rom[36561] = 12'h  0;
rom[36562] = 12'h  0;
rom[36563] = 12'h  0;
rom[36564] = 12'h  0;
rom[36565] = 12'h  0;
rom[36566] = 12'h  0;
rom[36567] = 12'h  0;
rom[36568] = 12'h  0;
rom[36569] = 12'h  0;
rom[36570] = 12'h  0;
rom[36571] = 12'h  0;
rom[36572] = 12'h  0;
rom[36573] = 12'h  0;
rom[36574] = 12'h  0;
rom[36575] = 12'h  0;
rom[36576] = 12'h  0;
rom[36577] = 12'h  0;
rom[36578] = 12'h  0;
rom[36579] = 12'h  0;
rom[36580] = 12'h  0;
rom[36581] = 12'h  0;
rom[36582] = 12'h  0;
rom[36583] = 12'h  0;
rom[36584] = 12'h  0;
rom[36585] = 12'h  0;
rom[36586] = 12'h  0;
rom[36587] = 12'h  0;
rom[36588] = 12'h  0;
rom[36589] = 12'h  0;
rom[36590] = 12'h  0;
rom[36591] = 12'h  0;
rom[36592] = 12'h  0;
rom[36593] = 12'h  0;
rom[36594] = 12'h111;
rom[36595] = 12'h111;
rom[36596] = 12'h111;
rom[36597] = 12'h222;
rom[36598] = 12'h222;
rom[36599] = 12'h333;
rom[36600] = 12'h444;
rom[36601] = 12'h444;
rom[36602] = 12'h444;
rom[36603] = 12'h444;
rom[36604] = 12'h444;
rom[36605] = 12'h444;
rom[36606] = 12'h444;
rom[36607] = 12'h555;
rom[36608] = 12'h555;
rom[36609] = 12'h555;
rom[36610] = 12'h555;
rom[36611] = 12'h555;
rom[36612] = 12'h555;
rom[36613] = 12'h555;
rom[36614] = 12'h555;
rom[36615] = 12'h444;
rom[36616] = 12'h444;
rom[36617] = 12'h444;
rom[36618] = 12'h444;
rom[36619] = 12'h444;
rom[36620] = 12'h444;
rom[36621] = 12'h444;
rom[36622] = 12'h444;
rom[36623] = 12'h444;
rom[36624] = 12'h444;
rom[36625] = 12'h444;
rom[36626] = 12'h444;
rom[36627] = 12'h444;
rom[36628] = 12'h555;
rom[36629] = 12'h555;
rom[36630] = 12'h555;
rom[36631] = 12'h555;
rom[36632] = 12'h555;
rom[36633] = 12'h555;
rom[36634] = 12'h444;
rom[36635] = 12'h444;
rom[36636] = 12'h333;
rom[36637] = 12'h333;
rom[36638] = 12'h333;
rom[36639] = 12'h333;
rom[36640] = 12'h222;
rom[36641] = 12'h222;
rom[36642] = 12'h222;
rom[36643] = 12'h222;
rom[36644] = 12'h222;
rom[36645] = 12'h222;
rom[36646] = 12'h111;
rom[36647] = 12'h111;
rom[36648] = 12'h111;
rom[36649] = 12'h111;
rom[36650] = 12'h  0;
rom[36651] = 12'h  0;
rom[36652] = 12'h  0;
rom[36653] = 12'h  0;
rom[36654] = 12'h  0;
rom[36655] = 12'h  0;
rom[36656] = 12'h  0;
rom[36657] = 12'h  0;
rom[36658] = 12'h  0;
rom[36659] = 12'h  0;
rom[36660] = 12'h  0;
rom[36661] = 12'h  0;
rom[36662] = 12'h  0;
rom[36663] = 12'h  0;
rom[36664] = 12'h  0;
rom[36665] = 12'h  0;
rom[36666] = 12'h  0;
rom[36667] = 12'h  0;
rom[36668] = 12'h  0;
rom[36669] = 12'h  0;
rom[36670] = 12'h  0;
rom[36671] = 12'h  0;
rom[36672] = 12'h  0;
rom[36673] = 12'h  0;
rom[36674] = 12'h  0;
rom[36675] = 12'h  0;
rom[36676] = 12'h  0;
rom[36677] = 12'h  0;
rom[36678] = 12'h111;
rom[36679] = 12'h111;
rom[36680] = 12'h111;
rom[36681] = 12'h111;
rom[36682] = 12'h111;
rom[36683] = 12'h222;
rom[36684] = 12'h333;
rom[36685] = 12'h333;
rom[36686] = 12'h444;
rom[36687] = 12'h444;
rom[36688] = 12'h333;
rom[36689] = 12'h333;
rom[36690] = 12'h444;
rom[36691] = 12'h555;
rom[36692] = 12'h666;
rom[36693] = 12'h666;
rom[36694] = 12'h777;
rom[36695] = 12'h888;
rom[36696] = 12'h999;
rom[36697] = 12'h999;
rom[36698] = 12'hbba;
rom[36699] = 12'hccb;
rom[36700] = 12'hccb;
rom[36701] = 12'hddc;
rom[36702] = 12'hfee;
rom[36703] = 12'hfed;
rom[36704] = 12'hdb9;
rom[36705] = 12'h753;
rom[36706] = 12'h520;
rom[36707] = 12'h621;
rom[36708] = 12'h621;
rom[36709] = 12'h510;
rom[36710] = 12'h510;
rom[36711] = 12'h510;
rom[36712] = 12'h400;
rom[36713] = 12'h300;
rom[36714] = 12'h200;
rom[36715] = 12'h200;
rom[36716] = 12'h100;
rom[36717] = 12'h  0;
rom[36718] = 12'h  0;
rom[36719] = 12'h  0;
rom[36720] = 12'h  0;
rom[36721] = 12'h  0;
rom[36722] = 12'h  0;
rom[36723] = 12'h  0;
rom[36724] = 12'h  0;
rom[36725] = 12'h  0;
rom[36726] = 12'h  0;
rom[36727] = 12'h  0;
rom[36728] = 12'h  0;
rom[36729] = 12'h  0;
rom[36730] = 12'h  0;
rom[36731] = 12'h  0;
rom[36732] = 12'h  0;
rom[36733] = 12'h100;
rom[36734] = 12'h100;
rom[36735] = 12'h100;
rom[36736] = 12'h200;
rom[36737] = 12'h200;
rom[36738] = 12'h200;
rom[36739] = 12'h300;
rom[36740] = 12'h400;
rom[36741] = 12'h610;
rom[36742] = 12'h710;
rom[36743] = 12'h920;
rom[36744] = 12'ha20;
rom[36745] = 12'hb30;
rom[36746] = 12'hd40;
rom[36747] = 12'hd50;
rom[36748] = 12'he60;
rom[36749] = 12'he60;
rom[36750] = 12'hf60;
rom[36751] = 12'he70;
rom[36752] = 12'hf91;
rom[36753] = 12'hfb3;
rom[36754] = 12'hfb4;
rom[36755] = 12'hc82;
rom[36756] = 12'h950;
rom[36757] = 12'h850;
rom[36758] = 12'h740;
rom[36759] = 12'h630;
rom[36760] = 12'h630;
rom[36761] = 12'h630;
rom[36762] = 12'h631;
rom[36763] = 12'h631;
rom[36764] = 12'h631;
rom[36765] = 12'h531;
rom[36766] = 12'h531;
rom[36767] = 12'h431;
rom[36768] = 12'h431;
rom[36769] = 12'h431;
rom[36770] = 12'h421;
rom[36771] = 12'h321;
rom[36772] = 12'h321;
rom[36773] = 12'h321;
rom[36774] = 12'h321;
rom[36775] = 12'h322;
rom[36776] = 12'h322;
rom[36777] = 12'h322;
rom[36778] = 12'h333;
rom[36779] = 12'h333;
rom[36780] = 12'h444;
rom[36781] = 12'h555;
rom[36782] = 12'h656;
rom[36783] = 12'h666;
rom[36784] = 12'h767;
rom[36785] = 12'h777;
rom[36786] = 12'h777;
rom[36787] = 12'h888;
rom[36788] = 12'h999;
rom[36789] = 12'h999;
rom[36790] = 12'h999;
rom[36791] = 12'h999;
rom[36792] = 12'haaa;
rom[36793] = 12'haaa;
rom[36794] = 12'haaa;
rom[36795] = 12'haaa;
rom[36796] = 12'haaa;
rom[36797] = 12'haaa;
rom[36798] = 12'haaa;
rom[36799] = 12'haaa;
rom[36800] = 12'h888;
rom[36801] = 12'h888;
rom[36802] = 12'h888;
rom[36803] = 12'h888;
rom[36804] = 12'h888;
rom[36805] = 12'h888;
rom[36806] = 12'h888;
rom[36807] = 12'h888;
rom[36808] = 12'h888;
rom[36809] = 12'h888;
rom[36810] = 12'h888;
rom[36811] = 12'h888;
rom[36812] = 12'h888;
rom[36813] = 12'h888;
rom[36814] = 12'h888;
rom[36815] = 12'h888;
rom[36816] = 12'h888;
rom[36817] = 12'h888;
rom[36818] = 12'h888;
rom[36819] = 12'h888;
rom[36820] = 12'h888;
rom[36821] = 12'h999;
rom[36822] = 12'h999;
rom[36823] = 12'h999;
rom[36824] = 12'h999;
rom[36825] = 12'h999;
rom[36826] = 12'h999;
rom[36827] = 12'haaa;
rom[36828] = 12'haaa;
rom[36829] = 12'haaa;
rom[36830] = 12'haaa;
rom[36831] = 12'haaa;
rom[36832] = 12'haaa;
rom[36833] = 12'haaa;
rom[36834] = 12'haaa;
rom[36835] = 12'haaa;
rom[36836] = 12'haaa;
rom[36837] = 12'haaa;
rom[36838] = 12'haaa;
rom[36839] = 12'haaa;
rom[36840] = 12'haaa;
rom[36841] = 12'haaa;
rom[36842] = 12'haaa;
rom[36843] = 12'haaa;
rom[36844] = 12'haaa;
rom[36845] = 12'haaa;
rom[36846] = 12'haaa;
rom[36847] = 12'haaa;
rom[36848] = 12'haaa;
rom[36849] = 12'haaa;
rom[36850] = 12'h999;
rom[36851] = 12'h999;
rom[36852] = 12'h999;
rom[36853] = 12'h999;
rom[36854] = 12'h888;
rom[36855] = 12'h888;
rom[36856] = 12'h888;
rom[36857] = 12'h888;
rom[36858] = 12'h888;
rom[36859] = 12'h888;
rom[36860] = 12'h888;
rom[36861] = 12'h888;
rom[36862] = 12'h888;
rom[36863] = 12'h888;
rom[36864] = 12'h777;
rom[36865] = 12'h777;
rom[36866] = 12'h777;
rom[36867] = 12'h777;
rom[36868] = 12'h777;
rom[36869] = 12'h777;
rom[36870] = 12'h777;
rom[36871] = 12'h777;
rom[36872] = 12'h777;
rom[36873] = 12'h777;
rom[36874] = 12'h777;
rom[36875] = 12'h888;
rom[36876] = 12'h999;
rom[36877] = 12'h999;
rom[36878] = 12'haaa;
rom[36879] = 12'haaa;
rom[36880] = 12'h999;
rom[36881] = 12'h888;
rom[36882] = 12'h777;
rom[36883] = 12'h666;
rom[36884] = 12'h555;
rom[36885] = 12'h555;
rom[36886] = 12'h555;
rom[36887] = 12'h444;
rom[36888] = 12'h444;
rom[36889] = 12'h333;
rom[36890] = 12'h333;
rom[36891] = 12'h333;
rom[36892] = 12'h222;
rom[36893] = 12'h222;
rom[36894] = 12'h222;
rom[36895] = 12'h222;
rom[36896] = 12'h222;
rom[36897] = 12'h222;
rom[36898] = 12'h111;
rom[36899] = 12'h111;
rom[36900] = 12'h111;
rom[36901] = 12'h111;
rom[36902] = 12'h111;
rom[36903] = 12'h  0;
rom[36904] = 12'h  0;
rom[36905] = 12'h  0;
rom[36906] = 12'h  0;
rom[36907] = 12'h  0;
rom[36908] = 12'h  0;
rom[36909] = 12'h  0;
rom[36910] = 12'h  0;
rom[36911] = 12'h  0;
rom[36912] = 12'h  0;
rom[36913] = 12'h  0;
rom[36914] = 12'h  0;
rom[36915] = 12'h  0;
rom[36916] = 12'h  0;
rom[36917] = 12'h  0;
rom[36918] = 12'h  0;
rom[36919] = 12'h  0;
rom[36920] = 12'h  0;
rom[36921] = 12'h  0;
rom[36922] = 12'h  0;
rom[36923] = 12'h  0;
rom[36924] = 12'h  0;
rom[36925] = 12'h  0;
rom[36926] = 12'h  0;
rom[36927] = 12'h  0;
rom[36928] = 12'h  0;
rom[36929] = 12'h  0;
rom[36930] = 12'h  0;
rom[36931] = 12'h  0;
rom[36932] = 12'h  0;
rom[36933] = 12'h  0;
rom[36934] = 12'h  0;
rom[36935] = 12'h  0;
rom[36936] = 12'h  0;
rom[36937] = 12'h  0;
rom[36938] = 12'h  0;
rom[36939] = 12'h  0;
rom[36940] = 12'h  0;
rom[36941] = 12'h  0;
rom[36942] = 12'h  0;
rom[36943] = 12'h  0;
rom[36944] = 12'h  0;
rom[36945] = 12'h  0;
rom[36946] = 12'h  0;
rom[36947] = 12'h  0;
rom[36948] = 12'h  0;
rom[36949] = 12'h  0;
rom[36950] = 12'h  0;
rom[36951] = 12'h  0;
rom[36952] = 12'h  0;
rom[36953] = 12'h  0;
rom[36954] = 12'h  0;
rom[36955] = 12'h  0;
rom[36956] = 12'h  0;
rom[36957] = 12'h  0;
rom[36958] = 12'h  0;
rom[36959] = 12'h  0;
rom[36960] = 12'h  0;
rom[36961] = 12'h  0;
rom[36962] = 12'h  0;
rom[36963] = 12'h  0;
rom[36964] = 12'h  0;
rom[36965] = 12'h  0;
rom[36966] = 12'h  0;
rom[36967] = 12'h  0;
rom[36968] = 12'h  0;
rom[36969] = 12'h  0;
rom[36970] = 12'h  0;
rom[36971] = 12'h  0;
rom[36972] = 12'h  0;
rom[36973] = 12'h  0;
rom[36974] = 12'h  0;
rom[36975] = 12'h  0;
rom[36976] = 12'h  0;
rom[36977] = 12'h  0;
rom[36978] = 12'h  0;
rom[36979] = 12'h  0;
rom[36980] = 12'h  0;
rom[36981] = 12'h  0;
rom[36982] = 12'h  0;
rom[36983] = 12'h  0;
rom[36984] = 12'h  0;
rom[36985] = 12'h  0;
rom[36986] = 12'h  0;
rom[36987] = 12'h  0;
rom[36988] = 12'h  0;
rom[36989] = 12'h  0;
rom[36990] = 12'h  0;
rom[36991] = 12'h  0;
rom[36992] = 12'h  0;
rom[36993] = 12'h  0;
rom[36994] = 12'h111;
rom[36995] = 12'h111;
rom[36996] = 12'h111;
rom[36997] = 12'h222;
rom[36998] = 12'h333;
rom[36999] = 12'h333;
rom[37000] = 12'h444;
rom[37001] = 12'h444;
rom[37002] = 12'h444;
rom[37003] = 12'h444;
rom[37004] = 12'h444;
rom[37005] = 12'h444;
rom[37006] = 12'h444;
rom[37007] = 12'h444;
rom[37008] = 12'h555;
rom[37009] = 12'h555;
rom[37010] = 12'h555;
rom[37011] = 12'h555;
rom[37012] = 12'h444;
rom[37013] = 12'h555;
rom[37014] = 12'h444;
rom[37015] = 12'h444;
rom[37016] = 12'h444;
rom[37017] = 12'h444;
rom[37018] = 12'h444;
rom[37019] = 12'h444;
rom[37020] = 12'h444;
rom[37021] = 12'h444;
rom[37022] = 12'h444;
rom[37023] = 12'h444;
rom[37024] = 12'h444;
rom[37025] = 12'h444;
rom[37026] = 12'h444;
rom[37027] = 12'h444;
rom[37028] = 12'h555;
rom[37029] = 12'h555;
rom[37030] = 12'h555;
rom[37031] = 12'h555;
rom[37032] = 12'h555;
rom[37033] = 12'h444;
rom[37034] = 12'h444;
rom[37035] = 12'h333;
rom[37036] = 12'h333;
rom[37037] = 12'h333;
rom[37038] = 12'h333;
rom[37039] = 12'h222;
rom[37040] = 12'h222;
rom[37041] = 12'h222;
rom[37042] = 12'h222;
rom[37043] = 12'h222;
rom[37044] = 12'h222;
rom[37045] = 12'h222;
rom[37046] = 12'h111;
rom[37047] = 12'h111;
rom[37048] = 12'h111;
rom[37049] = 12'h111;
rom[37050] = 12'h  0;
rom[37051] = 12'h  0;
rom[37052] = 12'h  0;
rom[37053] = 12'h  0;
rom[37054] = 12'h  0;
rom[37055] = 12'h  0;
rom[37056] = 12'h  0;
rom[37057] = 12'h  0;
rom[37058] = 12'h  0;
rom[37059] = 12'h  0;
rom[37060] = 12'h  0;
rom[37061] = 12'h  0;
rom[37062] = 12'h  0;
rom[37063] = 12'h  0;
rom[37064] = 12'h  0;
rom[37065] = 12'h  0;
rom[37066] = 12'h  0;
rom[37067] = 12'h  0;
rom[37068] = 12'h  0;
rom[37069] = 12'h  0;
rom[37070] = 12'h  0;
rom[37071] = 12'h  0;
rom[37072] = 12'h  0;
rom[37073] = 12'h  0;
rom[37074] = 12'h  0;
rom[37075] = 12'h  0;
rom[37076] = 12'h  0;
rom[37077] = 12'h  0;
rom[37078] = 12'h111;
rom[37079] = 12'h111;
rom[37080] = 12'h111;
rom[37081] = 12'h111;
rom[37082] = 12'h111;
rom[37083] = 12'h222;
rom[37084] = 12'h333;
rom[37085] = 12'h444;
rom[37086] = 12'h444;
rom[37087] = 12'h444;
rom[37088] = 12'h433;
rom[37089] = 12'h434;
rom[37090] = 12'h444;
rom[37091] = 12'h555;
rom[37092] = 12'h666;
rom[37093] = 12'h777;
rom[37094] = 12'h788;
rom[37095] = 12'h898;
rom[37096] = 12'h9a9;
rom[37097] = 12'haa9;
rom[37098] = 12'hbbb;
rom[37099] = 12'hccb;
rom[37100] = 12'hddc;
rom[37101] = 12'hffe;
rom[37102] = 12'hffe;
rom[37103] = 12'hdcb;
rom[37104] = 12'h864;
rom[37105] = 12'h621;
rom[37106] = 12'h510;
rom[37107] = 12'h621;
rom[37108] = 12'h620;
rom[37109] = 12'h510;
rom[37110] = 12'h510;
rom[37111] = 12'h500;
rom[37112] = 12'h400;
rom[37113] = 12'h400;
rom[37114] = 12'h300;
rom[37115] = 12'h200;
rom[37116] = 12'h100;
rom[37117] = 12'h  0;
rom[37118] = 12'h  0;
rom[37119] = 12'h  0;
rom[37120] = 12'h  0;
rom[37121] = 12'h  0;
rom[37122] = 12'h  0;
rom[37123] = 12'h  0;
rom[37124] = 12'h  0;
rom[37125] = 12'h  0;
rom[37126] = 12'h  0;
rom[37127] = 12'h  0;
rom[37128] = 12'h  0;
rom[37129] = 12'h  0;
rom[37130] = 12'h  0;
rom[37131] = 12'h  0;
rom[37132] = 12'h100;
rom[37133] = 12'h100;
rom[37134] = 12'h100;
rom[37135] = 12'h200;
rom[37136] = 12'h200;
rom[37137] = 12'h200;
rom[37138] = 12'h300;
rom[37139] = 12'h400;
rom[37140] = 12'h500;
rom[37141] = 12'h710;
rom[37142] = 12'h920;
rom[37143] = 12'ha20;
rom[37144] = 12'hb30;
rom[37145] = 12'hc40;
rom[37146] = 12'hd40;
rom[37147] = 12'he50;
rom[37148] = 12'he60;
rom[37149] = 12'he60;
rom[37150] = 12'he70;
rom[37151] = 12'he70;
rom[37152] = 12'hf92;
rom[37153] = 12'hfb3;
rom[37154] = 12'hea3;
rom[37155] = 12'hb71;
rom[37156] = 12'h850;
rom[37157] = 12'h840;
rom[37158] = 12'h740;
rom[37159] = 12'h630;
rom[37160] = 12'h630;
rom[37161] = 12'h630;
rom[37162] = 12'h631;
rom[37163] = 12'h631;
rom[37164] = 12'h631;
rom[37165] = 12'h531;
rom[37166] = 12'h531;
rom[37167] = 12'h531;
rom[37168] = 12'h531;
rom[37169] = 12'h431;
rom[37170] = 12'h431;
rom[37171] = 12'h431;
rom[37172] = 12'h431;
rom[37173] = 12'h321;
rom[37174] = 12'h322;
rom[37175] = 12'h322;
rom[37176] = 12'h332;
rom[37177] = 12'h333;
rom[37178] = 12'h333;
rom[37179] = 12'h434;
rom[37180] = 12'h444;
rom[37181] = 12'h555;
rom[37182] = 12'h656;
rom[37183] = 12'h666;
rom[37184] = 12'h777;
rom[37185] = 12'h777;
rom[37186] = 12'h888;
rom[37187] = 12'h888;
rom[37188] = 12'h999;
rom[37189] = 12'h999;
rom[37190] = 12'h999;
rom[37191] = 12'haaa;
rom[37192] = 12'haaa;
rom[37193] = 12'haaa;
rom[37194] = 12'haaa;
rom[37195] = 12'haaa;
rom[37196] = 12'haaa;
rom[37197] = 12'haaa;
rom[37198] = 12'haaa;
rom[37199] = 12'haaa;
rom[37200] = 12'h999;
rom[37201] = 12'h999;
rom[37202] = 12'h888;
rom[37203] = 12'h888;
rom[37204] = 12'h888;
rom[37205] = 12'h888;
rom[37206] = 12'h888;
rom[37207] = 12'h888;
rom[37208] = 12'h777;
rom[37209] = 12'h777;
rom[37210] = 12'h777;
rom[37211] = 12'h777;
rom[37212] = 12'h777;
rom[37213] = 12'h777;
rom[37214] = 12'h777;
rom[37215] = 12'h888;
rom[37216] = 12'h888;
rom[37217] = 12'h888;
rom[37218] = 12'h888;
rom[37219] = 12'h888;
rom[37220] = 12'h888;
rom[37221] = 12'h888;
rom[37222] = 12'h888;
rom[37223] = 12'h888;
rom[37224] = 12'h999;
rom[37225] = 12'h999;
rom[37226] = 12'h999;
rom[37227] = 12'h999;
rom[37228] = 12'h999;
rom[37229] = 12'haaa;
rom[37230] = 12'haaa;
rom[37231] = 12'haaa;
rom[37232] = 12'haaa;
rom[37233] = 12'haaa;
rom[37234] = 12'haaa;
rom[37235] = 12'haaa;
rom[37236] = 12'haaa;
rom[37237] = 12'haaa;
rom[37238] = 12'haaa;
rom[37239] = 12'haaa;
rom[37240] = 12'haaa;
rom[37241] = 12'haaa;
rom[37242] = 12'haaa;
rom[37243] = 12'haaa;
rom[37244] = 12'haaa;
rom[37245] = 12'haaa;
rom[37246] = 12'haaa;
rom[37247] = 12'haaa;
rom[37248] = 12'haaa;
rom[37249] = 12'haaa;
rom[37250] = 12'h999;
rom[37251] = 12'h999;
rom[37252] = 12'h999;
rom[37253] = 12'h999;
rom[37254] = 12'h888;
rom[37255] = 12'h888;
rom[37256] = 12'h888;
rom[37257] = 12'h888;
rom[37258] = 12'h888;
rom[37259] = 12'h888;
rom[37260] = 12'h777;
rom[37261] = 12'h777;
rom[37262] = 12'h777;
rom[37263] = 12'h777;
rom[37264] = 12'h888;
rom[37265] = 12'h777;
rom[37266] = 12'h777;
rom[37267] = 12'h777;
rom[37268] = 12'h777;
rom[37269] = 12'h777;
rom[37270] = 12'h777;
rom[37271] = 12'h777;
rom[37272] = 12'h777;
rom[37273] = 12'h777;
rom[37274] = 12'h777;
rom[37275] = 12'h777;
rom[37276] = 12'h888;
rom[37277] = 12'h888;
rom[37278] = 12'h999;
rom[37279] = 12'h999;
rom[37280] = 12'haaa;
rom[37281] = 12'h999;
rom[37282] = 12'h888;
rom[37283] = 12'h777;
rom[37284] = 12'h666;
rom[37285] = 12'h555;
rom[37286] = 12'h555;
rom[37287] = 12'h444;
rom[37288] = 12'h444;
rom[37289] = 12'h333;
rom[37290] = 12'h333;
rom[37291] = 12'h333;
rom[37292] = 12'h333;
rom[37293] = 12'h333;
rom[37294] = 12'h333;
rom[37295] = 12'h333;
rom[37296] = 12'h222;
rom[37297] = 12'h222;
rom[37298] = 12'h111;
rom[37299] = 12'h111;
rom[37300] = 12'h111;
rom[37301] = 12'h111;
rom[37302] = 12'h111;
rom[37303] = 12'h111;
rom[37304] = 12'h111;
rom[37305] = 12'h  0;
rom[37306] = 12'h  0;
rom[37307] = 12'h  0;
rom[37308] = 12'h  0;
rom[37309] = 12'h  0;
rom[37310] = 12'h  0;
rom[37311] = 12'h  0;
rom[37312] = 12'h  0;
rom[37313] = 12'h  0;
rom[37314] = 12'h  0;
rom[37315] = 12'h  0;
rom[37316] = 12'h  0;
rom[37317] = 12'h  0;
rom[37318] = 12'h  0;
rom[37319] = 12'h  0;
rom[37320] = 12'h  0;
rom[37321] = 12'h  0;
rom[37322] = 12'h  0;
rom[37323] = 12'h  0;
rom[37324] = 12'h  0;
rom[37325] = 12'h  0;
rom[37326] = 12'h  0;
rom[37327] = 12'h  0;
rom[37328] = 12'h  0;
rom[37329] = 12'h  0;
rom[37330] = 12'h  0;
rom[37331] = 12'h  0;
rom[37332] = 12'h  0;
rom[37333] = 12'h  0;
rom[37334] = 12'h  0;
rom[37335] = 12'h  0;
rom[37336] = 12'h  0;
rom[37337] = 12'h  0;
rom[37338] = 12'h  0;
rom[37339] = 12'h  0;
rom[37340] = 12'h  0;
rom[37341] = 12'h  0;
rom[37342] = 12'h  0;
rom[37343] = 12'h  0;
rom[37344] = 12'h  0;
rom[37345] = 12'h  0;
rom[37346] = 12'h  0;
rom[37347] = 12'h  0;
rom[37348] = 12'h  0;
rom[37349] = 12'h  0;
rom[37350] = 12'h  0;
rom[37351] = 12'h  0;
rom[37352] = 12'h  0;
rom[37353] = 12'h  0;
rom[37354] = 12'h  0;
rom[37355] = 12'h  0;
rom[37356] = 12'h  0;
rom[37357] = 12'h  0;
rom[37358] = 12'h  0;
rom[37359] = 12'h  0;
rom[37360] = 12'h  0;
rom[37361] = 12'h  0;
rom[37362] = 12'h  0;
rom[37363] = 12'h  0;
rom[37364] = 12'h  0;
rom[37365] = 12'h  0;
rom[37366] = 12'h  0;
rom[37367] = 12'h  0;
rom[37368] = 12'h  0;
rom[37369] = 12'h  0;
rom[37370] = 12'h  0;
rom[37371] = 12'h  0;
rom[37372] = 12'h  0;
rom[37373] = 12'h  0;
rom[37374] = 12'h  0;
rom[37375] = 12'h  0;
rom[37376] = 12'h  0;
rom[37377] = 12'h  0;
rom[37378] = 12'h  0;
rom[37379] = 12'h  0;
rom[37380] = 12'h  0;
rom[37381] = 12'h  0;
rom[37382] = 12'h  0;
rom[37383] = 12'h  0;
rom[37384] = 12'h  0;
rom[37385] = 12'h  0;
rom[37386] = 12'h  0;
rom[37387] = 12'h  0;
rom[37388] = 12'h  0;
rom[37389] = 12'h  0;
rom[37390] = 12'h  0;
rom[37391] = 12'h  0;
rom[37392] = 12'h  0;
rom[37393] = 12'h  0;
rom[37394] = 12'h111;
rom[37395] = 12'h111;
rom[37396] = 12'h222;
rom[37397] = 12'h222;
rom[37398] = 12'h333;
rom[37399] = 12'h333;
rom[37400] = 12'h444;
rom[37401] = 12'h444;
rom[37402] = 12'h444;
rom[37403] = 12'h444;
rom[37404] = 12'h444;
rom[37405] = 12'h444;
rom[37406] = 12'h444;
rom[37407] = 12'h444;
rom[37408] = 12'h444;
rom[37409] = 12'h555;
rom[37410] = 12'h555;
rom[37411] = 12'h444;
rom[37412] = 12'h444;
rom[37413] = 12'h555;
rom[37414] = 12'h444;
rom[37415] = 12'h444;
rom[37416] = 12'h444;
rom[37417] = 12'h444;
rom[37418] = 12'h444;
rom[37419] = 12'h444;
rom[37420] = 12'h444;
rom[37421] = 12'h444;
rom[37422] = 12'h444;
rom[37423] = 12'h444;
rom[37424] = 12'h444;
rom[37425] = 12'h444;
rom[37426] = 12'h444;
rom[37427] = 12'h555;
rom[37428] = 12'h555;
rom[37429] = 12'h555;
rom[37430] = 12'h555;
rom[37431] = 12'h555;
rom[37432] = 12'h444;
rom[37433] = 12'h444;
rom[37434] = 12'h444;
rom[37435] = 12'h333;
rom[37436] = 12'h333;
rom[37437] = 12'h333;
rom[37438] = 12'h333;
rom[37439] = 12'h222;
rom[37440] = 12'h222;
rom[37441] = 12'h222;
rom[37442] = 12'h222;
rom[37443] = 12'h222;
rom[37444] = 12'h222;
rom[37445] = 12'h222;
rom[37446] = 12'h111;
rom[37447] = 12'h111;
rom[37448] = 12'h111;
rom[37449] = 12'h111;
rom[37450] = 12'h  0;
rom[37451] = 12'h  0;
rom[37452] = 12'h  0;
rom[37453] = 12'h  0;
rom[37454] = 12'h  0;
rom[37455] = 12'h  0;
rom[37456] = 12'h  0;
rom[37457] = 12'h  0;
rom[37458] = 12'h  0;
rom[37459] = 12'h  0;
rom[37460] = 12'h  0;
rom[37461] = 12'h  0;
rom[37462] = 12'h  0;
rom[37463] = 12'h  0;
rom[37464] = 12'h  0;
rom[37465] = 12'h  0;
rom[37466] = 12'h  0;
rom[37467] = 12'h  0;
rom[37468] = 12'h  0;
rom[37469] = 12'h  0;
rom[37470] = 12'h  0;
rom[37471] = 12'h  0;
rom[37472] = 12'h  0;
rom[37473] = 12'h  0;
rom[37474] = 12'h  0;
rom[37475] = 12'h  0;
rom[37476] = 12'h  0;
rom[37477] = 12'h111;
rom[37478] = 12'h111;
rom[37479] = 12'h111;
rom[37480] = 12'h111;
rom[37481] = 12'h111;
rom[37482] = 12'h111;
rom[37483] = 12'h222;
rom[37484] = 12'h333;
rom[37485] = 12'h444;
rom[37486] = 12'h444;
rom[37487] = 12'h444;
rom[37488] = 12'h444;
rom[37489] = 12'h444;
rom[37490] = 12'h555;
rom[37491] = 12'h666;
rom[37492] = 12'h666;
rom[37493] = 12'h777;
rom[37494] = 12'h888;
rom[37495] = 12'h999;
rom[37496] = 12'haaa;
rom[37497] = 12'hbba;
rom[37498] = 12'hccb;
rom[37499] = 12'hdcc;
rom[37500] = 12'heed;
rom[37501] = 12'hfff;
rom[37502] = 12'hfed;
rom[37503] = 12'hb98;
rom[37504] = 12'h521;
rom[37505] = 12'h520;
rom[37506] = 12'h520;
rom[37507] = 12'h620;
rom[37508] = 12'h620;
rom[37509] = 12'h610;
rom[37510] = 12'h610;
rom[37511] = 12'h510;
rom[37512] = 12'h500;
rom[37513] = 12'h400;
rom[37514] = 12'h300;
rom[37515] = 12'h200;
rom[37516] = 12'h100;
rom[37517] = 12'h  0;
rom[37518] = 12'h  0;
rom[37519] = 12'h  0;
rom[37520] = 12'h  0;
rom[37521] = 12'h  0;
rom[37522] = 12'h  0;
rom[37523] = 12'h  0;
rom[37524] = 12'h  0;
rom[37525] = 12'h  0;
rom[37526] = 12'h  0;
rom[37527] = 12'h  0;
rom[37528] = 12'h  0;
rom[37529] = 12'h  0;
rom[37530] = 12'h  0;
rom[37531] = 12'h  0;
rom[37532] = 12'h100;
rom[37533] = 12'h100;
rom[37534] = 12'h200;
rom[37535] = 12'h200;
rom[37536] = 12'h200;
rom[37537] = 12'h300;
rom[37538] = 12'h400;
rom[37539] = 12'h500;
rom[37540] = 12'h710;
rom[37541] = 12'h810;
rom[37542] = 12'ha20;
rom[37543] = 12'hb30;
rom[37544] = 12'hc30;
rom[37545] = 12'hd40;
rom[37546] = 12'he50;
rom[37547] = 12'he50;
rom[37548] = 12'he60;
rom[37549] = 12'he60;
rom[37550] = 12'he70;
rom[37551] = 12'he81;
rom[37552] = 12'hfa2;
rom[37553] = 12'hfa3;
rom[37554] = 12'hd92;
rom[37555] = 12'ha60;
rom[37556] = 12'h840;
rom[37557] = 12'h740;
rom[37558] = 12'h740;
rom[37559] = 12'h630;
rom[37560] = 12'h620;
rom[37561] = 12'h620;
rom[37562] = 12'h630;
rom[37563] = 12'h631;
rom[37564] = 12'h631;
rom[37565] = 12'h531;
rom[37566] = 12'h531;
rom[37567] = 12'h531;
rom[37568] = 12'h541;
rom[37569] = 12'h531;
rom[37570] = 12'h531;
rom[37571] = 12'h431;
rom[37572] = 12'h432;
rom[37573] = 12'h432;
rom[37574] = 12'h432;
rom[37575] = 12'h332;
rom[37576] = 12'h333;
rom[37577] = 12'h333;
rom[37578] = 12'h433;
rom[37579] = 12'h444;
rom[37580] = 12'h544;
rom[37581] = 12'h555;
rom[37582] = 12'h666;
rom[37583] = 12'h666;
rom[37584] = 12'h777;
rom[37585] = 12'h777;
rom[37586] = 12'h888;
rom[37587] = 12'h888;
rom[37588] = 12'h999;
rom[37589] = 12'h999;
rom[37590] = 12'haaa;
rom[37591] = 12'haaa;
rom[37592] = 12'haaa;
rom[37593] = 12'haaa;
rom[37594] = 12'haaa;
rom[37595] = 12'haaa;
rom[37596] = 12'haaa;
rom[37597] = 12'haaa;
rom[37598] = 12'haaa;
rom[37599] = 12'haaa;
rom[37600] = 12'h999;
rom[37601] = 12'h999;
rom[37602] = 12'h888;
rom[37603] = 12'h888;
rom[37604] = 12'h888;
rom[37605] = 12'h888;
rom[37606] = 12'h888;
rom[37607] = 12'h888;
rom[37608] = 12'h777;
rom[37609] = 12'h777;
rom[37610] = 12'h777;
rom[37611] = 12'h888;
rom[37612] = 12'h888;
rom[37613] = 12'h888;
rom[37614] = 12'h888;
rom[37615] = 12'h888;
rom[37616] = 12'h888;
rom[37617] = 12'h888;
rom[37618] = 12'h888;
rom[37619] = 12'h888;
rom[37620] = 12'h888;
rom[37621] = 12'h888;
rom[37622] = 12'h888;
rom[37623] = 12'h888;
rom[37624] = 12'h888;
rom[37625] = 12'h888;
rom[37626] = 12'h888;
rom[37627] = 12'h999;
rom[37628] = 12'h999;
rom[37629] = 12'h999;
rom[37630] = 12'h999;
rom[37631] = 12'h999;
rom[37632] = 12'haaa;
rom[37633] = 12'haaa;
rom[37634] = 12'haaa;
rom[37635] = 12'haaa;
rom[37636] = 12'hbbb;
rom[37637] = 12'hbbb;
rom[37638] = 12'hbbb;
rom[37639] = 12'hbbb;
rom[37640] = 12'haaa;
rom[37641] = 12'haaa;
rom[37642] = 12'haaa;
rom[37643] = 12'haaa;
rom[37644] = 12'haaa;
rom[37645] = 12'haaa;
rom[37646] = 12'haaa;
rom[37647] = 12'haaa;
rom[37648] = 12'haaa;
rom[37649] = 12'haaa;
rom[37650] = 12'h999;
rom[37651] = 12'h999;
rom[37652] = 12'h999;
rom[37653] = 12'h999;
rom[37654] = 12'h888;
rom[37655] = 12'h888;
rom[37656] = 12'h888;
rom[37657] = 12'h888;
rom[37658] = 12'h888;
rom[37659] = 12'h888;
rom[37660] = 12'h777;
rom[37661] = 12'h777;
rom[37662] = 12'h777;
rom[37663] = 12'h777;
rom[37664] = 12'h888;
rom[37665] = 12'h777;
rom[37666] = 12'h777;
rom[37667] = 12'h777;
rom[37668] = 12'h777;
rom[37669] = 12'h777;
rom[37670] = 12'h777;
rom[37671] = 12'h777;
rom[37672] = 12'h777;
rom[37673] = 12'h777;
rom[37674] = 12'h777;
rom[37675] = 12'h777;
rom[37676] = 12'h777;
rom[37677] = 12'h888;
rom[37678] = 12'h888;
rom[37679] = 12'h999;
rom[37680] = 12'h999;
rom[37681] = 12'h999;
rom[37682] = 12'h999;
rom[37683] = 12'h888;
rom[37684] = 12'h777;
rom[37685] = 12'h666;
rom[37686] = 12'h666;
rom[37687] = 12'h555;
rom[37688] = 12'h444;
rom[37689] = 12'h444;
rom[37690] = 12'h444;
rom[37691] = 12'h333;
rom[37692] = 12'h333;
rom[37693] = 12'h333;
rom[37694] = 12'h333;
rom[37695] = 12'h333;
rom[37696] = 12'h222;
rom[37697] = 12'h222;
rom[37698] = 12'h111;
rom[37699] = 12'h111;
rom[37700] = 12'h111;
rom[37701] = 12'h111;
rom[37702] = 12'h111;
rom[37703] = 12'h111;
rom[37704] = 12'h111;
rom[37705] = 12'h  0;
rom[37706] = 12'h  0;
rom[37707] = 12'h  0;
rom[37708] = 12'h  0;
rom[37709] = 12'h  0;
rom[37710] = 12'h  0;
rom[37711] = 12'h  0;
rom[37712] = 12'h  0;
rom[37713] = 12'h  0;
rom[37714] = 12'h  0;
rom[37715] = 12'h  0;
rom[37716] = 12'h  0;
rom[37717] = 12'h  0;
rom[37718] = 12'h  0;
rom[37719] = 12'h  0;
rom[37720] = 12'h  0;
rom[37721] = 12'h  0;
rom[37722] = 12'h  0;
rom[37723] = 12'h  0;
rom[37724] = 12'h  0;
rom[37725] = 12'h  0;
rom[37726] = 12'h  0;
rom[37727] = 12'h  0;
rom[37728] = 12'h  0;
rom[37729] = 12'h  0;
rom[37730] = 12'h  0;
rom[37731] = 12'h  0;
rom[37732] = 12'h  0;
rom[37733] = 12'h  0;
rom[37734] = 12'h  0;
rom[37735] = 12'h  0;
rom[37736] = 12'h  0;
rom[37737] = 12'h  0;
rom[37738] = 12'h  0;
rom[37739] = 12'h  0;
rom[37740] = 12'h  0;
rom[37741] = 12'h  0;
rom[37742] = 12'h  0;
rom[37743] = 12'h  0;
rom[37744] = 12'h  0;
rom[37745] = 12'h  0;
rom[37746] = 12'h  0;
rom[37747] = 12'h  0;
rom[37748] = 12'h  0;
rom[37749] = 12'h  0;
rom[37750] = 12'h  0;
rom[37751] = 12'h  0;
rom[37752] = 12'h  0;
rom[37753] = 12'h  0;
rom[37754] = 12'h  0;
rom[37755] = 12'h  0;
rom[37756] = 12'h  0;
rom[37757] = 12'h  0;
rom[37758] = 12'h  0;
rom[37759] = 12'h  0;
rom[37760] = 12'h  0;
rom[37761] = 12'h  0;
rom[37762] = 12'h  0;
rom[37763] = 12'h  0;
rom[37764] = 12'h  0;
rom[37765] = 12'h  0;
rom[37766] = 12'h  0;
rom[37767] = 12'h  0;
rom[37768] = 12'h  0;
rom[37769] = 12'h  0;
rom[37770] = 12'h  0;
rom[37771] = 12'h  0;
rom[37772] = 12'h  0;
rom[37773] = 12'h  0;
rom[37774] = 12'h  0;
rom[37775] = 12'h  0;
rom[37776] = 12'h  0;
rom[37777] = 12'h  0;
rom[37778] = 12'h  0;
rom[37779] = 12'h  0;
rom[37780] = 12'h  0;
rom[37781] = 12'h  0;
rom[37782] = 12'h  0;
rom[37783] = 12'h  0;
rom[37784] = 12'h  0;
rom[37785] = 12'h  0;
rom[37786] = 12'h  0;
rom[37787] = 12'h  0;
rom[37788] = 12'h  0;
rom[37789] = 12'h  0;
rom[37790] = 12'h  0;
rom[37791] = 12'h  0;
rom[37792] = 12'h  0;
rom[37793] = 12'h111;
rom[37794] = 12'h111;
rom[37795] = 12'h111;
rom[37796] = 12'h222;
rom[37797] = 12'h333;
rom[37798] = 12'h333;
rom[37799] = 12'h333;
rom[37800] = 12'h333;
rom[37801] = 12'h444;
rom[37802] = 12'h444;
rom[37803] = 12'h444;
rom[37804] = 12'h444;
rom[37805] = 12'h444;
rom[37806] = 12'h444;
rom[37807] = 12'h444;
rom[37808] = 12'h444;
rom[37809] = 12'h555;
rom[37810] = 12'h555;
rom[37811] = 12'h444;
rom[37812] = 12'h444;
rom[37813] = 12'h555;
rom[37814] = 12'h444;
rom[37815] = 12'h444;
rom[37816] = 12'h444;
rom[37817] = 12'h444;
rom[37818] = 12'h444;
rom[37819] = 12'h444;
rom[37820] = 12'h444;
rom[37821] = 12'h444;
rom[37822] = 12'h444;
rom[37823] = 12'h444;
rom[37824] = 12'h444;
rom[37825] = 12'h444;
rom[37826] = 12'h444;
rom[37827] = 12'h555;
rom[37828] = 12'h555;
rom[37829] = 12'h555;
rom[37830] = 12'h555;
rom[37831] = 12'h555;
rom[37832] = 12'h444;
rom[37833] = 12'h444;
rom[37834] = 12'h444;
rom[37835] = 12'h333;
rom[37836] = 12'h333;
rom[37837] = 12'h333;
rom[37838] = 12'h333;
rom[37839] = 12'h222;
rom[37840] = 12'h222;
rom[37841] = 12'h222;
rom[37842] = 12'h222;
rom[37843] = 12'h222;
rom[37844] = 12'h222;
rom[37845] = 12'h222;
rom[37846] = 12'h111;
rom[37847] = 12'h111;
rom[37848] = 12'h111;
rom[37849] = 12'h111;
rom[37850] = 12'h111;
rom[37851] = 12'h  0;
rom[37852] = 12'h  0;
rom[37853] = 12'h  0;
rom[37854] = 12'h  0;
rom[37855] = 12'h  0;
rom[37856] = 12'h  0;
rom[37857] = 12'h  0;
rom[37858] = 12'h  0;
rom[37859] = 12'h  0;
rom[37860] = 12'h  0;
rom[37861] = 12'h  0;
rom[37862] = 12'h  0;
rom[37863] = 12'h  0;
rom[37864] = 12'h  0;
rom[37865] = 12'h  0;
rom[37866] = 12'h  0;
rom[37867] = 12'h  0;
rom[37868] = 12'h  0;
rom[37869] = 12'h  0;
rom[37870] = 12'h  0;
rom[37871] = 12'h  0;
rom[37872] = 12'h  0;
rom[37873] = 12'h  0;
rom[37874] = 12'h  0;
rom[37875] = 12'h  0;
rom[37876] = 12'h111;
rom[37877] = 12'h111;
rom[37878] = 12'h111;
rom[37879] = 12'h111;
rom[37880] = 12'h222;
rom[37881] = 12'h111;
rom[37882] = 12'h222;
rom[37883] = 12'h222;
rom[37884] = 12'h333;
rom[37885] = 12'h444;
rom[37886] = 12'h444;
rom[37887] = 12'h444;
rom[37888] = 12'h545;
rom[37889] = 12'h555;
rom[37890] = 12'h555;
rom[37891] = 12'h666;
rom[37892] = 12'h777;
rom[37893] = 12'h777;
rom[37894] = 12'h888;
rom[37895] = 12'h999;
rom[37896] = 12'haaa;
rom[37897] = 12'hbba;
rom[37898] = 12'hccb;
rom[37899] = 12'hedc;
rom[37900] = 12'hffe;
rom[37901] = 12'hffe;
rom[37902] = 12'hcba;
rom[37903] = 12'h865;
rom[37904] = 12'h520;
rom[37905] = 12'h620;
rom[37906] = 12'h620;
rom[37907] = 12'h620;
rom[37908] = 12'h721;
rom[37909] = 12'h720;
rom[37910] = 12'h610;
rom[37911] = 12'h610;
rom[37912] = 12'h500;
rom[37913] = 12'h400;
rom[37914] = 12'h300;
rom[37915] = 12'h200;
rom[37916] = 12'h100;
rom[37917] = 12'h100;
rom[37918] = 12'h  0;
rom[37919] = 12'h  0;
rom[37920] = 12'h  0;
rom[37921] = 12'h100;
rom[37922] = 12'h  0;
rom[37923] = 12'h  0;
rom[37924] = 12'h  0;
rom[37925] = 12'h  0;
rom[37926] = 12'h  0;
rom[37927] = 12'h  0;
rom[37928] = 12'h  0;
rom[37929] = 12'h  0;
rom[37930] = 12'h  0;
rom[37931] = 12'h100;
rom[37932] = 12'h100;
rom[37933] = 12'h100;
rom[37934] = 12'h200;
rom[37935] = 12'h200;
rom[37936] = 12'h200;
rom[37937] = 12'h300;
rom[37938] = 12'h400;
rom[37939] = 12'h610;
rom[37940] = 12'h810;
rom[37941] = 12'h920;
rom[37942] = 12'hb30;
rom[37943] = 12'hc30;
rom[37944] = 12'hd40;
rom[37945] = 12'he40;
rom[37946] = 12'he50;
rom[37947] = 12'he50;
rom[37948] = 12'he60;
rom[37949] = 12'he60;
rom[37950] = 12'he70;
rom[37951] = 12'he81;
rom[37952] = 12'hfa2;
rom[37953] = 12'he92;
rom[37954] = 12'hc81;
rom[37955] = 12'h950;
rom[37956] = 12'h840;
rom[37957] = 12'h740;
rom[37958] = 12'h740;
rom[37959] = 12'h620;
rom[37960] = 12'h620;
rom[37961] = 12'h620;
rom[37962] = 12'h620;
rom[37963] = 12'h520;
rom[37964] = 12'h530;
rom[37965] = 12'h531;
rom[37966] = 12'h541;
rom[37967] = 12'h541;
rom[37968] = 12'h541;
rom[37969] = 12'h531;
rom[37970] = 12'h542;
rom[37971] = 12'h532;
rom[37972] = 12'h532;
rom[37973] = 12'h432;
rom[37974] = 12'h432;
rom[37975] = 12'h433;
rom[37976] = 12'h433;
rom[37977] = 12'h443;
rom[37978] = 12'h444;
rom[37979] = 12'h544;
rom[37980] = 12'h555;
rom[37981] = 12'h655;
rom[37982] = 12'h666;
rom[37983] = 12'h666;
rom[37984] = 12'h777;
rom[37985] = 12'h777;
rom[37986] = 12'h888;
rom[37987] = 12'h999;
rom[37988] = 12'h999;
rom[37989] = 12'h999;
rom[37990] = 12'haaa;
rom[37991] = 12'haaa;
rom[37992] = 12'haaa;
rom[37993] = 12'haaa;
rom[37994] = 12'haaa;
rom[37995] = 12'haaa;
rom[37996] = 12'haaa;
rom[37997] = 12'haaa;
rom[37998] = 12'haaa;
rom[37999] = 12'haaa;
rom[38000] = 12'h999;
rom[38001] = 12'h888;
rom[38002] = 12'h888;
rom[38003] = 12'h888;
rom[38004] = 12'h888;
rom[38005] = 12'h888;
rom[38006] = 12'h888;
rom[38007] = 12'h888;
rom[38008] = 12'h888;
rom[38009] = 12'h888;
rom[38010] = 12'h888;
rom[38011] = 12'h888;
rom[38012] = 12'h888;
rom[38013] = 12'h888;
rom[38014] = 12'h999;
rom[38015] = 12'h999;
rom[38016] = 12'h888;
rom[38017] = 12'h888;
rom[38018] = 12'h888;
rom[38019] = 12'h888;
rom[38020] = 12'h888;
rom[38021] = 12'h888;
rom[38022] = 12'h888;
rom[38023] = 12'h888;
rom[38024] = 12'h888;
rom[38025] = 12'h888;
rom[38026] = 12'h888;
rom[38027] = 12'h888;
rom[38028] = 12'h999;
rom[38029] = 12'h999;
rom[38030] = 12'h999;
rom[38031] = 12'h999;
rom[38032] = 12'h999;
rom[38033] = 12'haaa;
rom[38034] = 12'haaa;
rom[38035] = 12'haaa;
rom[38036] = 12'hbbb;
rom[38037] = 12'hbbb;
rom[38038] = 12'hbbb;
rom[38039] = 12'hbbb;
rom[38040] = 12'haaa;
rom[38041] = 12'haaa;
rom[38042] = 12'haaa;
rom[38043] = 12'haaa;
rom[38044] = 12'haaa;
rom[38045] = 12'haaa;
rom[38046] = 12'haaa;
rom[38047] = 12'haaa;
rom[38048] = 12'haaa;
rom[38049] = 12'haaa;
rom[38050] = 12'haaa;
rom[38051] = 12'haaa;
rom[38052] = 12'h999;
rom[38053] = 12'h999;
rom[38054] = 12'h999;
rom[38055] = 12'h999;
rom[38056] = 12'h888;
rom[38057] = 12'h888;
rom[38058] = 12'h888;
rom[38059] = 12'h888;
rom[38060] = 12'h888;
rom[38061] = 12'h888;
rom[38062] = 12'h888;
rom[38063] = 12'h888;
rom[38064] = 12'h888;
rom[38065] = 12'h777;
rom[38066] = 12'h777;
rom[38067] = 12'h777;
rom[38068] = 12'h777;
rom[38069] = 12'h777;
rom[38070] = 12'h777;
rom[38071] = 12'h777;
rom[38072] = 12'h666;
rom[38073] = 12'h666;
rom[38074] = 12'h777;
rom[38075] = 12'h777;
rom[38076] = 12'h777;
rom[38077] = 12'h777;
rom[38078] = 12'h777;
rom[38079] = 12'h888;
rom[38080] = 12'h999;
rom[38081] = 12'h999;
rom[38082] = 12'haaa;
rom[38083] = 12'h999;
rom[38084] = 12'h999;
rom[38085] = 12'h888;
rom[38086] = 12'h777;
rom[38087] = 12'h666;
rom[38088] = 12'h555;
rom[38089] = 12'h555;
rom[38090] = 12'h444;
rom[38091] = 12'h444;
rom[38092] = 12'h333;
rom[38093] = 12'h333;
rom[38094] = 12'h333;
rom[38095] = 12'h222;
rom[38096] = 12'h222;
rom[38097] = 12'h222;
rom[38098] = 12'h222;
rom[38099] = 12'h111;
rom[38100] = 12'h111;
rom[38101] = 12'h111;
rom[38102] = 12'h111;
rom[38103] = 12'h  0;
rom[38104] = 12'h  0;
rom[38105] = 12'h  0;
rom[38106] = 12'h  0;
rom[38107] = 12'h  0;
rom[38108] = 12'h  0;
rom[38109] = 12'h  0;
rom[38110] = 12'h  0;
rom[38111] = 12'h  0;
rom[38112] = 12'h  0;
rom[38113] = 12'h  0;
rom[38114] = 12'h  0;
rom[38115] = 12'h  0;
rom[38116] = 12'h  0;
rom[38117] = 12'h  0;
rom[38118] = 12'h  0;
rom[38119] = 12'h  0;
rom[38120] = 12'h  0;
rom[38121] = 12'h  0;
rom[38122] = 12'h  0;
rom[38123] = 12'h  0;
rom[38124] = 12'h  0;
rom[38125] = 12'h  0;
rom[38126] = 12'h  0;
rom[38127] = 12'h  0;
rom[38128] = 12'h  0;
rom[38129] = 12'h  0;
rom[38130] = 12'h  0;
rom[38131] = 12'h  0;
rom[38132] = 12'h  0;
rom[38133] = 12'h  0;
rom[38134] = 12'h  0;
rom[38135] = 12'h  0;
rom[38136] = 12'h  0;
rom[38137] = 12'h  0;
rom[38138] = 12'h  0;
rom[38139] = 12'h  0;
rom[38140] = 12'h  0;
rom[38141] = 12'h  0;
rom[38142] = 12'h  0;
rom[38143] = 12'h  0;
rom[38144] = 12'h  0;
rom[38145] = 12'h  0;
rom[38146] = 12'h  0;
rom[38147] = 12'h  0;
rom[38148] = 12'h  0;
rom[38149] = 12'h  0;
rom[38150] = 12'h  0;
rom[38151] = 12'h  0;
rom[38152] = 12'h  0;
rom[38153] = 12'h  0;
rom[38154] = 12'h  0;
rom[38155] = 12'h  0;
rom[38156] = 12'h  0;
rom[38157] = 12'h  0;
rom[38158] = 12'h  0;
rom[38159] = 12'h  0;
rom[38160] = 12'h  0;
rom[38161] = 12'h  0;
rom[38162] = 12'h  0;
rom[38163] = 12'h  0;
rom[38164] = 12'h  0;
rom[38165] = 12'h  0;
rom[38166] = 12'h  0;
rom[38167] = 12'h  0;
rom[38168] = 12'h  0;
rom[38169] = 12'h  0;
rom[38170] = 12'h  0;
rom[38171] = 12'h  0;
rom[38172] = 12'h  0;
rom[38173] = 12'h  0;
rom[38174] = 12'h  0;
rom[38175] = 12'h  0;
rom[38176] = 12'h  0;
rom[38177] = 12'h  0;
rom[38178] = 12'h  0;
rom[38179] = 12'h  0;
rom[38180] = 12'h  0;
rom[38181] = 12'h  0;
rom[38182] = 12'h  0;
rom[38183] = 12'h  0;
rom[38184] = 12'h  0;
rom[38185] = 12'h  0;
rom[38186] = 12'h  0;
rom[38187] = 12'h  0;
rom[38188] = 12'h  0;
rom[38189] = 12'h  0;
rom[38190] = 12'h  0;
rom[38191] = 12'h  0;
rom[38192] = 12'h111;
rom[38193] = 12'h111;
rom[38194] = 12'h111;
rom[38195] = 12'h222;
rom[38196] = 12'h222;
rom[38197] = 12'h333;
rom[38198] = 12'h333;
rom[38199] = 12'h333;
rom[38200] = 12'h333;
rom[38201] = 12'h333;
rom[38202] = 12'h444;
rom[38203] = 12'h444;
rom[38204] = 12'h444;
rom[38205] = 12'h444;
rom[38206] = 12'h444;
rom[38207] = 12'h444;
rom[38208] = 12'h444;
rom[38209] = 12'h555;
rom[38210] = 12'h555;
rom[38211] = 12'h444;
rom[38212] = 12'h444;
rom[38213] = 12'h555;
rom[38214] = 12'h444;
rom[38215] = 12'h444;
rom[38216] = 12'h444;
rom[38217] = 12'h444;
rom[38218] = 12'h444;
rom[38219] = 12'h444;
rom[38220] = 12'h555;
rom[38221] = 12'h555;
rom[38222] = 12'h444;
rom[38223] = 12'h444;
rom[38224] = 12'h444;
rom[38225] = 12'h444;
rom[38226] = 12'h444;
rom[38227] = 12'h555;
rom[38228] = 12'h555;
rom[38229] = 12'h555;
rom[38230] = 12'h555;
rom[38231] = 12'h444;
rom[38232] = 12'h444;
rom[38233] = 12'h444;
rom[38234] = 12'h333;
rom[38235] = 12'h333;
rom[38236] = 12'h333;
rom[38237] = 12'h333;
rom[38238] = 12'h333;
rom[38239] = 12'h222;
rom[38240] = 12'h222;
rom[38241] = 12'h222;
rom[38242] = 12'h222;
rom[38243] = 12'h222;
rom[38244] = 12'h222;
rom[38245] = 12'h222;
rom[38246] = 12'h111;
rom[38247] = 12'h111;
rom[38248] = 12'h111;
rom[38249] = 12'h111;
rom[38250] = 12'h111;
rom[38251] = 12'h111;
rom[38252] = 12'h111;
rom[38253] = 12'h  0;
rom[38254] = 12'h  0;
rom[38255] = 12'h  0;
rom[38256] = 12'h  0;
rom[38257] = 12'h  0;
rom[38258] = 12'h  0;
rom[38259] = 12'h  0;
rom[38260] = 12'h  0;
rom[38261] = 12'h  0;
rom[38262] = 12'h  0;
rom[38263] = 12'h  0;
rom[38264] = 12'h  0;
rom[38265] = 12'h  0;
rom[38266] = 12'h  0;
rom[38267] = 12'h  0;
rom[38268] = 12'h  0;
rom[38269] = 12'h  0;
rom[38270] = 12'h  0;
rom[38271] = 12'h  0;
rom[38272] = 12'h  0;
rom[38273] = 12'h  0;
rom[38274] = 12'h111;
rom[38275] = 12'h111;
rom[38276] = 12'h111;
rom[38277] = 12'h111;
rom[38278] = 12'h111;
rom[38279] = 12'h111;
rom[38280] = 12'h222;
rom[38281] = 12'h222;
rom[38282] = 12'h222;
rom[38283] = 12'h333;
rom[38284] = 12'h444;
rom[38285] = 12'h444;
rom[38286] = 12'h444;
rom[38287] = 12'h444;
rom[38288] = 12'h555;
rom[38289] = 12'h555;
rom[38290] = 12'h666;
rom[38291] = 12'h667;
rom[38292] = 12'h777;
rom[38293] = 12'h788;
rom[38294] = 12'h898;
rom[38295] = 12'haa9;
rom[38296] = 12'hbbb;
rom[38297] = 12'hbbb;
rom[38298] = 12'hdcc;
rom[38299] = 12'hfed;
rom[38300] = 12'hffe;
rom[38301] = 12'hfed;
rom[38302] = 12'ha87;
rom[38303] = 12'h532;
rom[38304] = 12'h621;
rom[38305] = 12'h731;
rom[38306] = 12'h620;
rom[38307] = 12'h610;
rom[38308] = 12'h721;
rom[38309] = 12'h720;
rom[38310] = 12'h610;
rom[38311] = 12'h610;
rom[38312] = 12'h500;
rom[38313] = 12'h500;
rom[38314] = 12'h400;
rom[38315] = 12'h300;
rom[38316] = 12'h200;
rom[38317] = 12'h100;
rom[38318] = 12'h  0;
rom[38319] = 12'h  0;
rom[38320] = 12'h  0;
rom[38321] = 12'h  0;
rom[38322] = 12'h  0;
rom[38323] = 12'h  0;
rom[38324] = 12'h  0;
rom[38325] = 12'h  0;
rom[38326] = 12'h  0;
rom[38327] = 12'h  0;
rom[38328] = 12'h  0;
rom[38329] = 12'h  0;
rom[38330] = 12'h100;
rom[38331] = 12'h100;
rom[38332] = 12'h200;
rom[38333] = 12'h200;
rom[38334] = 12'h200;
rom[38335] = 12'h300;
rom[38336] = 12'h300;
rom[38337] = 12'h400;
rom[38338] = 12'h500;
rom[38339] = 12'h710;
rom[38340] = 12'h910;
rom[38341] = 12'hb20;
rom[38342] = 12'hc30;
rom[38343] = 12'hd30;
rom[38344] = 12'he40;
rom[38345] = 12'he40;
rom[38346] = 12'he50;
rom[38347] = 12'he50;
rom[38348] = 12'he60;
rom[38349] = 12'hd60;
rom[38350] = 12'he71;
rom[38351] = 12'he82;
rom[38352] = 12'he93;
rom[38353] = 12'hd92;
rom[38354] = 12'hb71;
rom[38355] = 12'h950;
rom[38356] = 12'h740;
rom[38357] = 12'h740;
rom[38358] = 12'h630;
rom[38359] = 12'h520;
rom[38360] = 12'h630;
rom[38361] = 12'h620;
rom[38362] = 12'h520;
rom[38363] = 12'h520;
rom[38364] = 12'h530;
rom[38365] = 12'h531;
rom[38366] = 12'h541;
rom[38367] = 12'h541;
rom[38368] = 12'h541;
rom[38369] = 12'h542;
rom[38370] = 12'h542;
rom[38371] = 12'h542;
rom[38372] = 12'h542;
rom[38373] = 12'h543;
rom[38374] = 12'h443;
rom[38375] = 12'h443;
rom[38376] = 12'h443;
rom[38377] = 12'h443;
rom[38378] = 12'h444;
rom[38379] = 12'h544;
rom[38380] = 12'h555;
rom[38381] = 12'h655;
rom[38382] = 12'h666;
rom[38383] = 12'h666;
rom[38384] = 12'h777;
rom[38385] = 12'h777;
rom[38386] = 12'h888;
rom[38387] = 12'h999;
rom[38388] = 12'h999;
rom[38389] = 12'h999;
rom[38390] = 12'haaa;
rom[38391] = 12'haaa;
rom[38392] = 12'haaa;
rom[38393] = 12'haaa;
rom[38394] = 12'haaa;
rom[38395] = 12'haaa;
rom[38396] = 12'haaa;
rom[38397] = 12'haaa;
rom[38398] = 12'haaa;
rom[38399] = 12'haaa;
rom[38400] = 12'h888;
rom[38401] = 12'h888;
rom[38402] = 12'h888;
rom[38403] = 12'h888;
rom[38404] = 12'h888;
rom[38405] = 12'h888;
rom[38406] = 12'h888;
rom[38407] = 12'h888;
rom[38408] = 12'h888;
rom[38409] = 12'h888;
rom[38410] = 12'h888;
rom[38411] = 12'h888;
rom[38412] = 12'h888;
rom[38413] = 12'h888;
rom[38414] = 12'h888;
rom[38415] = 12'h888;
rom[38416] = 12'h888;
rom[38417] = 12'h888;
rom[38418] = 12'h888;
rom[38419] = 12'h888;
rom[38420] = 12'h888;
rom[38421] = 12'h888;
rom[38422] = 12'h888;
rom[38423] = 12'h888;
rom[38424] = 12'h888;
rom[38425] = 12'h888;
rom[38426] = 12'h888;
rom[38427] = 12'h888;
rom[38428] = 12'h888;
rom[38429] = 12'h888;
rom[38430] = 12'h999;
rom[38431] = 12'h999;
rom[38432] = 12'h999;
rom[38433] = 12'h999;
rom[38434] = 12'h999;
rom[38435] = 12'haaa;
rom[38436] = 12'haaa;
rom[38437] = 12'haaa;
rom[38438] = 12'hbbb;
rom[38439] = 12'hbbb;
rom[38440] = 12'hbbb;
rom[38441] = 12'hbbb;
rom[38442] = 12'haaa;
rom[38443] = 12'haaa;
rom[38444] = 12'haaa;
rom[38445] = 12'haaa;
rom[38446] = 12'haaa;
rom[38447] = 12'haaa;
rom[38448] = 12'haaa;
rom[38449] = 12'haaa;
rom[38450] = 12'haaa;
rom[38451] = 12'haaa;
rom[38452] = 12'haaa;
rom[38453] = 12'haaa;
rom[38454] = 12'h999;
rom[38455] = 12'h888;
rom[38456] = 12'h888;
rom[38457] = 12'h888;
rom[38458] = 12'h888;
rom[38459] = 12'h888;
rom[38460] = 12'h888;
rom[38461] = 12'h888;
rom[38462] = 12'h888;
rom[38463] = 12'h888;
rom[38464] = 12'h888;
rom[38465] = 12'h777;
rom[38466] = 12'h777;
rom[38467] = 12'h777;
rom[38468] = 12'h777;
rom[38469] = 12'h777;
rom[38470] = 12'h777;
rom[38471] = 12'h777;
rom[38472] = 12'h666;
rom[38473] = 12'h666;
rom[38474] = 12'h666;
rom[38475] = 12'h666;
rom[38476] = 12'h666;
rom[38477] = 12'h777;
rom[38478] = 12'h777;
rom[38479] = 12'h777;
rom[38480] = 12'h888;
rom[38481] = 12'h888;
rom[38482] = 12'h999;
rom[38483] = 12'h999;
rom[38484] = 12'h888;
rom[38485] = 12'h888;
rom[38486] = 12'h777;
rom[38487] = 12'h777;
rom[38488] = 12'h666;
rom[38489] = 12'h666;
rom[38490] = 12'h555;
rom[38491] = 12'h444;
rom[38492] = 12'h444;
rom[38493] = 12'h333;
rom[38494] = 12'h333;
rom[38495] = 12'h333;
rom[38496] = 12'h333;
rom[38497] = 12'h222;
rom[38498] = 12'h222;
rom[38499] = 12'h222;
rom[38500] = 12'h222;
rom[38501] = 12'h222;
rom[38502] = 12'h111;
rom[38503] = 12'h  0;
rom[38504] = 12'h  0;
rom[38505] = 12'h  0;
rom[38506] = 12'h  0;
rom[38507] = 12'h  0;
rom[38508] = 12'h  0;
rom[38509] = 12'h  0;
rom[38510] = 12'h  0;
rom[38511] = 12'h  0;
rom[38512] = 12'h  0;
rom[38513] = 12'h  0;
rom[38514] = 12'h  0;
rom[38515] = 12'h  0;
rom[38516] = 12'h  0;
rom[38517] = 12'h  0;
rom[38518] = 12'h  0;
rom[38519] = 12'h  0;
rom[38520] = 12'h  0;
rom[38521] = 12'h  0;
rom[38522] = 12'h  0;
rom[38523] = 12'h  0;
rom[38524] = 12'h  0;
rom[38525] = 12'h  0;
rom[38526] = 12'h  0;
rom[38527] = 12'h  0;
rom[38528] = 12'h  0;
rom[38529] = 12'h  0;
rom[38530] = 12'h  0;
rom[38531] = 12'h  0;
rom[38532] = 12'h  0;
rom[38533] = 12'h  0;
rom[38534] = 12'h  0;
rom[38535] = 12'h  0;
rom[38536] = 12'h  0;
rom[38537] = 12'h  0;
rom[38538] = 12'h  0;
rom[38539] = 12'h  0;
rom[38540] = 12'h  0;
rom[38541] = 12'h  0;
rom[38542] = 12'h  0;
rom[38543] = 12'h  0;
rom[38544] = 12'h  0;
rom[38545] = 12'h  0;
rom[38546] = 12'h  0;
rom[38547] = 12'h  0;
rom[38548] = 12'h  0;
rom[38549] = 12'h  0;
rom[38550] = 12'h  0;
rom[38551] = 12'h  0;
rom[38552] = 12'h  0;
rom[38553] = 12'h  0;
rom[38554] = 12'h  0;
rom[38555] = 12'h  0;
rom[38556] = 12'h  0;
rom[38557] = 12'h  0;
rom[38558] = 12'h  0;
rom[38559] = 12'h  0;
rom[38560] = 12'h  0;
rom[38561] = 12'h  0;
rom[38562] = 12'h  0;
rom[38563] = 12'h  0;
rom[38564] = 12'h  0;
rom[38565] = 12'h  0;
rom[38566] = 12'h  0;
rom[38567] = 12'h  0;
rom[38568] = 12'h  0;
rom[38569] = 12'h  0;
rom[38570] = 12'h  0;
rom[38571] = 12'h  0;
rom[38572] = 12'h  0;
rom[38573] = 12'h  0;
rom[38574] = 12'h  0;
rom[38575] = 12'h  0;
rom[38576] = 12'h  0;
rom[38577] = 12'h  0;
rom[38578] = 12'h  0;
rom[38579] = 12'h  0;
rom[38580] = 12'h  0;
rom[38581] = 12'h  0;
rom[38582] = 12'h  0;
rom[38583] = 12'h  0;
rom[38584] = 12'h  0;
rom[38585] = 12'h  0;
rom[38586] = 12'h  0;
rom[38587] = 12'h  0;
rom[38588] = 12'h  0;
rom[38589] = 12'h  0;
rom[38590] = 12'h  0;
rom[38591] = 12'h111;
rom[38592] = 12'h111;
rom[38593] = 12'h111;
rom[38594] = 12'h222;
rom[38595] = 12'h222;
rom[38596] = 12'h333;
rom[38597] = 12'h333;
rom[38598] = 12'h333;
rom[38599] = 12'h333;
rom[38600] = 12'h444;
rom[38601] = 12'h444;
rom[38602] = 12'h444;
rom[38603] = 12'h444;
rom[38604] = 12'h444;
rom[38605] = 12'h444;
rom[38606] = 12'h444;
rom[38607] = 12'h444;
rom[38608] = 12'h444;
rom[38609] = 12'h444;
rom[38610] = 12'h444;
rom[38611] = 12'h444;
rom[38612] = 12'h444;
rom[38613] = 12'h555;
rom[38614] = 12'h555;
rom[38615] = 12'h555;
rom[38616] = 12'h555;
rom[38617] = 12'h444;
rom[38618] = 12'h444;
rom[38619] = 12'h444;
rom[38620] = 12'h444;
rom[38621] = 12'h444;
rom[38622] = 12'h444;
rom[38623] = 12'h444;
rom[38624] = 12'h444;
rom[38625] = 12'h444;
rom[38626] = 12'h555;
rom[38627] = 12'h555;
rom[38628] = 12'h444;
rom[38629] = 12'h444;
rom[38630] = 12'h444;
rom[38631] = 12'h444;
rom[38632] = 12'h444;
rom[38633] = 12'h444;
rom[38634] = 12'h333;
rom[38635] = 12'h333;
rom[38636] = 12'h333;
rom[38637] = 12'h333;
rom[38638] = 12'h222;
rom[38639] = 12'h222;
rom[38640] = 12'h222;
rom[38641] = 12'h222;
rom[38642] = 12'h222;
rom[38643] = 12'h222;
rom[38644] = 12'h222;
rom[38645] = 12'h111;
rom[38646] = 12'h111;
rom[38647] = 12'h111;
rom[38648] = 12'h111;
rom[38649] = 12'h111;
rom[38650] = 12'h111;
rom[38651] = 12'h111;
rom[38652] = 12'h111;
rom[38653] = 12'h111;
rom[38654] = 12'h  0;
rom[38655] = 12'h  0;
rom[38656] = 12'h  0;
rom[38657] = 12'h  0;
rom[38658] = 12'h  0;
rom[38659] = 12'h  0;
rom[38660] = 12'h  0;
rom[38661] = 12'h  0;
rom[38662] = 12'h  0;
rom[38663] = 12'h  0;
rom[38664] = 12'h  0;
rom[38665] = 12'h  0;
rom[38666] = 12'h  0;
rom[38667] = 12'h  0;
rom[38668] = 12'h  0;
rom[38669] = 12'h  0;
rom[38670] = 12'h  0;
rom[38671] = 12'h  0;
rom[38672] = 12'h  0;
rom[38673] = 12'h  0;
rom[38674] = 12'h  0;
rom[38675] = 12'h  0;
rom[38676] = 12'h111;
rom[38677] = 12'h111;
rom[38678] = 12'h111;
rom[38679] = 12'h222;
rom[38680] = 12'h222;
rom[38681] = 12'h222;
rom[38682] = 12'h222;
rom[38683] = 12'h333;
rom[38684] = 12'h444;
rom[38685] = 12'h444;
rom[38686] = 12'h444;
rom[38687] = 12'h444;
rom[38688] = 12'h555;
rom[38689] = 12'h555;
rom[38690] = 12'h666;
rom[38691] = 12'h777;
rom[38692] = 12'h888;
rom[38693] = 12'h888;
rom[38694] = 12'h999;
rom[38695] = 12'h9aa;
rom[38696] = 12'hbbb;
rom[38697] = 12'hccc;
rom[38698] = 12'hdcc;
rom[38699] = 12'hfed;
rom[38700] = 12'hfff;
rom[38701] = 12'hca9;
rom[38702] = 12'h543;
rom[38703] = 12'h521;
rom[38704] = 12'h621;
rom[38705] = 12'h620;
rom[38706] = 12'h610;
rom[38707] = 12'h710;
rom[38708] = 12'h720;
rom[38709] = 12'h720;
rom[38710] = 12'h710;
rom[38711] = 12'h710;
rom[38712] = 12'h610;
rom[38713] = 12'h500;
rom[38714] = 12'h500;
rom[38715] = 12'h400;
rom[38716] = 12'h300;
rom[38717] = 12'h200;
rom[38718] = 12'h100;
rom[38719] = 12'h100;
rom[38720] = 12'h  0;
rom[38721] = 12'h  0;
rom[38722] = 12'h  0;
rom[38723] = 12'h  0;
rom[38724] = 12'h  0;
rom[38725] = 12'h  0;
rom[38726] = 12'h  0;
rom[38727] = 12'h  0;
rom[38728] = 12'h100;
rom[38729] = 12'h100;
rom[38730] = 12'h200;
rom[38731] = 12'h200;
rom[38732] = 12'h300;
rom[38733] = 12'h300;
rom[38734] = 12'h400;
rom[38735] = 12'h400;
rom[38736] = 12'h600;
rom[38737] = 12'h710;
rom[38738] = 12'h810;
rom[38739] = 12'h920;
rom[38740] = 12'hb20;
rom[38741] = 12'hc30;
rom[38742] = 12'hd30;
rom[38743] = 12'hd40;
rom[38744] = 12'he40;
rom[38745] = 12'he50;
rom[38746] = 12'he50;
rom[38747] = 12'he50;
rom[38748] = 12'hd50;
rom[38749] = 12'hd60;
rom[38750] = 12'he71;
rom[38751] = 12'he82;
rom[38752] = 12'hd82;
rom[38753] = 12'hb71;
rom[38754] = 12'ha60;
rom[38755] = 12'h840;
rom[38756] = 12'h740;
rom[38757] = 12'h730;
rom[38758] = 12'h630;
rom[38759] = 12'h630;
rom[38760] = 12'h520;
rom[38761] = 12'h520;
rom[38762] = 12'h520;
rom[38763] = 12'h420;
rom[38764] = 12'h520;
rom[38765] = 12'h530;
rom[38766] = 12'h531;
rom[38767] = 12'h531;
rom[38768] = 12'h531;
rom[38769] = 12'h532;
rom[38770] = 12'h542;
rom[38771] = 12'h543;
rom[38772] = 12'h543;
rom[38773] = 12'h543;
rom[38774] = 12'h544;
rom[38775] = 12'h544;
rom[38776] = 12'h544;
rom[38777] = 12'h544;
rom[38778] = 12'h544;
rom[38779] = 12'h544;
rom[38780] = 12'h555;
rom[38781] = 12'h655;
rom[38782] = 12'h766;
rom[38783] = 12'h766;
rom[38784] = 12'h777;
rom[38785] = 12'h888;
rom[38786] = 12'h888;
rom[38787] = 12'h999;
rom[38788] = 12'h999;
rom[38789] = 12'h999;
rom[38790] = 12'h999;
rom[38791] = 12'h999;
rom[38792] = 12'haaa;
rom[38793] = 12'haaa;
rom[38794] = 12'h999;
rom[38795] = 12'haaa;
rom[38796] = 12'haaa;
rom[38797] = 12'haaa;
rom[38798] = 12'haaa;
rom[38799] = 12'haaa;
rom[38800] = 12'h999;
rom[38801] = 12'h999;
rom[38802] = 12'h888;
rom[38803] = 12'h888;
rom[38804] = 12'h888;
rom[38805] = 12'h888;
rom[38806] = 12'h888;
rom[38807] = 12'h888;
rom[38808] = 12'h888;
rom[38809] = 12'h888;
rom[38810] = 12'h888;
rom[38811] = 12'h888;
rom[38812] = 12'h888;
rom[38813] = 12'h888;
rom[38814] = 12'h888;
rom[38815] = 12'h888;
rom[38816] = 12'h888;
rom[38817] = 12'h888;
rom[38818] = 12'h888;
rom[38819] = 12'h888;
rom[38820] = 12'h888;
rom[38821] = 12'h888;
rom[38822] = 12'h888;
rom[38823] = 12'h888;
rom[38824] = 12'h888;
rom[38825] = 12'h888;
rom[38826] = 12'h888;
rom[38827] = 12'h888;
rom[38828] = 12'h888;
rom[38829] = 12'h888;
rom[38830] = 12'h888;
rom[38831] = 12'h888;
rom[38832] = 12'h888;
rom[38833] = 12'h888;
rom[38834] = 12'h999;
rom[38835] = 12'h999;
rom[38836] = 12'haaa;
rom[38837] = 12'haaa;
rom[38838] = 12'haaa;
rom[38839] = 12'hbbb;
rom[38840] = 12'hbbb;
rom[38841] = 12'hbbb;
rom[38842] = 12'hbbb;
rom[38843] = 12'hbbb;
rom[38844] = 12'hbbb;
rom[38845] = 12'hbbb;
rom[38846] = 12'hbbb;
rom[38847] = 12'hbbb;
rom[38848] = 12'haaa;
rom[38849] = 12'haaa;
rom[38850] = 12'haaa;
rom[38851] = 12'haaa;
rom[38852] = 12'haaa;
rom[38853] = 12'haaa;
rom[38854] = 12'h999;
rom[38855] = 12'h999;
rom[38856] = 12'h888;
rom[38857] = 12'h888;
rom[38858] = 12'h888;
rom[38859] = 12'h888;
rom[38860] = 12'h888;
rom[38861] = 12'h888;
rom[38862] = 12'h888;
rom[38863] = 12'h888;
rom[38864] = 12'h888;
rom[38865] = 12'h777;
rom[38866] = 12'h777;
rom[38867] = 12'h777;
rom[38868] = 12'h777;
rom[38869] = 12'h777;
rom[38870] = 12'h777;
rom[38871] = 12'h777;
rom[38872] = 12'h666;
rom[38873] = 12'h666;
rom[38874] = 12'h666;
rom[38875] = 12'h666;
rom[38876] = 12'h666;
rom[38877] = 12'h666;
rom[38878] = 12'h777;
rom[38879] = 12'h777;
rom[38880] = 12'h777;
rom[38881] = 12'h888;
rom[38882] = 12'h999;
rom[38883] = 12'h999;
rom[38884] = 12'h888;
rom[38885] = 12'h888;
rom[38886] = 12'h777;
rom[38887] = 12'h777;
rom[38888] = 12'h666;
rom[38889] = 12'h666;
rom[38890] = 12'h555;
rom[38891] = 12'h555;
rom[38892] = 12'h555;
rom[38893] = 12'h444;
rom[38894] = 12'h444;
rom[38895] = 12'h333;
rom[38896] = 12'h333;
rom[38897] = 12'h333;
rom[38898] = 12'h222;
rom[38899] = 12'h222;
rom[38900] = 12'h222;
rom[38901] = 12'h111;
rom[38902] = 12'h111;
rom[38903] = 12'h111;
rom[38904] = 12'h111;
rom[38905] = 12'h  0;
rom[38906] = 12'h  0;
rom[38907] = 12'h  0;
rom[38908] = 12'h  0;
rom[38909] = 12'h  0;
rom[38910] = 12'h  0;
rom[38911] = 12'h  0;
rom[38912] = 12'h  0;
rom[38913] = 12'h  0;
rom[38914] = 12'h  0;
rom[38915] = 12'h  0;
rom[38916] = 12'h  0;
rom[38917] = 12'h  0;
rom[38918] = 12'h  0;
rom[38919] = 12'h  0;
rom[38920] = 12'h  0;
rom[38921] = 12'h  0;
rom[38922] = 12'h  0;
rom[38923] = 12'h  0;
rom[38924] = 12'h  0;
rom[38925] = 12'h  0;
rom[38926] = 12'h  0;
rom[38927] = 12'h  0;
rom[38928] = 12'h  0;
rom[38929] = 12'h  0;
rom[38930] = 12'h  0;
rom[38931] = 12'h  0;
rom[38932] = 12'h  0;
rom[38933] = 12'h  0;
rom[38934] = 12'h  0;
rom[38935] = 12'h  0;
rom[38936] = 12'h  0;
rom[38937] = 12'h  0;
rom[38938] = 12'h  0;
rom[38939] = 12'h  0;
rom[38940] = 12'h  0;
rom[38941] = 12'h  0;
rom[38942] = 12'h  0;
rom[38943] = 12'h  0;
rom[38944] = 12'h  0;
rom[38945] = 12'h  0;
rom[38946] = 12'h  0;
rom[38947] = 12'h  0;
rom[38948] = 12'h  0;
rom[38949] = 12'h  0;
rom[38950] = 12'h  0;
rom[38951] = 12'h  0;
rom[38952] = 12'h  0;
rom[38953] = 12'h  0;
rom[38954] = 12'h  0;
rom[38955] = 12'h  0;
rom[38956] = 12'h  0;
rom[38957] = 12'h  0;
rom[38958] = 12'h  0;
rom[38959] = 12'h  0;
rom[38960] = 12'h  0;
rom[38961] = 12'h  0;
rom[38962] = 12'h  0;
rom[38963] = 12'h  0;
rom[38964] = 12'h  0;
rom[38965] = 12'h  0;
rom[38966] = 12'h  0;
rom[38967] = 12'h  0;
rom[38968] = 12'h  0;
rom[38969] = 12'h  0;
rom[38970] = 12'h  0;
rom[38971] = 12'h  0;
rom[38972] = 12'h  0;
rom[38973] = 12'h  0;
rom[38974] = 12'h  0;
rom[38975] = 12'h  0;
rom[38976] = 12'h  0;
rom[38977] = 12'h  0;
rom[38978] = 12'h  0;
rom[38979] = 12'h  0;
rom[38980] = 12'h  0;
rom[38981] = 12'h  0;
rom[38982] = 12'h  0;
rom[38983] = 12'h  0;
rom[38984] = 12'h  0;
rom[38985] = 12'h  0;
rom[38986] = 12'h  0;
rom[38987] = 12'h  0;
rom[38988] = 12'h  0;
rom[38989] = 12'h111;
rom[38990] = 12'h111;
rom[38991] = 12'h111;
rom[38992] = 12'h111;
rom[38993] = 12'h222;
rom[38994] = 12'h222;
rom[38995] = 12'h333;
rom[38996] = 12'h333;
rom[38997] = 12'h333;
rom[38998] = 12'h333;
rom[38999] = 12'h333;
rom[39000] = 12'h444;
rom[39001] = 12'h444;
rom[39002] = 12'h444;
rom[39003] = 12'h444;
rom[39004] = 12'h444;
rom[39005] = 12'h444;
rom[39006] = 12'h444;
rom[39007] = 12'h444;
rom[39008] = 12'h444;
rom[39009] = 12'h444;
rom[39010] = 12'h444;
rom[39011] = 12'h444;
rom[39012] = 12'h444;
rom[39013] = 12'h444;
rom[39014] = 12'h444;
rom[39015] = 12'h555;
rom[39016] = 12'h444;
rom[39017] = 12'h444;
rom[39018] = 12'h444;
rom[39019] = 12'h444;
rom[39020] = 12'h444;
rom[39021] = 12'h444;
rom[39022] = 12'h444;
rom[39023] = 12'h444;
rom[39024] = 12'h444;
rom[39025] = 12'h444;
rom[39026] = 12'h444;
rom[39027] = 12'h444;
rom[39028] = 12'h444;
rom[39029] = 12'h444;
rom[39030] = 12'h444;
rom[39031] = 12'h444;
rom[39032] = 12'h444;
rom[39033] = 12'h444;
rom[39034] = 12'h333;
rom[39035] = 12'h333;
rom[39036] = 12'h333;
rom[39037] = 12'h333;
rom[39038] = 12'h222;
rom[39039] = 12'h222;
rom[39040] = 12'h222;
rom[39041] = 12'h222;
rom[39042] = 12'h222;
rom[39043] = 12'h222;
rom[39044] = 12'h111;
rom[39045] = 12'h111;
rom[39046] = 12'h111;
rom[39047] = 12'h111;
rom[39048] = 12'h111;
rom[39049] = 12'h111;
rom[39050] = 12'h111;
rom[39051] = 12'h111;
rom[39052] = 12'h111;
rom[39053] = 12'h111;
rom[39054] = 12'h  0;
rom[39055] = 12'h  0;
rom[39056] = 12'h  0;
rom[39057] = 12'h  0;
rom[39058] = 12'h  0;
rom[39059] = 12'h  0;
rom[39060] = 12'h  0;
rom[39061] = 12'h  0;
rom[39062] = 12'h  0;
rom[39063] = 12'h  0;
rom[39064] = 12'h  0;
rom[39065] = 12'h  0;
rom[39066] = 12'h  0;
rom[39067] = 12'h  0;
rom[39068] = 12'h  0;
rom[39069] = 12'h  0;
rom[39070] = 12'h  0;
rom[39071] = 12'h  0;
rom[39072] = 12'h  0;
rom[39073] = 12'h111;
rom[39074] = 12'h111;
rom[39075] = 12'h111;
rom[39076] = 12'h111;
rom[39077] = 12'h111;
rom[39078] = 12'h111;
rom[39079] = 12'h222;
rom[39080] = 12'h222;
rom[39081] = 12'h222;
rom[39082] = 12'h222;
rom[39083] = 12'h333;
rom[39084] = 12'h444;
rom[39085] = 12'h444;
rom[39086] = 12'h555;
rom[39087] = 12'h444;
rom[39088] = 12'h655;
rom[39089] = 12'h655;
rom[39090] = 12'h666;
rom[39091] = 12'h777;
rom[39092] = 12'h888;
rom[39093] = 12'h899;
rom[39094] = 12'h999;
rom[39095] = 12'haaa;
rom[39096] = 12'hbbb;
rom[39097] = 12'hccc;
rom[39098] = 12'hedd;
rom[39099] = 12'hfee;
rom[39100] = 12'hfed;
rom[39101] = 12'ha97;
rom[39102] = 12'h632;
rom[39103] = 12'h521;
rom[39104] = 12'h621;
rom[39105] = 12'h620;
rom[39106] = 12'h710;
rom[39107] = 12'h710;
rom[39108] = 12'h710;
rom[39109] = 12'h820;
rom[39110] = 12'h810;
rom[39111] = 12'h710;
rom[39112] = 12'h710;
rom[39113] = 12'h610;
rom[39114] = 12'h500;
rom[39115] = 12'h400;
rom[39116] = 12'h300;
rom[39117] = 12'h200;
rom[39118] = 12'h200;
rom[39119] = 12'h100;
rom[39120] = 12'h100;
rom[39121] = 12'h100;
rom[39122] = 12'h  0;
rom[39123] = 12'h  0;
rom[39124] = 12'h  0;
rom[39125] = 12'h  0;
rom[39126] = 12'h100;
rom[39127] = 12'h100;
rom[39128] = 12'h100;
rom[39129] = 12'h200;
rom[39130] = 12'h200;
rom[39131] = 12'h300;
rom[39132] = 12'h400;
rom[39133] = 12'h400;
rom[39134] = 12'h500;
rom[39135] = 12'h600;
rom[39136] = 12'h710;
rom[39137] = 12'h810;
rom[39138] = 12'h920;
rom[39139] = 12'ha20;
rom[39140] = 12'hc30;
rom[39141] = 12'hc30;
rom[39142] = 12'hd30;
rom[39143] = 12'he40;
rom[39144] = 12'he40;
rom[39145] = 12'he40;
rom[39146] = 12'he50;
rom[39147] = 12'hd50;
rom[39148] = 12'hd50;
rom[39149] = 12'hd60;
rom[39150] = 12'he71;
rom[39151] = 12'he82;
rom[39152] = 12'hc71;
rom[39153] = 12'ha61;
rom[39154] = 12'h950;
rom[39155] = 12'h840;
rom[39156] = 12'h740;
rom[39157] = 12'h630;
rom[39158] = 12'h630;
rom[39159] = 12'h530;
rom[39160] = 12'h520;
rom[39161] = 12'h520;
rom[39162] = 12'h420;
rom[39163] = 12'h420;
rom[39164] = 12'h420;
rom[39165] = 12'h430;
rom[39166] = 12'h531;
rom[39167] = 12'h531;
rom[39168] = 12'h532;
rom[39169] = 12'h532;
rom[39170] = 12'h543;
rom[39171] = 12'h543;
rom[39172] = 12'h543;
rom[39173] = 12'h543;
rom[39174] = 12'h544;
rom[39175] = 12'h544;
rom[39176] = 12'h544;
rom[39177] = 12'h544;
rom[39178] = 12'h544;
rom[39179] = 12'h555;
rom[39180] = 12'h555;
rom[39181] = 12'h666;
rom[39182] = 12'h766;
rom[39183] = 12'h777;
rom[39184] = 12'h877;
rom[39185] = 12'h888;
rom[39186] = 12'h999;
rom[39187] = 12'h999;
rom[39188] = 12'h999;
rom[39189] = 12'h999;
rom[39190] = 12'h999;
rom[39191] = 12'h999;
rom[39192] = 12'haaa;
rom[39193] = 12'haaa;
rom[39194] = 12'h999;
rom[39195] = 12'haaa;
rom[39196] = 12'haaa;
rom[39197] = 12'haaa;
rom[39198] = 12'haaa;
rom[39199] = 12'haaa;
rom[39200] = 12'h999;
rom[39201] = 12'h999;
rom[39202] = 12'h999;
rom[39203] = 12'h888;
rom[39204] = 12'h888;
rom[39205] = 12'h888;
rom[39206] = 12'h888;
rom[39207] = 12'h888;
rom[39208] = 12'h888;
rom[39209] = 12'h888;
rom[39210] = 12'h888;
rom[39211] = 12'h777;
rom[39212] = 12'h777;
rom[39213] = 12'h777;
rom[39214] = 12'h777;
rom[39215] = 12'h777;
rom[39216] = 12'h888;
rom[39217] = 12'h888;
rom[39218] = 12'h888;
rom[39219] = 12'h888;
rom[39220] = 12'h888;
rom[39221] = 12'h888;
rom[39222] = 12'h888;
rom[39223] = 12'h888;
rom[39224] = 12'h888;
rom[39225] = 12'h888;
rom[39226] = 12'h888;
rom[39227] = 12'h888;
rom[39228] = 12'h888;
rom[39229] = 12'h888;
rom[39230] = 12'h888;
rom[39231] = 12'h999;
rom[39232] = 12'h999;
rom[39233] = 12'h999;
rom[39234] = 12'h999;
rom[39235] = 12'h999;
rom[39236] = 12'haaa;
rom[39237] = 12'haaa;
rom[39238] = 12'haaa;
rom[39239] = 12'hbbb;
rom[39240] = 12'hbbb;
rom[39241] = 12'hbbb;
rom[39242] = 12'hbbb;
rom[39243] = 12'hbbb;
rom[39244] = 12'hbbb;
rom[39245] = 12'hbbb;
rom[39246] = 12'hbbb;
rom[39247] = 12'hbbb;
rom[39248] = 12'hbbb;
rom[39249] = 12'haaa;
rom[39250] = 12'haaa;
rom[39251] = 12'haaa;
rom[39252] = 12'haaa;
rom[39253] = 12'haaa;
rom[39254] = 12'haaa;
rom[39255] = 12'haaa;
rom[39256] = 12'h999;
rom[39257] = 12'h999;
rom[39258] = 12'h888;
rom[39259] = 12'h888;
rom[39260] = 12'h888;
rom[39261] = 12'h888;
rom[39262] = 12'h888;
rom[39263] = 12'h888;
rom[39264] = 12'h888;
rom[39265] = 12'h888;
rom[39266] = 12'h777;
rom[39267] = 12'h777;
rom[39268] = 12'h777;
rom[39269] = 12'h777;
rom[39270] = 12'h777;
rom[39271] = 12'h777;
rom[39272] = 12'h777;
rom[39273] = 12'h666;
rom[39274] = 12'h666;
rom[39275] = 12'h666;
rom[39276] = 12'h666;
rom[39277] = 12'h666;
rom[39278] = 12'h666;
rom[39279] = 12'h666;
rom[39280] = 12'h777;
rom[39281] = 12'h777;
rom[39282] = 12'h888;
rom[39283] = 12'h888;
rom[39284] = 12'h888;
rom[39285] = 12'h888;
rom[39286] = 12'h888;
rom[39287] = 12'h777;
rom[39288] = 12'h666;
rom[39289] = 12'h666;
rom[39290] = 12'h666;
rom[39291] = 12'h666;
rom[39292] = 12'h555;
rom[39293] = 12'h555;
rom[39294] = 12'h444;
rom[39295] = 12'h444;
rom[39296] = 12'h333;
rom[39297] = 12'h333;
rom[39298] = 12'h333;
rom[39299] = 12'h333;
rom[39300] = 12'h222;
rom[39301] = 12'h111;
rom[39302] = 12'h111;
rom[39303] = 12'h111;
rom[39304] = 12'h111;
rom[39305] = 12'h111;
rom[39306] = 12'h  0;
rom[39307] = 12'h  0;
rom[39308] = 12'h  0;
rom[39309] = 12'h  0;
rom[39310] = 12'h  0;
rom[39311] = 12'h  0;
rom[39312] = 12'h  0;
rom[39313] = 12'h  0;
rom[39314] = 12'h  0;
rom[39315] = 12'h  0;
rom[39316] = 12'h  0;
rom[39317] = 12'h  0;
rom[39318] = 12'h  0;
rom[39319] = 12'h  0;
rom[39320] = 12'h  0;
rom[39321] = 12'h  0;
rom[39322] = 12'h  0;
rom[39323] = 12'h  0;
rom[39324] = 12'h  0;
rom[39325] = 12'h  0;
rom[39326] = 12'h  0;
rom[39327] = 12'h  0;
rom[39328] = 12'h  0;
rom[39329] = 12'h  0;
rom[39330] = 12'h  0;
rom[39331] = 12'h  0;
rom[39332] = 12'h  0;
rom[39333] = 12'h  0;
rom[39334] = 12'h  0;
rom[39335] = 12'h  0;
rom[39336] = 12'h  0;
rom[39337] = 12'h  0;
rom[39338] = 12'h  0;
rom[39339] = 12'h  0;
rom[39340] = 12'h  0;
rom[39341] = 12'h  0;
rom[39342] = 12'h  0;
rom[39343] = 12'h  0;
rom[39344] = 12'h  0;
rom[39345] = 12'h  0;
rom[39346] = 12'h  0;
rom[39347] = 12'h  0;
rom[39348] = 12'h  0;
rom[39349] = 12'h  0;
rom[39350] = 12'h  0;
rom[39351] = 12'h  0;
rom[39352] = 12'h  0;
rom[39353] = 12'h  0;
rom[39354] = 12'h  0;
rom[39355] = 12'h  0;
rom[39356] = 12'h  0;
rom[39357] = 12'h  0;
rom[39358] = 12'h  0;
rom[39359] = 12'h  0;
rom[39360] = 12'h  0;
rom[39361] = 12'h  0;
rom[39362] = 12'h  0;
rom[39363] = 12'h  0;
rom[39364] = 12'h  0;
rom[39365] = 12'h  0;
rom[39366] = 12'h  0;
rom[39367] = 12'h  0;
rom[39368] = 12'h  0;
rom[39369] = 12'h  0;
rom[39370] = 12'h  0;
rom[39371] = 12'h  0;
rom[39372] = 12'h  0;
rom[39373] = 12'h  0;
rom[39374] = 12'h  0;
rom[39375] = 12'h  0;
rom[39376] = 12'h  0;
rom[39377] = 12'h  0;
rom[39378] = 12'h  0;
rom[39379] = 12'h  0;
rom[39380] = 12'h  0;
rom[39381] = 12'h  0;
rom[39382] = 12'h  0;
rom[39383] = 12'h  0;
rom[39384] = 12'h  0;
rom[39385] = 12'h  0;
rom[39386] = 12'h  0;
rom[39387] = 12'h111;
rom[39388] = 12'h111;
rom[39389] = 12'h111;
rom[39390] = 12'h222;
rom[39391] = 12'h222;
rom[39392] = 12'h222;
rom[39393] = 12'h222;
rom[39394] = 12'h222;
rom[39395] = 12'h333;
rom[39396] = 12'h333;
rom[39397] = 12'h333;
rom[39398] = 12'h333;
rom[39399] = 12'h444;
rom[39400] = 12'h444;
rom[39401] = 12'h444;
rom[39402] = 12'h444;
rom[39403] = 12'h444;
rom[39404] = 12'h444;
rom[39405] = 12'h444;
rom[39406] = 12'h444;
rom[39407] = 12'h444;
rom[39408] = 12'h444;
rom[39409] = 12'h444;
rom[39410] = 12'h444;
rom[39411] = 12'h444;
rom[39412] = 12'h444;
rom[39413] = 12'h444;
rom[39414] = 12'h444;
rom[39415] = 12'h444;
rom[39416] = 12'h444;
rom[39417] = 12'h444;
rom[39418] = 12'h444;
rom[39419] = 12'h444;
rom[39420] = 12'h444;
rom[39421] = 12'h444;
rom[39422] = 12'h444;
rom[39423] = 12'h444;
rom[39424] = 12'h444;
rom[39425] = 12'h444;
rom[39426] = 12'h444;
rom[39427] = 12'h444;
rom[39428] = 12'h444;
rom[39429] = 12'h444;
rom[39430] = 12'h444;
rom[39431] = 12'h444;
rom[39432] = 12'h444;
rom[39433] = 12'h444;
rom[39434] = 12'h333;
rom[39435] = 12'h333;
rom[39436] = 12'h333;
rom[39437] = 12'h222;
rom[39438] = 12'h222;
rom[39439] = 12'h222;
rom[39440] = 12'h222;
rom[39441] = 12'h222;
rom[39442] = 12'h222;
rom[39443] = 12'h111;
rom[39444] = 12'h111;
rom[39445] = 12'h111;
rom[39446] = 12'h111;
rom[39447] = 12'h111;
rom[39448] = 12'h111;
rom[39449] = 12'h111;
rom[39450] = 12'h111;
rom[39451] = 12'h111;
rom[39452] = 12'h111;
rom[39453] = 12'h111;
rom[39454] = 12'h  0;
rom[39455] = 12'h  0;
rom[39456] = 12'h  0;
rom[39457] = 12'h  0;
rom[39458] = 12'h  0;
rom[39459] = 12'h  0;
rom[39460] = 12'h  0;
rom[39461] = 12'h  0;
rom[39462] = 12'h  0;
rom[39463] = 12'h  0;
rom[39464] = 12'h  0;
rom[39465] = 12'h  0;
rom[39466] = 12'h  0;
rom[39467] = 12'h  0;
rom[39468] = 12'h  0;
rom[39469] = 12'h  0;
rom[39470] = 12'h  0;
rom[39471] = 12'h  0;
rom[39472] = 12'h111;
rom[39473] = 12'h111;
rom[39474] = 12'h111;
rom[39475] = 12'h111;
rom[39476] = 12'h111;
rom[39477] = 12'h111;
rom[39478] = 12'h111;
rom[39479] = 12'h222;
rom[39480] = 12'h222;
rom[39481] = 12'h222;
rom[39482] = 12'h333;
rom[39483] = 12'h444;
rom[39484] = 12'h444;
rom[39485] = 12'h444;
rom[39486] = 12'h555;
rom[39487] = 12'h555;
rom[39488] = 12'h666;
rom[39489] = 12'h666;
rom[39490] = 12'h767;
rom[39491] = 12'h777;
rom[39492] = 12'h888;
rom[39493] = 12'h999;
rom[39494] = 12'h9aa;
rom[39495] = 12'haba;
rom[39496] = 12'hbbb;
rom[39497] = 12'hdcc;
rom[39498] = 12'hfed;
rom[39499] = 12'hfee;
rom[39500] = 12'hdba;
rom[39501] = 12'h865;
rom[39502] = 12'h532;
rom[39503] = 12'h631;
rom[39504] = 12'h620;
rom[39505] = 12'h620;
rom[39506] = 12'h710;
rom[39507] = 12'h710;
rom[39508] = 12'h720;
rom[39509] = 12'h820;
rom[39510] = 12'h810;
rom[39511] = 12'h810;
rom[39512] = 12'h710;
rom[39513] = 12'h710;
rom[39514] = 12'h610;
rom[39515] = 12'h500;
rom[39516] = 12'h400;
rom[39517] = 12'h300;
rom[39518] = 12'h200;
rom[39519] = 12'h200;
rom[39520] = 12'h200;
rom[39521] = 12'h100;
rom[39522] = 12'h100;
rom[39523] = 12'h100;
rom[39524] = 12'h100;
rom[39525] = 12'h100;
rom[39526] = 12'h200;
rom[39527] = 12'h200;
rom[39528] = 12'h200;
rom[39529] = 12'h300;
rom[39530] = 12'h300;
rom[39531] = 12'h400;
rom[39532] = 12'h500;
rom[39533] = 12'h500;
rom[39534] = 12'h610;
rom[39535] = 12'h710;
rom[39536] = 12'h810;
rom[39537] = 12'h920;
rom[39538] = 12'ha20;
rom[39539] = 12'hb31;
rom[39540] = 12'hc31;
rom[39541] = 12'hd41;
rom[39542] = 12'hd40;
rom[39543] = 12'hd40;
rom[39544] = 12'hd40;
rom[39545] = 12'hd40;
rom[39546] = 12'hd40;
rom[39547] = 12'hd50;
rom[39548] = 12'hd60;
rom[39549] = 12'hd71;
rom[39550] = 12'he71;
rom[39551] = 12'hd82;
rom[39552] = 12'hb61;
rom[39553] = 12'ha60;
rom[39554] = 12'h840;
rom[39555] = 12'h740;
rom[39556] = 12'h730;
rom[39557] = 12'h630;
rom[39558] = 12'h630;
rom[39559] = 12'h520;
rom[39560] = 12'h520;
rom[39561] = 12'h420;
rom[39562] = 12'h420;
rom[39563] = 12'h420;
rom[39564] = 12'h420;
rom[39565] = 12'h420;
rom[39566] = 12'h531;
rom[39567] = 12'h531;
rom[39568] = 12'h532;
rom[39569] = 12'h532;
rom[39570] = 12'h543;
rom[39571] = 12'h543;
rom[39572] = 12'h543;
rom[39573] = 12'h544;
rom[39574] = 12'h544;
rom[39575] = 12'h544;
rom[39576] = 12'h544;
rom[39577] = 12'h544;
rom[39578] = 12'h555;
rom[39579] = 12'h555;
rom[39580] = 12'h655;
rom[39581] = 12'h766;
rom[39582] = 12'h777;
rom[39583] = 12'h777;
rom[39584] = 12'h888;
rom[39585] = 12'h888;
rom[39586] = 12'h999;
rom[39587] = 12'h999;
rom[39588] = 12'haaa;
rom[39589] = 12'haaa;
rom[39590] = 12'haaa;
rom[39591] = 12'haaa;
rom[39592] = 12'haaa;
rom[39593] = 12'haaa;
rom[39594] = 12'h999;
rom[39595] = 12'haaa;
rom[39596] = 12'haaa;
rom[39597] = 12'haaa;
rom[39598] = 12'haaa;
rom[39599] = 12'haaa;
rom[39600] = 12'h999;
rom[39601] = 12'h999;
rom[39602] = 12'h888;
rom[39603] = 12'h888;
rom[39604] = 12'h888;
rom[39605] = 12'h888;
rom[39606] = 12'h888;
rom[39607] = 12'h888;
rom[39608] = 12'h777;
rom[39609] = 12'h777;
rom[39610] = 12'h777;
rom[39611] = 12'h777;
rom[39612] = 12'h777;
rom[39613] = 12'h777;
rom[39614] = 12'h777;
rom[39615] = 12'h888;
rom[39616] = 12'h888;
rom[39617] = 12'h888;
rom[39618] = 12'h888;
rom[39619] = 12'h888;
rom[39620] = 12'h888;
rom[39621] = 12'h888;
rom[39622] = 12'h888;
rom[39623] = 12'h888;
rom[39624] = 12'h888;
rom[39625] = 12'h888;
rom[39626] = 12'h888;
rom[39627] = 12'h999;
rom[39628] = 12'h999;
rom[39629] = 12'h999;
rom[39630] = 12'h999;
rom[39631] = 12'h999;
rom[39632] = 12'h999;
rom[39633] = 12'h999;
rom[39634] = 12'h999;
rom[39635] = 12'h999;
rom[39636] = 12'haaa;
rom[39637] = 12'haaa;
rom[39638] = 12'haaa;
rom[39639] = 12'haaa;
rom[39640] = 12'haaa;
rom[39641] = 12'haaa;
rom[39642] = 12'hbbb;
rom[39643] = 12'hbbb;
rom[39644] = 12'hbbb;
rom[39645] = 12'hbbb;
rom[39646] = 12'hbbb;
rom[39647] = 12'hbbb;
rom[39648] = 12'hbbb;
rom[39649] = 12'hbbb;
rom[39650] = 12'haaa;
rom[39651] = 12'haaa;
rom[39652] = 12'hbbb;
rom[39653] = 12'haaa;
rom[39654] = 12'haaa;
rom[39655] = 12'haaa;
rom[39656] = 12'h999;
rom[39657] = 12'h999;
rom[39658] = 12'h888;
rom[39659] = 12'h888;
rom[39660] = 12'h888;
rom[39661] = 12'h888;
rom[39662] = 12'h888;
rom[39663] = 12'h888;
rom[39664] = 12'h888;
rom[39665] = 12'h888;
rom[39666] = 12'h888;
rom[39667] = 12'h777;
rom[39668] = 12'h777;
rom[39669] = 12'h777;
rom[39670] = 12'h777;
rom[39671] = 12'h777;
rom[39672] = 12'h666;
rom[39673] = 12'h666;
rom[39674] = 12'h666;
rom[39675] = 12'h666;
rom[39676] = 12'h666;
rom[39677] = 12'h666;
rom[39678] = 12'h666;
rom[39679] = 12'h666;
rom[39680] = 12'h666;
rom[39681] = 12'h777;
rom[39682] = 12'h888;
rom[39683] = 12'h888;
rom[39684] = 12'h888;
rom[39685] = 12'h888;
rom[39686] = 12'h888;
rom[39687] = 12'h777;
rom[39688] = 12'h666;
rom[39689] = 12'h666;
rom[39690] = 12'h666;
rom[39691] = 12'h666;
rom[39692] = 12'h666;
rom[39693] = 12'h555;
rom[39694] = 12'h555;
rom[39695] = 12'h555;
rom[39696] = 12'h444;
rom[39697] = 12'h444;
rom[39698] = 12'h444;
rom[39699] = 12'h333;
rom[39700] = 12'h222;
rom[39701] = 12'h111;
rom[39702] = 12'h111;
rom[39703] = 12'h111;
rom[39704] = 12'h111;
rom[39705] = 12'h111;
rom[39706] = 12'h111;
rom[39707] = 12'h  0;
rom[39708] = 12'h  0;
rom[39709] = 12'h  0;
rom[39710] = 12'h  0;
rom[39711] = 12'h  0;
rom[39712] = 12'h  0;
rom[39713] = 12'h  0;
rom[39714] = 12'h  0;
rom[39715] = 12'h  0;
rom[39716] = 12'h  0;
rom[39717] = 12'h  0;
rom[39718] = 12'h  0;
rom[39719] = 12'h  0;
rom[39720] = 12'h  0;
rom[39721] = 12'h  0;
rom[39722] = 12'h  0;
rom[39723] = 12'h  0;
rom[39724] = 12'h  0;
rom[39725] = 12'h  0;
rom[39726] = 12'h  0;
rom[39727] = 12'h  0;
rom[39728] = 12'h  0;
rom[39729] = 12'h  0;
rom[39730] = 12'h  0;
rom[39731] = 12'h  0;
rom[39732] = 12'h  0;
rom[39733] = 12'h  0;
rom[39734] = 12'h  0;
rom[39735] = 12'h  0;
rom[39736] = 12'h  0;
rom[39737] = 12'h  0;
rom[39738] = 12'h  0;
rom[39739] = 12'h  0;
rom[39740] = 12'h  0;
rom[39741] = 12'h  0;
rom[39742] = 12'h  0;
rom[39743] = 12'h  0;
rom[39744] = 12'h  0;
rom[39745] = 12'h  0;
rom[39746] = 12'h  0;
rom[39747] = 12'h  0;
rom[39748] = 12'h  0;
rom[39749] = 12'h  0;
rom[39750] = 12'h  0;
rom[39751] = 12'h  0;
rom[39752] = 12'h  0;
rom[39753] = 12'h  0;
rom[39754] = 12'h  0;
rom[39755] = 12'h  0;
rom[39756] = 12'h  0;
rom[39757] = 12'h  0;
rom[39758] = 12'h  0;
rom[39759] = 12'h  0;
rom[39760] = 12'h  0;
rom[39761] = 12'h  0;
rom[39762] = 12'h  0;
rom[39763] = 12'h  0;
rom[39764] = 12'h  0;
rom[39765] = 12'h  0;
rom[39766] = 12'h  0;
rom[39767] = 12'h  0;
rom[39768] = 12'h  0;
rom[39769] = 12'h  0;
rom[39770] = 12'h  0;
rom[39771] = 12'h  0;
rom[39772] = 12'h  0;
rom[39773] = 12'h  0;
rom[39774] = 12'h  0;
rom[39775] = 12'h  0;
rom[39776] = 12'h  0;
rom[39777] = 12'h  0;
rom[39778] = 12'h  0;
rom[39779] = 12'h  0;
rom[39780] = 12'h  0;
rom[39781] = 12'h  0;
rom[39782] = 12'h  0;
rom[39783] = 12'h  0;
rom[39784] = 12'h111;
rom[39785] = 12'h111;
rom[39786] = 12'h111;
rom[39787] = 12'h111;
rom[39788] = 12'h222;
rom[39789] = 12'h222;
rom[39790] = 12'h222;
rom[39791] = 12'h222;
rom[39792] = 12'h222;
rom[39793] = 12'h222;
rom[39794] = 12'h333;
rom[39795] = 12'h333;
rom[39796] = 12'h333;
rom[39797] = 12'h333;
rom[39798] = 12'h333;
rom[39799] = 12'h333;
rom[39800] = 12'h333;
rom[39801] = 12'h333;
rom[39802] = 12'h444;
rom[39803] = 12'h444;
rom[39804] = 12'h444;
rom[39805] = 12'h444;
rom[39806] = 12'h444;
rom[39807] = 12'h444;
rom[39808] = 12'h444;
rom[39809] = 12'h444;
rom[39810] = 12'h444;
rom[39811] = 12'h444;
rom[39812] = 12'h444;
rom[39813] = 12'h444;
rom[39814] = 12'h444;
rom[39815] = 12'h444;
rom[39816] = 12'h444;
rom[39817] = 12'h444;
rom[39818] = 12'h444;
rom[39819] = 12'h444;
rom[39820] = 12'h444;
rom[39821] = 12'h444;
rom[39822] = 12'h444;
rom[39823] = 12'h444;
rom[39824] = 12'h444;
rom[39825] = 12'h444;
rom[39826] = 12'h444;
rom[39827] = 12'h444;
rom[39828] = 12'h444;
rom[39829] = 12'h444;
rom[39830] = 12'h444;
rom[39831] = 12'h444;
rom[39832] = 12'h444;
rom[39833] = 12'h333;
rom[39834] = 12'h333;
rom[39835] = 12'h333;
rom[39836] = 12'h333;
rom[39837] = 12'h222;
rom[39838] = 12'h222;
rom[39839] = 12'h222;
rom[39840] = 12'h222;
rom[39841] = 12'h222;
rom[39842] = 12'h222;
rom[39843] = 12'h111;
rom[39844] = 12'h111;
rom[39845] = 12'h111;
rom[39846] = 12'h111;
rom[39847] = 12'h111;
rom[39848] = 12'h111;
rom[39849] = 12'h111;
rom[39850] = 12'h111;
rom[39851] = 12'h111;
rom[39852] = 12'h111;
rom[39853] = 12'h  0;
rom[39854] = 12'h  0;
rom[39855] = 12'h  0;
rom[39856] = 12'h  0;
rom[39857] = 12'h  0;
rom[39858] = 12'h  0;
rom[39859] = 12'h  0;
rom[39860] = 12'h  0;
rom[39861] = 12'h  0;
rom[39862] = 12'h  0;
rom[39863] = 12'h  0;
rom[39864] = 12'h  0;
rom[39865] = 12'h  0;
rom[39866] = 12'h  0;
rom[39867] = 12'h  0;
rom[39868] = 12'h  0;
rom[39869] = 12'h  0;
rom[39870] = 12'h  0;
rom[39871] = 12'h  0;
rom[39872] = 12'h  0;
rom[39873] = 12'h111;
rom[39874] = 12'h111;
rom[39875] = 12'h111;
rom[39876] = 12'h111;
rom[39877] = 12'h111;
rom[39878] = 12'h111;
rom[39879] = 12'h111;
rom[39880] = 12'h222;
rom[39881] = 12'h333;
rom[39882] = 12'h333;
rom[39883] = 12'h444;
rom[39884] = 12'h444;
rom[39885] = 12'h444;
rom[39886] = 12'h555;
rom[39887] = 12'h555;
rom[39888] = 12'h666;
rom[39889] = 12'h766;
rom[39890] = 12'h777;
rom[39891] = 12'h888;
rom[39892] = 12'h888;
rom[39893] = 12'h999;
rom[39894] = 12'haaa;
rom[39895] = 12'hbbb;
rom[39896] = 12'hccb;
rom[39897] = 12'hdcc;
rom[39898] = 12'hffe;
rom[39899] = 12'hfed;
rom[39900] = 12'ha88;
rom[39901] = 12'h632;
rom[39902] = 12'h521;
rom[39903] = 12'h621;
rom[39904] = 12'h620;
rom[39905] = 12'h720;
rom[39906] = 12'h720;
rom[39907] = 12'h720;
rom[39908] = 12'h820;
rom[39909] = 12'h820;
rom[39910] = 12'h820;
rom[39911] = 12'h820;
rom[39912] = 12'h810;
rom[39913] = 12'h710;
rom[39914] = 12'h710;
rom[39915] = 12'h610;
rom[39916] = 12'h500;
rom[39917] = 12'h400;
rom[39918] = 12'h300;
rom[39919] = 12'h300;
rom[39920] = 12'h300;
rom[39921] = 12'h200;
rom[39922] = 12'h200;
rom[39923] = 12'h200;
rom[39924] = 12'h200;
rom[39925] = 12'h200;
rom[39926] = 12'h300;
rom[39927] = 12'h300;
rom[39928] = 12'h300;
rom[39929] = 12'h400;
rom[39930] = 12'h400;
rom[39931] = 12'h500;
rom[39932] = 12'h600;
rom[39933] = 12'h710;
rom[39934] = 12'h710;
rom[39935] = 12'h820;
rom[39936] = 12'h920;
rom[39937] = 12'ha30;
rom[39938] = 12'hb31;
rom[39939] = 12'hc41;
rom[39940] = 12'hd41;
rom[39941] = 12'hd41;
rom[39942] = 12'hd40;
rom[39943] = 12'hd40;
rom[39944] = 12'hd40;
rom[39945] = 12'hd40;
rom[39946] = 12'hc40;
rom[39947] = 12'hd50;
rom[39948] = 12'hd61;
rom[39949] = 12'hd71;
rom[39950] = 12'hd71;
rom[39951] = 12'hc71;
rom[39952] = 12'ha50;
rom[39953] = 12'h950;
rom[39954] = 12'h840;
rom[39955] = 12'h730;
rom[39956] = 12'h630;
rom[39957] = 12'h630;
rom[39958] = 12'h530;
rom[39959] = 12'h520;
rom[39960] = 12'h520;
rom[39961] = 12'h420;
rom[39962] = 12'h420;
rom[39963] = 12'h420;
rom[39964] = 12'h420;
rom[39965] = 12'h430;
rom[39966] = 12'h531;
rom[39967] = 12'h531;
rom[39968] = 12'h532;
rom[39969] = 12'h532;
rom[39970] = 12'h543;
rom[39971] = 12'h543;
rom[39972] = 12'h543;
rom[39973] = 12'h544;
rom[39974] = 12'h544;
rom[39975] = 12'h554;
rom[39976] = 12'h544;
rom[39977] = 12'h555;
rom[39978] = 12'h555;
rom[39979] = 12'h655;
rom[39980] = 12'h666;
rom[39981] = 12'h766;
rom[39982] = 12'h877;
rom[39983] = 12'h877;
rom[39984] = 12'h888;
rom[39985] = 12'h999;
rom[39986] = 12'h999;
rom[39987] = 12'haaa;
rom[39988] = 12'haaa;
rom[39989] = 12'haaa;
rom[39990] = 12'haaa;
rom[39991] = 12'haaa;
rom[39992] = 12'haaa;
rom[39993] = 12'haaa;
rom[39994] = 12'h999;
rom[39995] = 12'haaa;
rom[39996] = 12'haaa;
rom[39997] = 12'haaa;
rom[39998] = 12'haaa;
rom[39999] = 12'haaa;
rom[40000] = 12'h999;
rom[40001] = 12'h888;
rom[40002] = 12'h888;
rom[40003] = 12'h888;
rom[40004] = 12'h888;
rom[40005] = 12'h888;
rom[40006] = 12'h888;
rom[40007] = 12'h888;
rom[40008] = 12'h777;
rom[40009] = 12'h777;
rom[40010] = 12'h777;
rom[40011] = 12'h777;
rom[40012] = 12'h777;
rom[40013] = 12'h777;
rom[40014] = 12'h888;
rom[40015] = 12'h888;
rom[40016] = 12'h888;
rom[40017] = 12'h888;
rom[40018] = 12'h888;
rom[40019] = 12'h888;
rom[40020] = 12'h888;
rom[40021] = 12'h888;
rom[40022] = 12'h888;
rom[40023] = 12'h888;
rom[40024] = 12'h888;
rom[40025] = 12'h888;
rom[40026] = 12'h999;
rom[40027] = 12'h999;
rom[40028] = 12'h999;
rom[40029] = 12'h999;
rom[40030] = 12'h999;
rom[40031] = 12'h999;
rom[40032] = 12'h999;
rom[40033] = 12'h999;
rom[40034] = 12'h999;
rom[40035] = 12'h999;
rom[40036] = 12'h999;
rom[40037] = 12'h999;
rom[40038] = 12'h999;
rom[40039] = 12'haaa;
rom[40040] = 12'haaa;
rom[40041] = 12'haaa;
rom[40042] = 12'haaa;
rom[40043] = 12'hbbb;
rom[40044] = 12'hbbb;
rom[40045] = 12'hbbb;
rom[40046] = 12'hbbb;
rom[40047] = 12'hbbb;
rom[40048] = 12'hbbb;
rom[40049] = 12'hbbb;
rom[40050] = 12'hbbb;
rom[40051] = 12'hbbb;
rom[40052] = 12'hbbb;
rom[40053] = 12'haaa;
rom[40054] = 12'haaa;
rom[40055] = 12'haaa;
rom[40056] = 12'haaa;
rom[40057] = 12'h999;
rom[40058] = 12'h999;
rom[40059] = 12'h888;
rom[40060] = 12'h888;
rom[40061] = 12'h888;
rom[40062] = 12'h888;
rom[40063] = 12'h888;
rom[40064] = 12'h888;
rom[40065] = 12'h888;
rom[40066] = 12'h888;
rom[40067] = 12'h777;
rom[40068] = 12'h777;
rom[40069] = 12'h777;
rom[40070] = 12'h777;
rom[40071] = 12'h777;
rom[40072] = 12'h666;
rom[40073] = 12'h666;
rom[40074] = 12'h666;
rom[40075] = 12'h666;
rom[40076] = 12'h666;
rom[40077] = 12'h666;
rom[40078] = 12'h666;
rom[40079] = 12'h666;
rom[40080] = 12'h666;
rom[40081] = 12'h666;
rom[40082] = 12'h777;
rom[40083] = 12'h777;
rom[40084] = 12'h888;
rom[40085] = 12'h888;
rom[40086] = 12'h888;
rom[40087] = 12'h888;
rom[40088] = 12'h777;
rom[40089] = 12'h666;
rom[40090] = 12'h666;
rom[40091] = 12'h555;
rom[40092] = 12'h555;
rom[40093] = 12'h555;
rom[40094] = 12'h555;
rom[40095] = 12'h555;
rom[40096] = 12'h444;
rom[40097] = 12'h444;
rom[40098] = 12'h444;
rom[40099] = 12'h444;
rom[40100] = 12'h333;
rom[40101] = 12'h222;
rom[40102] = 12'h222;
rom[40103] = 12'h222;
rom[40104] = 12'h111;
rom[40105] = 12'h111;
rom[40106] = 12'h111;
rom[40107] = 12'h111;
rom[40108] = 12'h111;
rom[40109] = 12'h  0;
rom[40110] = 12'h  0;
rom[40111] = 12'h  0;
rom[40112] = 12'h  0;
rom[40113] = 12'h  0;
rom[40114] = 12'h  0;
rom[40115] = 12'h  0;
rom[40116] = 12'h  0;
rom[40117] = 12'h  0;
rom[40118] = 12'h  0;
rom[40119] = 12'h  0;
rom[40120] = 12'h  0;
rom[40121] = 12'h  0;
rom[40122] = 12'h  0;
rom[40123] = 12'h  0;
rom[40124] = 12'h  0;
rom[40125] = 12'h  0;
rom[40126] = 12'h  0;
rom[40127] = 12'h  0;
rom[40128] = 12'h  0;
rom[40129] = 12'h  0;
rom[40130] = 12'h  0;
rom[40131] = 12'h  0;
rom[40132] = 12'h  0;
rom[40133] = 12'h  0;
rom[40134] = 12'h  0;
rom[40135] = 12'h  0;
rom[40136] = 12'h  0;
rom[40137] = 12'h  0;
rom[40138] = 12'h  0;
rom[40139] = 12'h  0;
rom[40140] = 12'h  0;
rom[40141] = 12'h  0;
rom[40142] = 12'h  0;
rom[40143] = 12'h  0;
rom[40144] = 12'h  0;
rom[40145] = 12'h  0;
rom[40146] = 12'h  0;
rom[40147] = 12'h  0;
rom[40148] = 12'h  0;
rom[40149] = 12'h  0;
rom[40150] = 12'h  0;
rom[40151] = 12'h  0;
rom[40152] = 12'h  0;
rom[40153] = 12'h  0;
rom[40154] = 12'h  0;
rom[40155] = 12'h  0;
rom[40156] = 12'h  0;
rom[40157] = 12'h  0;
rom[40158] = 12'h  0;
rom[40159] = 12'h  0;
rom[40160] = 12'h  0;
rom[40161] = 12'h  0;
rom[40162] = 12'h  0;
rom[40163] = 12'h  0;
rom[40164] = 12'h  0;
rom[40165] = 12'h  0;
rom[40166] = 12'h  0;
rom[40167] = 12'h  0;
rom[40168] = 12'h  0;
rom[40169] = 12'h  0;
rom[40170] = 12'h  0;
rom[40171] = 12'h  0;
rom[40172] = 12'h  0;
rom[40173] = 12'h  0;
rom[40174] = 12'h  0;
rom[40175] = 12'h  0;
rom[40176] = 12'h  0;
rom[40177] = 12'h  0;
rom[40178] = 12'h  0;
rom[40179] = 12'h  0;
rom[40180] = 12'h  0;
rom[40181] = 12'h  0;
rom[40182] = 12'h111;
rom[40183] = 12'h111;
rom[40184] = 12'h111;
rom[40185] = 12'h111;
rom[40186] = 12'h111;
rom[40187] = 12'h222;
rom[40188] = 12'h222;
rom[40189] = 12'h222;
rom[40190] = 12'h222;
rom[40191] = 12'h222;
rom[40192] = 12'h333;
rom[40193] = 12'h333;
rom[40194] = 12'h333;
rom[40195] = 12'h333;
rom[40196] = 12'h333;
rom[40197] = 12'h333;
rom[40198] = 12'h333;
rom[40199] = 12'h333;
rom[40200] = 12'h333;
rom[40201] = 12'h333;
rom[40202] = 12'h444;
rom[40203] = 12'h444;
rom[40204] = 12'h444;
rom[40205] = 12'h444;
rom[40206] = 12'h444;
rom[40207] = 12'h444;
rom[40208] = 12'h444;
rom[40209] = 12'h444;
rom[40210] = 12'h444;
rom[40211] = 12'h444;
rom[40212] = 12'h444;
rom[40213] = 12'h444;
rom[40214] = 12'h444;
rom[40215] = 12'h444;
rom[40216] = 12'h444;
rom[40217] = 12'h444;
rom[40218] = 12'h444;
rom[40219] = 12'h444;
rom[40220] = 12'h444;
rom[40221] = 12'h444;
rom[40222] = 12'h444;
rom[40223] = 12'h333;
rom[40224] = 12'h444;
rom[40225] = 12'h444;
rom[40226] = 12'h444;
rom[40227] = 12'h444;
rom[40228] = 12'h444;
rom[40229] = 12'h444;
rom[40230] = 12'h444;
rom[40231] = 12'h444;
rom[40232] = 12'h444;
rom[40233] = 12'h333;
rom[40234] = 12'h333;
rom[40235] = 12'h333;
rom[40236] = 12'h222;
rom[40237] = 12'h222;
rom[40238] = 12'h222;
rom[40239] = 12'h222;
rom[40240] = 12'h222;
rom[40241] = 12'h222;
rom[40242] = 12'h111;
rom[40243] = 12'h111;
rom[40244] = 12'h111;
rom[40245] = 12'h111;
rom[40246] = 12'h111;
rom[40247] = 12'h111;
rom[40248] = 12'h111;
rom[40249] = 12'h111;
rom[40250] = 12'h111;
rom[40251] = 12'h111;
rom[40252] = 12'h111;
rom[40253] = 12'h  0;
rom[40254] = 12'h  0;
rom[40255] = 12'h  0;
rom[40256] = 12'h  0;
rom[40257] = 12'h  0;
rom[40258] = 12'h  0;
rom[40259] = 12'h  0;
rom[40260] = 12'h  0;
rom[40261] = 12'h  0;
rom[40262] = 12'h  0;
rom[40263] = 12'h  0;
rom[40264] = 12'h  0;
rom[40265] = 12'h  0;
rom[40266] = 12'h  0;
rom[40267] = 12'h  0;
rom[40268] = 12'h  0;
rom[40269] = 12'h  0;
rom[40270] = 12'h  0;
rom[40271] = 12'h  0;
rom[40272] = 12'h  0;
rom[40273] = 12'h111;
rom[40274] = 12'h111;
rom[40275] = 12'h111;
rom[40276] = 12'h111;
rom[40277] = 12'h111;
rom[40278] = 12'h111;
rom[40279] = 12'h111;
rom[40280] = 12'h222;
rom[40281] = 12'h333;
rom[40282] = 12'h444;
rom[40283] = 12'h444;
rom[40284] = 12'h444;
rom[40285] = 12'h444;
rom[40286] = 12'h555;
rom[40287] = 12'h655;
rom[40288] = 12'h666;
rom[40289] = 12'h777;
rom[40290] = 12'h888;
rom[40291] = 12'h888;
rom[40292] = 12'h899;
rom[40293] = 12'h999;
rom[40294] = 12'haaa;
rom[40295] = 12'hbbb;
rom[40296] = 12'hccc;
rom[40297] = 12'hedd;
rom[40298] = 12'hfff;
rom[40299] = 12'hfdc;
rom[40300] = 12'h966;
rom[40301] = 12'h521;
rom[40302] = 12'h521;
rom[40303] = 12'h621;
rom[40304] = 12'h610;
rom[40305] = 12'h720;
rom[40306] = 12'h720;
rom[40307] = 12'h820;
rom[40308] = 12'h820;
rom[40309] = 12'h820;
rom[40310] = 12'h920;
rom[40311] = 12'h920;
rom[40312] = 12'h820;
rom[40313] = 12'h820;
rom[40314] = 12'h710;
rom[40315] = 12'h710;
rom[40316] = 12'h610;
rom[40317] = 12'h500;
rom[40318] = 12'h500;
rom[40319] = 12'h400;
rom[40320] = 12'h400;
rom[40321] = 12'h400;
rom[40322] = 12'h400;
rom[40323] = 12'h300;
rom[40324] = 12'h300;
rom[40325] = 12'h400;
rom[40326] = 12'h400;
rom[40327] = 12'h400;
rom[40328] = 12'h500;
rom[40329] = 12'h500;
rom[40330] = 12'h600;
rom[40331] = 12'h610;
rom[40332] = 12'h710;
rom[40333] = 12'h820;
rom[40334] = 12'h920;
rom[40335] = 12'h920;
rom[40336] = 12'ha31;
rom[40337] = 12'hb31;
rom[40338] = 12'hc41;
rom[40339] = 12'hc41;
rom[40340] = 12'hd41;
rom[40341] = 12'hd41;
rom[40342] = 12'hd30;
rom[40343] = 12'hd30;
rom[40344] = 12'hc30;
rom[40345] = 12'hc30;
rom[40346] = 12'hc40;
rom[40347] = 12'hc50;
rom[40348] = 12'hd61;
rom[40349] = 12'hd72;
rom[40350] = 12'hc71;
rom[40351] = 12'hb61;
rom[40352] = 12'h950;
rom[40353] = 12'h840;
rom[40354] = 12'h730;
rom[40355] = 12'h730;
rom[40356] = 12'h630;
rom[40357] = 12'h630;
rom[40358] = 12'h630;
rom[40359] = 12'h520;
rom[40360] = 12'h520;
rom[40361] = 12'h420;
rom[40362] = 12'h420;
rom[40363] = 12'h420;
rom[40364] = 12'h420;
rom[40365] = 12'h430;
rom[40366] = 12'h531;
rom[40367] = 12'h531;
rom[40368] = 12'h532;
rom[40369] = 12'h532;
rom[40370] = 12'h543;
rom[40371] = 12'h543;
rom[40372] = 12'h543;
rom[40373] = 12'h544;
rom[40374] = 12'h554;
rom[40375] = 12'h554;
rom[40376] = 12'h555;
rom[40377] = 12'h555;
rom[40378] = 12'h555;
rom[40379] = 12'h666;
rom[40380] = 12'h666;
rom[40381] = 12'h777;
rom[40382] = 12'h877;
rom[40383] = 12'h888;
rom[40384] = 12'h988;
rom[40385] = 12'h999;
rom[40386] = 12'h999;
rom[40387] = 12'haaa;
rom[40388] = 12'haaa;
rom[40389] = 12'haaa;
rom[40390] = 12'haaa;
rom[40391] = 12'haaa;
rom[40392] = 12'haaa;
rom[40393] = 12'h999;
rom[40394] = 12'h999;
rom[40395] = 12'haaa;
rom[40396] = 12'haaa;
rom[40397] = 12'haaa;
rom[40398] = 12'haaa;
rom[40399] = 12'haaa;
rom[40400] = 12'h999;
rom[40401] = 12'h999;
rom[40402] = 12'h999;
rom[40403] = 12'h888;
rom[40404] = 12'h888;
rom[40405] = 12'h888;
rom[40406] = 12'h888;
rom[40407] = 12'h888;
rom[40408] = 12'h888;
rom[40409] = 12'h888;
rom[40410] = 12'h888;
rom[40411] = 12'h888;
rom[40412] = 12'h888;
rom[40413] = 12'h888;
rom[40414] = 12'h888;
rom[40415] = 12'h888;
rom[40416] = 12'h888;
rom[40417] = 12'h888;
rom[40418] = 12'h888;
rom[40419] = 12'h888;
rom[40420] = 12'h888;
rom[40421] = 12'h888;
rom[40422] = 12'h888;
rom[40423] = 12'h888;
rom[40424] = 12'h999;
rom[40425] = 12'h999;
rom[40426] = 12'h999;
rom[40427] = 12'h999;
rom[40428] = 12'h999;
rom[40429] = 12'h999;
rom[40430] = 12'h999;
rom[40431] = 12'h999;
rom[40432] = 12'h999;
rom[40433] = 12'h999;
rom[40434] = 12'h999;
rom[40435] = 12'h999;
rom[40436] = 12'h999;
rom[40437] = 12'h999;
rom[40438] = 12'h999;
rom[40439] = 12'h999;
rom[40440] = 12'haaa;
rom[40441] = 12'haaa;
rom[40442] = 12'haaa;
rom[40443] = 12'haaa;
rom[40444] = 12'hbbb;
rom[40445] = 12'hbbb;
rom[40446] = 12'hbbb;
rom[40447] = 12'hbbb;
rom[40448] = 12'hbbb;
rom[40449] = 12'hbbb;
rom[40450] = 12'hbbb;
rom[40451] = 12'hbbb;
rom[40452] = 12'hbbb;
rom[40453] = 12'hbbb;
rom[40454] = 12'haaa;
rom[40455] = 12'haaa;
rom[40456] = 12'haaa;
rom[40457] = 12'haaa;
rom[40458] = 12'h999;
rom[40459] = 12'h999;
rom[40460] = 12'h888;
rom[40461] = 12'h888;
rom[40462] = 12'h888;
rom[40463] = 12'h888;
rom[40464] = 12'h888;
rom[40465] = 12'h888;
rom[40466] = 12'h888;
rom[40467] = 12'h777;
rom[40468] = 12'h777;
rom[40469] = 12'h777;
rom[40470] = 12'h777;
rom[40471] = 12'h777;
rom[40472] = 12'h666;
rom[40473] = 12'h666;
rom[40474] = 12'h666;
rom[40475] = 12'h666;
rom[40476] = 12'h666;
rom[40477] = 12'h666;
rom[40478] = 12'h666;
rom[40479] = 12'h666;
rom[40480] = 12'h555;
rom[40481] = 12'h666;
rom[40482] = 12'h666;
rom[40483] = 12'h777;
rom[40484] = 12'h777;
rom[40485] = 12'h888;
rom[40486] = 12'h888;
rom[40487] = 12'h888;
rom[40488] = 12'h777;
rom[40489] = 12'h666;
rom[40490] = 12'h666;
rom[40491] = 12'h555;
rom[40492] = 12'h555;
rom[40493] = 12'h555;
rom[40494] = 12'h555;
rom[40495] = 12'h555;
rom[40496] = 12'h444;
rom[40497] = 12'h444;
rom[40498] = 12'h444;
rom[40499] = 12'h444;
rom[40500] = 12'h333;
rom[40501] = 12'h333;
rom[40502] = 12'h333;
rom[40503] = 12'h222;
rom[40504] = 12'h222;
rom[40505] = 12'h111;
rom[40506] = 12'h111;
rom[40507] = 12'h111;
rom[40508] = 12'h111;
rom[40509] = 12'h111;
rom[40510] = 12'h  0;
rom[40511] = 12'h  0;
rom[40512] = 12'h  0;
rom[40513] = 12'h  0;
rom[40514] = 12'h  0;
rom[40515] = 12'h  0;
rom[40516] = 12'h  0;
rom[40517] = 12'h  0;
rom[40518] = 12'h  0;
rom[40519] = 12'h  0;
rom[40520] = 12'h  0;
rom[40521] = 12'h  0;
rom[40522] = 12'h  0;
rom[40523] = 12'h  0;
rom[40524] = 12'h  0;
rom[40525] = 12'h  0;
rom[40526] = 12'h  0;
rom[40527] = 12'h  0;
rom[40528] = 12'h  0;
rom[40529] = 12'h  0;
rom[40530] = 12'h  0;
rom[40531] = 12'h  0;
rom[40532] = 12'h  0;
rom[40533] = 12'h  0;
rom[40534] = 12'h  0;
rom[40535] = 12'h  0;
rom[40536] = 12'h  0;
rom[40537] = 12'h  0;
rom[40538] = 12'h  0;
rom[40539] = 12'h  0;
rom[40540] = 12'h  0;
rom[40541] = 12'h  0;
rom[40542] = 12'h  0;
rom[40543] = 12'h  0;
rom[40544] = 12'h  0;
rom[40545] = 12'h  0;
rom[40546] = 12'h  0;
rom[40547] = 12'h  0;
rom[40548] = 12'h  0;
rom[40549] = 12'h  0;
rom[40550] = 12'h  0;
rom[40551] = 12'h  0;
rom[40552] = 12'h  0;
rom[40553] = 12'h  0;
rom[40554] = 12'h  0;
rom[40555] = 12'h  0;
rom[40556] = 12'h  0;
rom[40557] = 12'h  0;
rom[40558] = 12'h  0;
rom[40559] = 12'h  0;
rom[40560] = 12'h  0;
rom[40561] = 12'h  0;
rom[40562] = 12'h  0;
rom[40563] = 12'h  0;
rom[40564] = 12'h  0;
rom[40565] = 12'h  0;
rom[40566] = 12'h  0;
rom[40567] = 12'h  0;
rom[40568] = 12'h  0;
rom[40569] = 12'h  0;
rom[40570] = 12'h  0;
rom[40571] = 12'h  0;
rom[40572] = 12'h  0;
rom[40573] = 12'h  0;
rom[40574] = 12'h  0;
rom[40575] = 12'h  0;
rom[40576] = 12'h  0;
rom[40577] = 12'h  0;
rom[40578] = 12'h  0;
rom[40579] = 12'h  0;
rom[40580] = 12'h111;
rom[40581] = 12'h111;
rom[40582] = 12'h111;
rom[40583] = 12'h111;
rom[40584] = 12'h222;
rom[40585] = 12'h222;
rom[40586] = 12'h222;
rom[40587] = 12'h222;
rom[40588] = 12'h222;
rom[40589] = 12'h222;
rom[40590] = 12'h222;
rom[40591] = 12'h222;
rom[40592] = 12'h333;
rom[40593] = 12'h333;
rom[40594] = 12'h333;
rom[40595] = 12'h333;
rom[40596] = 12'h333;
rom[40597] = 12'h333;
rom[40598] = 12'h333;
rom[40599] = 12'h333;
rom[40600] = 12'h333;
rom[40601] = 12'h444;
rom[40602] = 12'h444;
rom[40603] = 12'h444;
rom[40604] = 12'h444;
rom[40605] = 12'h444;
rom[40606] = 12'h444;
rom[40607] = 12'h444;
rom[40608] = 12'h444;
rom[40609] = 12'h444;
rom[40610] = 12'h444;
rom[40611] = 12'h444;
rom[40612] = 12'h444;
rom[40613] = 12'h444;
rom[40614] = 12'h444;
rom[40615] = 12'h444;
rom[40616] = 12'h444;
rom[40617] = 12'h444;
rom[40618] = 12'h444;
rom[40619] = 12'h444;
rom[40620] = 12'h444;
rom[40621] = 12'h444;
rom[40622] = 12'h333;
rom[40623] = 12'h333;
rom[40624] = 12'h444;
rom[40625] = 12'h444;
rom[40626] = 12'h444;
rom[40627] = 12'h444;
rom[40628] = 12'h444;
rom[40629] = 12'h444;
rom[40630] = 12'h444;
rom[40631] = 12'h444;
rom[40632] = 12'h333;
rom[40633] = 12'h333;
rom[40634] = 12'h333;
rom[40635] = 12'h222;
rom[40636] = 12'h222;
rom[40637] = 12'h222;
rom[40638] = 12'h222;
rom[40639] = 12'h222;
rom[40640] = 12'h222;
rom[40641] = 12'h222;
rom[40642] = 12'h111;
rom[40643] = 12'h111;
rom[40644] = 12'h111;
rom[40645] = 12'h111;
rom[40646] = 12'h111;
rom[40647] = 12'h111;
rom[40648] = 12'h111;
rom[40649] = 12'h111;
rom[40650] = 12'h111;
rom[40651] = 12'h  0;
rom[40652] = 12'h  0;
rom[40653] = 12'h  0;
rom[40654] = 12'h  0;
rom[40655] = 12'h  0;
rom[40656] = 12'h  0;
rom[40657] = 12'h  0;
rom[40658] = 12'h  0;
rom[40659] = 12'h  0;
rom[40660] = 12'h  0;
rom[40661] = 12'h  0;
rom[40662] = 12'h  0;
rom[40663] = 12'h  0;
rom[40664] = 12'h  0;
rom[40665] = 12'h  0;
rom[40666] = 12'h  0;
rom[40667] = 12'h  0;
rom[40668] = 12'h  0;
rom[40669] = 12'h  0;
rom[40670] = 12'h  0;
rom[40671] = 12'h  0;
rom[40672] = 12'h  0;
rom[40673] = 12'h111;
rom[40674] = 12'h111;
rom[40675] = 12'h111;
rom[40676] = 12'h111;
rom[40677] = 12'h111;
rom[40678] = 12'h111;
rom[40679] = 12'h222;
rom[40680] = 12'h222;
rom[40681] = 12'h333;
rom[40682] = 12'h444;
rom[40683] = 12'h444;
rom[40684] = 12'h444;
rom[40685] = 12'h444;
rom[40686] = 12'h555;
rom[40687] = 12'h666;
rom[40688] = 12'h666;
rom[40689] = 12'h777;
rom[40690] = 12'h888;
rom[40691] = 12'h888;
rom[40692] = 12'h899;
rom[40693] = 12'h9a9;
rom[40694] = 12'habb;
rom[40695] = 12'hbbb;
rom[40696] = 12'hddd;
rom[40697] = 12'hfee;
rom[40698] = 12'hffe;
rom[40699] = 12'hdbb;
rom[40700] = 12'h854;
rom[40701] = 12'h511;
rom[40702] = 12'h521;
rom[40703] = 12'h621;
rom[40704] = 12'h610;
rom[40705] = 12'h710;
rom[40706] = 12'h720;
rom[40707] = 12'h820;
rom[40708] = 12'h820;
rom[40709] = 12'h820;
rom[40710] = 12'h920;
rom[40711] = 12'h920;
rom[40712] = 12'h920;
rom[40713] = 12'h820;
rom[40714] = 12'h820;
rom[40715] = 12'h810;
rom[40716] = 12'h710;
rom[40717] = 12'h610;
rom[40718] = 12'h610;
rom[40719] = 12'h610;
rom[40720] = 12'h500;
rom[40721] = 12'h500;
rom[40722] = 12'h500;
rom[40723] = 12'h500;
rom[40724] = 12'h500;
rom[40725] = 12'h500;
rom[40726] = 12'h500;
rom[40727] = 12'h600;
rom[40728] = 12'h600;
rom[40729] = 12'h710;
rom[40730] = 12'h710;
rom[40731] = 12'h810;
rom[40732] = 12'h920;
rom[40733] = 12'ha21;
rom[40734] = 12'ha21;
rom[40735] = 12'hb31;
rom[40736] = 12'hb31;
rom[40737] = 12'hb31;
rom[40738] = 12'hc31;
rom[40739] = 12'hc31;
rom[40740] = 12'hc31;
rom[40741] = 12'hc30;
rom[40742] = 12'hc30;
rom[40743] = 12'hc30;
rom[40744] = 12'hc30;
rom[40745] = 12'hb30;
rom[40746] = 12'hb40;
rom[40747] = 12'hc50;
rom[40748] = 12'hc61;
rom[40749] = 12'hc62;
rom[40750] = 12'hb61;
rom[40751] = 12'ha50;
rom[40752] = 12'h940;
rom[40753] = 12'h840;
rom[40754] = 12'h730;
rom[40755] = 12'h730;
rom[40756] = 12'h630;
rom[40757] = 12'h630;
rom[40758] = 12'h630;
rom[40759] = 12'h520;
rom[40760] = 12'h520;
rom[40761] = 12'h420;
rom[40762] = 12'h420;
rom[40763] = 12'h420;
rom[40764] = 12'h430;
rom[40765] = 12'h431;
rom[40766] = 12'h531;
rom[40767] = 12'h531;
rom[40768] = 12'h432;
rom[40769] = 12'h532;
rom[40770] = 12'h543;
rom[40771] = 12'h543;
rom[40772] = 12'h544;
rom[40773] = 12'h544;
rom[40774] = 12'h554;
rom[40775] = 12'h555;
rom[40776] = 12'h555;
rom[40777] = 12'h555;
rom[40778] = 12'h656;
rom[40779] = 12'h666;
rom[40780] = 12'h777;
rom[40781] = 12'h777;
rom[40782] = 12'h888;
rom[40783] = 12'h888;
rom[40784] = 12'h999;
rom[40785] = 12'h999;
rom[40786] = 12'h999;
rom[40787] = 12'haaa;
rom[40788] = 12'haaa;
rom[40789] = 12'haaa;
rom[40790] = 12'haaa;
rom[40791] = 12'haaa;
rom[40792] = 12'haaa;
rom[40793] = 12'h999;
rom[40794] = 12'h999;
rom[40795] = 12'h999;
rom[40796] = 12'haaa;
rom[40797] = 12'haaa;
rom[40798] = 12'haaa;
rom[40799] = 12'haaa;
rom[40800] = 12'h999;
rom[40801] = 12'h999;
rom[40802] = 12'h999;
rom[40803] = 12'h888;
rom[40804] = 12'h888;
rom[40805] = 12'h888;
rom[40806] = 12'h888;
rom[40807] = 12'h999;
rom[40808] = 12'h999;
rom[40809] = 12'h999;
rom[40810] = 12'h888;
rom[40811] = 12'h888;
rom[40812] = 12'h888;
rom[40813] = 12'h888;
rom[40814] = 12'h888;
rom[40815] = 12'h888;
rom[40816] = 12'h999;
rom[40817] = 12'h999;
rom[40818] = 12'h999;
rom[40819] = 12'h999;
rom[40820] = 12'h999;
rom[40821] = 12'h999;
rom[40822] = 12'h999;
rom[40823] = 12'h999;
rom[40824] = 12'h999;
rom[40825] = 12'h999;
rom[40826] = 12'h999;
rom[40827] = 12'h999;
rom[40828] = 12'h999;
rom[40829] = 12'h999;
rom[40830] = 12'h999;
rom[40831] = 12'h999;
rom[40832] = 12'h999;
rom[40833] = 12'h999;
rom[40834] = 12'h999;
rom[40835] = 12'h999;
rom[40836] = 12'h999;
rom[40837] = 12'h999;
rom[40838] = 12'haaa;
rom[40839] = 12'haaa;
rom[40840] = 12'haaa;
rom[40841] = 12'haaa;
rom[40842] = 12'haaa;
rom[40843] = 12'haaa;
rom[40844] = 12'hbbb;
rom[40845] = 12'hbbb;
rom[40846] = 12'hbbb;
rom[40847] = 12'hbbb;
rom[40848] = 12'hbbb;
rom[40849] = 12'hbbb;
rom[40850] = 12'hbbb;
rom[40851] = 12'hbbb;
rom[40852] = 12'hbbb;
rom[40853] = 12'hbbb;
rom[40854] = 12'haaa;
rom[40855] = 12'haaa;
rom[40856] = 12'haaa;
rom[40857] = 12'haaa;
rom[40858] = 12'h999;
rom[40859] = 12'h999;
rom[40860] = 12'h999;
rom[40861] = 12'h888;
rom[40862] = 12'h888;
rom[40863] = 12'h888;
rom[40864] = 12'h888;
rom[40865] = 12'h888;
rom[40866] = 12'h888;
rom[40867] = 12'h777;
rom[40868] = 12'h777;
rom[40869] = 12'h777;
rom[40870] = 12'h777;
rom[40871] = 12'h777;
rom[40872] = 12'h666;
rom[40873] = 12'h666;
rom[40874] = 12'h666;
rom[40875] = 12'h666;
rom[40876] = 12'h666;
rom[40877] = 12'h666;
rom[40878] = 12'h666;
rom[40879] = 12'h666;
rom[40880] = 12'h555;
rom[40881] = 12'h555;
rom[40882] = 12'h666;
rom[40883] = 12'h666;
rom[40884] = 12'h666;
rom[40885] = 12'h777;
rom[40886] = 12'h888;
rom[40887] = 12'h888;
rom[40888] = 12'h777;
rom[40889] = 12'h777;
rom[40890] = 12'h666;
rom[40891] = 12'h555;
rom[40892] = 12'h555;
rom[40893] = 12'h555;
rom[40894] = 12'h444;
rom[40895] = 12'h444;
rom[40896] = 12'h444;
rom[40897] = 12'h444;
rom[40898] = 12'h444;
rom[40899] = 12'h444;
rom[40900] = 12'h444;
rom[40901] = 12'h444;
rom[40902] = 12'h333;
rom[40903] = 12'h222;
rom[40904] = 12'h222;
rom[40905] = 12'h222;
rom[40906] = 12'h111;
rom[40907] = 12'h111;
rom[40908] = 12'h111;
rom[40909] = 12'h111;
rom[40910] = 12'h  0;
rom[40911] = 12'h  0;
rom[40912] = 12'h  0;
rom[40913] = 12'h  0;
rom[40914] = 12'h  0;
rom[40915] = 12'h  0;
rom[40916] = 12'h  0;
rom[40917] = 12'h  0;
rom[40918] = 12'h  0;
rom[40919] = 12'h  0;
rom[40920] = 12'h  0;
rom[40921] = 12'h  0;
rom[40922] = 12'h  0;
rom[40923] = 12'h  0;
rom[40924] = 12'h  0;
rom[40925] = 12'h  0;
rom[40926] = 12'h  0;
rom[40927] = 12'h  0;
rom[40928] = 12'h  0;
rom[40929] = 12'h  0;
rom[40930] = 12'h  0;
rom[40931] = 12'h  0;
rom[40932] = 12'h  0;
rom[40933] = 12'h  0;
rom[40934] = 12'h  0;
rom[40935] = 12'h  0;
rom[40936] = 12'h  0;
rom[40937] = 12'h  0;
rom[40938] = 12'h  0;
rom[40939] = 12'h  0;
rom[40940] = 12'h  0;
rom[40941] = 12'h  0;
rom[40942] = 12'h  0;
rom[40943] = 12'h  0;
rom[40944] = 12'h  0;
rom[40945] = 12'h  0;
rom[40946] = 12'h  0;
rom[40947] = 12'h  0;
rom[40948] = 12'h  0;
rom[40949] = 12'h  0;
rom[40950] = 12'h  0;
rom[40951] = 12'h  0;
rom[40952] = 12'h  0;
rom[40953] = 12'h  0;
rom[40954] = 12'h  0;
rom[40955] = 12'h  0;
rom[40956] = 12'h  0;
rom[40957] = 12'h  0;
rom[40958] = 12'h  0;
rom[40959] = 12'h  0;
rom[40960] = 12'h  0;
rom[40961] = 12'h  0;
rom[40962] = 12'h  0;
rom[40963] = 12'h  0;
rom[40964] = 12'h  0;
rom[40965] = 12'h  0;
rom[40966] = 12'h  0;
rom[40967] = 12'h  0;
rom[40968] = 12'h  0;
rom[40969] = 12'h  0;
rom[40970] = 12'h  0;
rom[40971] = 12'h  0;
rom[40972] = 12'h  0;
rom[40973] = 12'h  0;
rom[40974] = 12'h  0;
rom[40975] = 12'h  0;
rom[40976] = 12'h111;
rom[40977] = 12'h111;
rom[40978] = 12'h111;
rom[40979] = 12'h111;
rom[40980] = 12'h111;
rom[40981] = 12'h111;
rom[40982] = 12'h222;
rom[40983] = 12'h222;
rom[40984] = 12'h222;
rom[40985] = 12'h222;
rom[40986] = 12'h222;
rom[40987] = 12'h222;
rom[40988] = 12'h222;
rom[40989] = 12'h222;
rom[40990] = 12'h222;
rom[40991] = 12'h222;
rom[40992] = 12'h333;
rom[40993] = 12'h333;
rom[40994] = 12'h333;
rom[40995] = 12'h333;
rom[40996] = 12'h333;
rom[40997] = 12'h333;
rom[40998] = 12'h333;
rom[40999] = 12'h333;
rom[41000] = 12'h444;
rom[41001] = 12'h444;
rom[41002] = 12'h444;
rom[41003] = 12'h444;
rom[41004] = 12'h444;
rom[41005] = 12'h444;
rom[41006] = 12'h444;
rom[41007] = 12'h444;
rom[41008] = 12'h444;
rom[41009] = 12'h444;
rom[41010] = 12'h444;
rom[41011] = 12'h444;
rom[41012] = 12'h444;
rom[41013] = 12'h444;
rom[41014] = 12'h444;
rom[41015] = 12'h444;
rom[41016] = 12'h444;
rom[41017] = 12'h444;
rom[41018] = 12'h444;
rom[41019] = 12'h444;
rom[41020] = 12'h444;
rom[41021] = 12'h333;
rom[41022] = 12'h333;
rom[41023] = 12'h333;
rom[41024] = 12'h444;
rom[41025] = 12'h444;
rom[41026] = 12'h444;
rom[41027] = 12'h444;
rom[41028] = 12'h444;
rom[41029] = 12'h444;
rom[41030] = 12'h444;
rom[41031] = 12'h444;
rom[41032] = 12'h333;
rom[41033] = 12'h333;
rom[41034] = 12'h333;
rom[41035] = 12'h222;
rom[41036] = 12'h222;
rom[41037] = 12'h222;
rom[41038] = 12'h222;
rom[41039] = 12'h222;
rom[41040] = 12'h222;
rom[41041] = 12'h222;
rom[41042] = 12'h111;
rom[41043] = 12'h111;
rom[41044] = 12'h111;
rom[41045] = 12'h111;
rom[41046] = 12'h111;
rom[41047] = 12'h111;
rom[41048] = 12'h111;
rom[41049] = 12'h111;
rom[41050] = 12'h  0;
rom[41051] = 12'h  0;
rom[41052] = 12'h  0;
rom[41053] = 12'h  0;
rom[41054] = 12'h  0;
rom[41055] = 12'h  0;
rom[41056] = 12'h  0;
rom[41057] = 12'h  0;
rom[41058] = 12'h  0;
rom[41059] = 12'h  0;
rom[41060] = 12'h  0;
rom[41061] = 12'h  0;
rom[41062] = 12'h  0;
rom[41063] = 12'h  0;
rom[41064] = 12'h  0;
rom[41065] = 12'h  0;
rom[41066] = 12'h  0;
rom[41067] = 12'h  0;
rom[41068] = 12'h  0;
rom[41069] = 12'h  0;
rom[41070] = 12'h  0;
rom[41071] = 12'h  0;
rom[41072] = 12'h  0;
rom[41073] = 12'h111;
rom[41074] = 12'h111;
rom[41075] = 12'h111;
rom[41076] = 12'h111;
rom[41077] = 12'h222;
rom[41078] = 12'h222;
rom[41079] = 12'h222;
rom[41080] = 12'h333;
rom[41081] = 12'h444;
rom[41082] = 12'h444;
rom[41083] = 12'h444;
rom[41084] = 12'h444;
rom[41085] = 12'h555;
rom[41086] = 12'h555;
rom[41087] = 12'h666;
rom[41088] = 12'h666;
rom[41089] = 12'h877;
rom[41090] = 12'h888;
rom[41091] = 12'h999;
rom[41092] = 12'h999;
rom[41093] = 12'haaa;
rom[41094] = 12'hbbb;
rom[41095] = 12'hccb;
rom[41096] = 12'hedd;
rom[41097] = 12'hfee;
rom[41098] = 12'hfed;
rom[41099] = 12'hb98;
rom[41100] = 12'h633;
rom[41101] = 12'h511;
rom[41102] = 12'h621;
rom[41103] = 12'h610;
rom[41104] = 12'h610;
rom[41105] = 12'h710;
rom[41106] = 12'h710;
rom[41107] = 12'h820;
rom[41108] = 12'h810;
rom[41109] = 12'h810;
rom[41110] = 12'h810;
rom[41111] = 12'h920;
rom[41112] = 12'h920;
rom[41113] = 12'h920;
rom[41114] = 12'h920;
rom[41115] = 12'h820;
rom[41116] = 12'h820;
rom[41117] = 12'h720;
rom[41118] = 12'h710;
rom[41119] = 12'h710;
rom[41120] = 12'h710;
rom[41121] = 12'h710;
rom[41122] = 12'h710;
rom[41123] = 12'h710;
rom[41124] = 12'h710;
rom[41125] = 12'h710;
rom[41126] = 12'h710;
rom[41127] = 12'h810;
rom[41128] = 12'h810;
rom[41129] = 12'h920;
rom[41130] = 12'h921;
rom[41131] = 12'ha21;
rom[41132] = 12'ha31;
rom[41133] = 12'hb31;
rom[41134] = 12'hb31;
rom[41135] = 12'hb31;
rom[41136] = 12'hb31;
rom[41137] = 12'hb31;
rom[41138] = 12'hb31;
rom[41139] = 12'hb30;
rom[41140] = 12'hb30;
rom[41141] = 12'hb30;
rom[41142] = 12'hb30;
rom[41143] = 12'hb30;
rom[41144] = 12'hb30;
rom[41145] = 12'hb30;
rom[41146] = 12'hb40;
rom[41147] = 12'hb51;
rom[41148] = 12'hc61;
rom[41149] = 12'hb61;
rom[41150] = 12'ha50;
rom[41151] = 12'h940;
rom[41152] = 12'h840;
rom[41153] = 12'h730;
rom[41154] = 12'h730;
rom[41155] = 12'h630;
rom[41156] = 12'h630;
rom[41157] = 12'h630;
rom[41158] = 12'h530;
rom[41159] = 12'h520;
rom[41160] = 12'h420;
rom[41161] = 12'h420;
rom[41162] = 12'h430;
rom[41163] = 12'h430;
rom[41164] = 12'h431;
rom[41165] = 12'h431;
rom[41166] = 12'h431;
rom[41167] = 12'h431;
rom[41168] = 12'h432;
rom[41169] = 12'h532;
rom[41170] = 12'h543;
rom[41171] = 12'h543;
rom[41172] = 12'h544;
rom[41173] = 12'h554;
rom[41174] = 12'h555;
rom[41175] = 12'h555;
rom[41176] = 12'h665;
rom[41177] = 12'h666;
rom[41178] = 12'h666;
rom[41179] = 12'h777;
rom[41180] = 12'h777;
rom[41181] = 12'h888;
rom[41182] = 12'h888;
rom[41183] = 12'h888;
rom[41184] = 12'h999;
rom[41185] = 12'h999;
rom[41186] = 12'haaa;
rom[41187] = 12'haaa;
rom[41188] = 12'haaa;
rom[41189] = 12'haaa;
rom[41190] = 12'haaa;
rom[41191] = 12'haaa;
rom[41192] = 12'haaa;
rom[41193] = 12'h999;
rom[41194] = 12'h999;
rom[41195] = 12'h999;
rom[41196] = 12'haaa;
rom[41197] = 12'haaa;
rom[41198] = 12'haaa;
rom[41199] = 12'haaa;
rom[41200] = 12'h999;
rom[41201] = 12'h999;
rom[41202] = 12'h888;
rom[41203] = 12'h888;
rom[41204] = 12'h888;
rom[41205] = 12'h888;
rom[41206] = 12'h888;
rom[41207] = 12'h999;
rom[41208] = 12'h999;
rom[41209] = 12'h999;
rom[41210] = 12'h999;
rom[41211] = 12'h999;
rom[41212] = 12'h999;
rom[41213] = 12'h999;
rom[41214] = 12'h999;
rom[41215] = 12'h999;
rom[41216] = 12'h999;
rom[41217] = 12'h999;
rom[41218] = 12'h999;
rom[41219] = 12'h999;
rom[41220] = 12'h999;
rom[41221] = 12'h999;
rom[41222] = 12'h999;
rom[41223] = 12'h999;
rom[41224] = 12'h999;
rom[41225] = 12'h999;
rom[41226] = 12'h999;
rom[41227] = 12'h999;
rom[41228] = 12'h999;
rom[41229] = 12'h999;
rom[41230] = 12'h999;
rom[41231] = 12'h999;
rom[41232] = 12'h999;
rom[41233] = 12'h999;
rom[41234] = 12'h999;
rom[41235] = 12'h999;
rom[41236] = 12'h999;
rom[41237] = 12'h999;
rom[41238] = 12'h999;
rom[41239] = 12'h999;
rom[41240] = 12'haaa;
rom[41241] = 12'haaa;
rom[41242] = 12'haaa;
rom[41243] = 12'haaa;
rom[41244] = 12'haaa;
rom[41245] = 12'haaa;
rom[41246] = 12'hbbb;
rom[41247] = 12'hbbb;
rom[41248] = 12'hbbb;
rom[41249] = 12'hbbb;
rom[41250] = 12'hbbb;
rom[41251] = 12'hbbb;
rom[41252] = 12'hbbb;
rom[41253] = 12'hbbb;
rom[41254] = 12'hbbb;
rom[41255] = 12'haaa;
rom[41256] = 12'hbbb;
rom[41257] = 12'haaa;
rom[41258] = 12'haaa;
rom[41259] = 12'h999;
rom[41260] = 12'h999;
rom[41261] = 12'h999;
rom[41262] = 12'h888;
rom[41263] = 12'h888;
rom[41264] = 12'h888;
rom[41265] = 12'h888;
rom[41266] = 12'h888;
rom[41267] = 12'h777;
rom[41268] = 12'h777;
rom[41269] = 12'h777;
rom[41270] = 12'h777;
rom[41271] = 12'h777;
rom[41272] = 12'h666;
rom[41273] = 12'h666;
rom[41274] = 12'h666;
rom[41275] = 12'h666;
rom[41276] = 12'h666;
rom[41277] = 12'h666;
rom[41278] = 12'h555;
rom[41279] = 12'h555;
rom[41280] = 12'h555;
rom[41281] = 12'h555;
rom[41282] = 12'h555;
rom[41283] = 12'h555;
rom[41284] = 12'h666;
rom[41285] = 12'h777;
rom[41286] = 12'h777;
rom[41287] = 12'h777;
rom[41288] = 12'h888;
rom[41289] = 12'h777;
rom[41290] = 12'h666;
rom[41291] = 12'h666;
rom[41292] = 12'h555;
rom[41293] = 12'h555;
rom[41294] = 12'h444;
rom[41295] = 12'h444;
rom[41296] = 12'h444;
rom[41297] = 12'h333;
rom[41298] = 12'h333;
rom[41299] = 12'h333;
rom[41300] = 12'h444;
rom[41301] = 12'h444;
rom[41302] = 12'h333;
rom[41303] = 12'h222;
rom[41304] = 12'h222;
rom[41305] = 12'h222;
rom[41306] = 12'h222;
rom[41307] = 12'h111;
rom[41308] = 12'h111;
rom[41309] = 12'h111;
rom[41310] = 12'h111;
rom[41311] = 12'h  0;
rom[41312] = 12'h  0;
rom[41313] = 12'h  0;
rom[41314] = 12'h  0;
rom[41315] = 12'h  0;
rom[41316] = 12'h  0;
rom[41317] = 12'h  0;
rom[41318] = 12'h  0;
rom[41319] = 12'h  0;
rom[41320] = 12'h  0;
rom[41321] = 12'h  0;
rom[41322] = 12'h  0;
rom[41323] = 12'h  0;
rom[41324] = 12'h  0;
rom[41325] = 12'h  0;
rom[41326] = 12'h  0;
rom[41327] = 12'h  0;
rom[41328] = 12'h  0;
rom[41329] = 12'h  0;
rom[41330] = 12'h  0;
rom[41331] = 12'h  0;
rom[41332] = 12'h  0;
rom[41333] = 12'h  0;
rom[41334] = 12'h  0;
rom[41335] = 12'h  0;
rom[41336] = 12'h  0;
rom[41337] = 12'h  0;
rom[41338] = 12'h  0;
rom[41339] = 12'h  0;
rom[41340] = 12'h  0;
rom[41341] = 12'h  0;
rom[41342] = 12'h  0;
rom[41343] = 12'h  0;
rom[41344] = 12'h  0;
rom[41345] = 12'h  0;
rom[41346] = 12'h  0;
rom[41347] = 12'h  0;
rom[41348] = 12'h  0;
rom[41349] = 12'h  0;
rom[41350] = 12'h  0;
rom[41351] = 12'h  0;
rom[41352] = 12'h  0;
rom[41353] = 12'h  0;
rom[41354] = 12'h  0;
rom[41355] = 12'h  0;
rom[41356] = 12'h  0;
rom[41357] = 12'h  0;
rom[41358] = 12'h  0;
rom[41359] = 12'h  0;
rom[41360] = 12'h  0;
rom[41361] = 12'h  0;
rom[41362] = 12'h  0;
rom[41363] = 12'h  0;
rom[41364] = 12'h  0;
rom[41365] = 12'h  0;
rom[41366] = 12'h  0;
rom[41367] = 12'h  0;
rom[41368] = 12'h  0;
rom[41369] = 12'h  0;
rom[41370] = 12'h  0;
rom[41371] = 12'h  0;
rom[41372] = 12'h  0;
rom[41373] = 12'h  0;
rom[41374] = 12'h  0;
rom[41375] = 12'h  0;
rom[41376] = 12'h111;
rom[41377] = 12'h111;
rom[41378] = 12'h111;
rom[41379] = 12'h111;
rom[41380] = 12'h111;
rom[41381] = 12'h222;
rom[41382] = 12'h222;
rom[41383] = 12'h222;
rom[41384] = 12'h222;
rom[41385] = 12'h222;
rom[41386] = 12'h222;
rom[41387] = 12'h222;
rom[41388] = 12'h333;
rom[41389] = 12'h333;
rom[41390] = 12'h333;
rom[41391] = 12'h333;
rom[41392] = 12'h333;
rom[41393] = 12'h333;
rom[41394] = 12'h333;
rom[41395] = 12'h333;
rom[41396] = 12'h333;
rom[41397] = 12'h444;
rom[41398] = 12'h333;
rom[41399] = 12'h333;
rom[41400] = 12'h444;
rom[41401] = 12'h444;
rom[41402] = 12'h444;
rom[41403] = 12'h444;
rom[41404] = 12'h444;
rom[41405] = 12'h444;
rom[41406] = 12'h444;
rom[41407] = 12'h444;
rom[41408] = 12'h444;
rom[41409] = 12'h444;
rom[41410] = 12'h444;
rom[41411] = 12'h444;
rom[41412] = 12'h444;
rom[41413] = 12'h444;
rom[41414] = 12'h444;
rom[41415] = 12'h444;
rom[41416] = 12'h444;
rom[41417] = 12'h444;
rom[41418] = 12'h444;
rom[41419] = 12'h444;
rom[41420] = 12'h444;
rom[41421] = 12'h333;
rom[41422] = 12'h333;
rom[41423] = 12'h333;
rom[41424] = 12'h444;
rom[41425] = 12'h444;
rom[41426] = 12'h444;
rom[41427] = 12'h333;
rom[41428] = 12'h444;
rom[41429] = 12'h444;
rom[41430] = 12'h444;
rom[41431] = 12'h444;
rom[41432] = 12'h333;
rom[41433] = 12'h333;
rom[41434] = 12'h333;
rom[41435] = 12'h222;
rom[41436] = 12'h222;
rom[41437] = 12'h222;
rom[41438] = 12'h222;
rom[41439] = 12'h222;
rom[41440] = 12'h222;
rom[41441] = 12'h222;
rom[41442] = 12'h111;
rom[41443] = 12'h111;
rom[41444] = 12'h111;
rom[41445] = 12'h111;
rom[41446] = 12'h111;
rom[41447] = 12'h111;
rom[41448] = 12'h111;
rom[41449] = 12'h111;
rom[41450] = 12'h  0;
rom[41451] = 12'h  0;
rom[41452] = 12'h  0;
rom[41453] = 12'h  0;
rom[41454] = 12'h  0;
rom[41455] = 12'h  0;
rom[41456] = 12'h  0;
rom[41457] = 12'h  0;
rom[41458] = 12'h  0;
rom[41459] = 12'h  0;
rom[41460] = 12'h  0;
rom[41461] = 12'h  0;
rom[41462] = 12'h  0;
rom[41463] = 12'h  0;
rom[41464] = 12'h  0;
rom[41465] = 12'h  0;
rom[41466] = 12'h  0;
rom[41467] = 12'h  0;
rom[41468] = 12'h  0;
rom[41469] = 12'h  0;
rom[41470] = 12'h  0;
rom[41471] = 12'h  0;
rom[41472] = 12'h111;
rom[41473] = 12'h111;
rom[41474] = 12'h111;
rom[41475] = 12'h111;
rom[41476] = 12'h111;
rom[41477] = 12'h222;
rom[41478] = 12'h222;
rom[41479] = 12'h222;
rom[41480] = 12'h333;
rom[41481] = 12'h444;
rom[41482] = 12'h444;
rom[41483] = 12'h444;
rom[41484] = 12'h444;
rom[41485] = 12'h555;
rom[41486] = 12'h666;
rom[41487] = 12'h666;
rom[41488] = 12'h666;
rom[41489] = 12'h888;
rom[41490] = 12'h999;
rom[41491] = 12'h999;
rom[41492] = 12'h999;
rom[41493] = 12'haaa;
rom[41494] = 12'hbbb;
rom[41495] = 12'hccc;
rom[41496] = 12'hedd;
rom[41497] = 12'hfee;
rom[41498] = 12'hfdc;
rom[41499] = 12'h976;
rom[41500] = 12'h521;
rom[41501] = 12'h510;
rom[41502] = 12'h611;
rom[41503] = 12'h610;
rom[41504] = 12'h600;
rom[41505] = 12'h610;
rom[41506] = 12'h710;
rom[41507] = 12'h710;
rom[41508] = 12'h810;
rom[41509] = 12'h810;
rom[41510] = 12'h810;
rom[41511] = 12'h810;
rom[41512] = 12'h910;
rom[41513] = 12'h920;
rom[41514] = 12'h920;
rom[41515] = 12'h920;
rom[41516] = 12'h920;
rom[41517] = 12'h820;
rom[41518] = 12'h820;
rom[41519] = 12'h820;
rom[41520] = 12'h920;
rom[41521] = 12'h920;
rom[41522] = 12'h920;
rom[41523] = 12'h920;
rom[41524] = 12'h920;
rom[41525] = 12'h920;
rom[41526] = 12'h921;
rom[41527] = 12'h921;
rom[41528] = 12'h921;
rom[41529] = 12'ha21;
rom[41530] = 12'ha31;
rom[41531] = 12'hb31;
rom[41532] = 12'hb31;
rom[41533] = 12'hc31;
rom[41534] = 12'hc31;
rom[41535] = 12'hb31;
rom[41536] = 12'hb31;
rom[41537] = 12'hb31;
rom[41538] = 12'hb30;
rom[41539] = 12'hb20;
rom[41540] = 12'hb20;
rom[41541] = 12'ha20;
rom[41542] = 12'ha20;
rom[41543] = 12'ha20;
rom[41544] = 12'ha30;
rom[41545] = 12'ha30;
rom[41546] = 12'ha40;
rom[41547] = 12'hb51;
rom[41548] = 12'hb51;
rom[41549] = 12'ha51;
rom[41550] = 12'h940;
rom[41551] = 12'h830;
rom[41552] = 12'h830;
rom[41553] = 12'h730;
rom[41554] = 12'h730;
rom[41555] = 12'h630;
rom[41556] = 12'h630;
rom[41557] = 12'h630;
rom[41558] = 12'h520;
rom[41559] = 12'h520;
rom[41560] = 12'h420;
rom[41561] = 12'h420;
rom[41562] = 12'h430;
rom[41563] = 12'h431;
rom[41564] = 12'h431;
rom[41565] = 12'h431;
rom[41566] = 12'h431;
rom[41567] = 12'h431;
rom[41568] = 12'h432;
rom[41569] = 12'h542;
rom[41570] = 12'h543;
rom[41571] = 12'h543;
rom[41572] = 12'h554;
rom[41573] = 12'h554;
rom[41574] = 12'h555;
rom[41575] = 12'h555;
rom[41576] = 12'h666;
rom[41577] = 12'h666;
rom[41578] = 12'h767;
rom[41579] = 12'h777;
rom[41580] = 12'h877;
rom[41581] = 12'h888;
rom[41582] = 12'h888;
rom[41583] = 12'h888;
rom[41584] = 12'h999;
rom[41585] = 12'h999;
rom[41586] = 12'haaa;
rom[41587] = 12'haaa;
rom[41588] = 12'haaa;
rom[41589] = 12'haaa;
rom[41590] = 12'haaa;
rom[41591] = 12'haaa;
rom[41592] = 12'haaa;
rom[41593] = 12'h999;
rom[41594] = 12'h999;
rom[41595] = 12'h999;
rom[41596] = 12'haaa;
rom[41597] = 12'haaa;
rom[41598] = 12'haaa;
rom[41599] = 12'haaa;
rom[41600] = 12'h999;
rom[41601] = 12'h999;
rom[41602] = 12'h999;
rom[41603] = 12'h999;
rom[41604] = 12'h999;
rom[41605] = 12'h999;
rom[41606] = 12'h999;
rom[41607] = 12'h999;
rom[41608] = 12'h999;
rom[41609] = 12'h999;
rom[41610] = 12'h999;
rom[41611] = 12'h999;
rom[41612] = 12'h999;
rom[41613] = 12'h999;
rom[41614] = 12'h999;
rom[41615] = 12'h999;
rom[41616] = 12'h999;
rom[41617] = 12'h999;
rom[41618] = 12'h999;
rom[41619] = 12'h999;
rom[41620] = 12'h999;
rom[41621] = 12'h999;
rom[41622] = 12'h888;
rom[41623] = 12'h888;
rom[41624] = 12'h888;
rom[41625] = 12'h888;
rom[41626] = 12'h888;
rom[41627] = 12'h888;
rom[41628] = 12'h888;
rom[41629] = 12'h888;
rom[41630] = 12'h888;
rom[41631] = 12'h888;
rom[41632] = 12'h888;
rom[41633] = 12'h888;
rom[41634] = 12'h888;
rom[41635] = 12'h888;
rom[41636] = 12'h888;
rom[41637] = 12'h888;
rom[41638] = 12'h999;
rom[41639] = 12'h999;
rom[41640] = 12'h999;
rom[41641] = 12'h999;
rom[41642] = 12'h999;
rom[41643] = 12'h999;
rom[41644] = 12'haaa;
rom[41645] = 12'haaa;
rom[41646] = 12'haaa;
rom[41647] = 12'haaa;
rom[41648] = 12'haaa;
rom[41649] = 12'hbbb;
rom[41650] = 12'hbbb;
rom[41651] = 12'hbbb;
rom[41652] = 12'hbbb;
rom[41653] = 12'hbbb;
rom[41654] = 12'hbbb;
rom[41655] = 12'haaa;
rom[41656] = 12'hbbb;
rom[41657] = 12'haaa;
rom[41658] = 12'haaa;
rom[41659] = 12'haaa;
rom[41660] = 12'h999;
rom[41661] = 12'h999;
rom[41662] = 12'h999;
rom[41663] = 12'h888;
rom[41664] = 12'h888;
rom[41665] = 12'h888;
rom[41666] = 12'h888;
rom[41667] = 12'h888;
rom[41668] = 12'h888;
rom[41669] = 12'h777;
rom[41670] = 12'h777;
rom[41671] = 12'h777;
rom[41672] = 12'h777;
rom[41673] = 12'h666;
rom[41674] = 12'h666;
rom[41675] = 12'h666;
rom[41676] = 12'h666;
rom[41677] = 12'h666;
rom[41678] = 12'h666;
rom[41679] = 12'h555;
rom[41680] = 12'h555;
rom[41681] = 12'h555;
rom[41682] = 12'h555;
rom[41683] = 12'h555;
rom[41684] = 12'h555;
rom[41685] = 12'h666;
rom[41686] = 12'h777;
rom[41687] = 12'h777;
rom[41688] = 12'h777;
rom[41689] = 12'h777;
rom[41690] = 12'h777;
rom[41691] = 12'h666;
rom[41692] = 12'h666;
rom[41693] = 12'h555;
rom[41694] = 12'h444;
rom[41695] = 12'h444;
rom[41696] = 12'h444;
rom[41697] = 12'h444;
rom[41698] = 12'h333;
rom[41699] = 12'h333;
rom[41700] = 12'h333;
rom[41701] = 12'h333;
rom[41702] = 12'h333;
rom[41703] = 12'h333;
rom[41704] = 12'h333;
rom[41705] = 12'h222;
rom[41706] = 12'h222;
rom[41707] = 12'h111;
rom[41708] = 12'h111;
rom[41709] = 12'h111;
rom[41710] = 12'h111;
rom[41711] = 12'h111;
rom[41712] = 12'h111;
rom[41713] = 12'h  0;
rom[41714] = 12'h  0;
rom[41715] = 12'h  0;
rom[41716] = 12'h  0;
rom[41717] = 12'h  0;
rom[41718] = 12'h  0;
rom[41719] = 12'h  0;
rom[41720] = 12'h  0;
rom[41721] = 12'h  0;
rom[41722] = 12'h  0;
rom[41723] = 12'h  0;
rom[41724] = 12'h  0;
rom[41725] = 12'h  0;
rom[41726] = 12'h  0;
rom[41727] = 12'h  0;
rom[41728] = 12'h  0;
rom[41729] = 12'h  0;
rom[41730] = 12'h  0;
rom[41731] = 12'h  0;
rom[41732] = 12'h  0;
rom[41733] = 12'h  0;
rom[41734] = 12'h  0;
rom[41735] = 12'h  0;
rom[41736] = 12'h  0;
rom[41737] = 12'h  0;
rom[41738] = 12'h  0;
rom[41739] = 12'h  0;
rom[41740] = 12'h  0;
rom[41741] = 12'h  0;
rom[41742] = 12'h  0;
rom[41743] = 12'h  0;
rom[41744] = 12'h  0;
rom[41745] = 12'h  0;
rom[41746] = 12'h  0;
rom[41747] = 12'h  0;
rom[41748] = 12'h  0;
rom[41749] = 12'h  0;
rom[41750] = 12'h  0;
rom[41751] = 12'h  0;
rom[41752] = 12'h  0;
rom[41753] = 12'h  0;
rom[41754] = 12'h  0;
rom[41755] = 12'h  0;
rom[41756] = 12'h  0;
rom[41757] = 12'h  0;
rom[41758] = 12'h  0;
rom[41759] = 12'h  0;
rom[41760] = 12'h  0;
rom[41761] = 12'h  0;
rom[41762] = 12'h  0;
rom[41763] = 12'h  0;
rom[41764] = 12'h  0;
rom[41765] = 12'h  0;
rom[41766] = 12'h  0;
rom[41767] = 12'h  0;
rom[41768] = 12'h  0;
rom[41769] = 12'h  0;
rom[41770] = 12'h  0;
rom[41771] = 12'h111;
rom[41772] = 12'h111;
rom[41773] = 12'h111;
rom[41774] = 12'h111;
rom[41775] = 12'h111;
rom[41776] = 12'h111;
rom[41777] = 12'h111;
rom[41778] = 12'h222;
rom[41779] = 12'h222;
rom[41780] = 12'h222;
rom[41781] = 12'h222;
rom[41782] = 12'h222;
rom[41783] = 12'h222;
rom[41784] = 12'h222;
rom[41785] = 12'h222;
rom[41786] = 12'h222;
rom[41787] = 12'h333;
rom[41788] = 12'h333;
rom[41789] = 12'h333;
rom[41790] = 12'h333;
rom[41791] = 12'h333;
rom[41792] = 12'h333;
rom[41793] = 12'h333;
rom[41794] = 12'h333;
rom[41795] = 12'h333;
rom[41796] = 12'h333;
rom[41797] = 12'h333;
rom[41798] = 12'h333;
rom[41799] = 12'h333;
rom[41800] = 12'h444;
rom[41801] = 12'h444;
rom[41802] = 12'h444;
rom[41803] = 12'h444;
rom[41804] = 12'h444;
rom[41805] = 12'h444;
rom[41806] = 12'h444;
rom[41807] = 12'h444;
rom[41808] = 12'h444;
rom[41809] = 12'h444;
rom[41810] = 12'h444;
rom[41811] = 12'h444;
rom[41812] = 12'h444;
rom[41813] = 12'h444;
rom[41814] = 12'h444;
rom[41815] = 12'h444;
rom[41816] = 12'h444;
rom[41817] = 12'h444;
rom[41818] = 12'h444;
rom[41819] = 12'h444;
rom[41820] = 12'h444;
rom[41821] = 12'h444;
rom[41822] = 12'h333;
rom[41823] = 12'h333;
rom[41824] = 12'h444;
rom[41825] = 12'h444;
rom[41826] = 12'h333;
rom[41827] = 12'h333;
rom[41828] = 12'h333;
rom[41829] = 12'h333;
rom[41830] = 12'h333;
rom[41831] = 12'h333;
rom[41832] = 12'h333;
rom[41833] = 12'h333;
rom[41834] = 12'h222;
rom[41835] = 12'h222;
rom[41836] = 12'h222;
rom[41837] = 12'h222;
rom[41838] = 12'h222;
rom[41839] = 12'h222;
rom[41840] = 12'h222;
rom[41841] = 12'h222;
rom[41842] = 12'h111;
rom[41843] = 12'h111;
rom[41844] = 12'h111;
rom[41845] = 12'h111;
rom[41846] = 12'h111;
rom[41847] = 12'h111;
rom[41848] = 12'h111;
rom[41849] = 12'h111;
rom[41850] = 12'h  0;
rom[41851] = 12'h  0;
rom[41852] = 12'h  0;
rom[41853] = 12'h  0;
rom[41854] = 12'h  0;
rom[41855] = 12'h  0;
rom[41856] = 12'h  0;
rom[41857] = 12'h  0;
rom[41858] = 12'h  0;
rom[41859] = 12'h  0;
rom[41860] = 12'h  0;
rom[41861] = 12'h  0;
rom[41862] = 12'h  0;
rom[41863] = 12'h  0;
rom[41864] = 12'h  0;
rom[41865] = 12'h  0;
rom[41866] = 12'h  0;
rom[41867] = 12'h  0;
rom[41868] = 12'h  0;
rom[41869] = 12'h  0;
rom[41870] = 12'h  0;
rom[41871] = 12'h  0;
rom[41872] = 12'h111;
rom[41873] = 12'h111;
rom[41874] = 12'h111;
rom[41875] = 12'h222;
rom[41876] = 12'h222;
rom[41877] = 12'h222;
rom[41878] = 12'h222;
rom[41879] = 12'h333;
rom[41880] = 12'h444;
rom[41881] = 12'h444;
rom[41882] = 12'h444;
rom[41883] = 12'h444;
rom[41884] = 12'h555;
rom[41885] = 12'h555;
rom[41886] = 12'h666;
rom[41887] = 12'h666;
rom[41888] = 12'h887;
rom[41889] = 12'h887;
rom[41890] = 12'h777;
rom[41891] = 12'h888;
rom[41892] = 12'h999;
rom[41893] = 12'haaa;
rom[41894] = 12'hbbb;
rom[41895] = 12'hddc;
rom[41896] = 12'hedd;
rom[41897] = 12'hfff;
rom[41898] = 12'hdbb;
rom[41899] = 12'h743;
rom[41900] = 12'h521;
rom[41901] = 12'h621;
rom[41902] = 12'h510;
rom[41903] = 12'h500;
rom[41904] = 12'h610;
rom[41905] = 12'h610;
rom[41906] = 12'h610;
rom[41907] = 12'h710;
rom[41908] = 12'h710;
rom[41909] = 12'h710;
rom[41910] = 12'h810;
rom[41911] = 12'h810;
rom[41912] = 12'h810;
rom[41913] = 12'h810;
rom[41914] = 12'h810;
rom[41915] = 12'h810;
rom[41916] = 12'h810;
rom[41917] = 12'h820;
rom[41918] = 12'h820;
rom[41919] = 12'h820;
rom[41920] = 12'h920;
rom[41921] = 12'h920;
rom[41922] = 12'h920;
rom[41923] = 12'h920;
rom[41924] = 12'h921;
rom[41925] = 12'ha21;
rom[41926] = 12'ha21;
rom[41927] = 12'ha21;
rom[41928] = 12'ha31;
rom[41929] = 12'ha31;
rom[41930] = 12'ha21;
rom[41931] = 12'ha21;
rom[41932] = 12'hb20;
rom[41933] = 12'hb20;
rom[41934] = 12'hb20;
rom[41935] = 12'hb20;
rom[41936] = 12'ha20;
rom[41937] = 12'ha20;
rom[41938] = 12'ha20;
rom[41939] = 12'ha20;
rom[41940] = 12'ha20;
rom[41941] = 12'ha20;
rom[41942] = 12'ha20;
rom[41943] = 12'h920;
rom[41944] = 12'h920;
rom[41945] = 12'ha30;
rom[41946] = 12'ha41;
rom[41947] = 12'ha51;
rom[41948] = 12'ha51;
rom[41949] = 12'h940;
rom[41950] = 12'h840;
rom[41951] = 12'h830;
rom[41952] = 12'h730;
rom[41953] = 12'h720;
rom[41954] = 12'h620;
rom[41955] = 12'h620;
rom[41956] = 12'h620;
rom[41957] = 12'h630;
rom[41958] = 12'h530;
rom[41959] = 12'h530;
rom[41960] = 12'h420;
rom[41961] = 12'h430;
rom[41962] = 12'h431;
rom[41963] = 12'h431;
rom[41964] = 12'h431;
rom[41965] = 12'h431;
rom[41966] = 12'h431;
rom[41967] = 12'h432;
rom[41968] = 12'h532;
rom[41969] = 12'h543;
rom[41970] = 12'h543;
rom[41971] = 12'h544;
rom[41972] = 12'h554;
rom[41973] = 12'h555;
rom[41974] = 12'h655;
rom[41975] = 12'h655;
rom[41976] = 12'h777;
rom[41977] = 12'h777;
rom[41978] = 12'h777;
rom[41979] = 12'h777;
rom[41980] = 12'h878;
rom[41981] = 12'h888;
rom[41982] = 12'h999;
rom[41983] = 12'h999;
rom[41984] = 12'haaa;
rom[41985] = 12'haaa;
rom[41986] = 12'haaa;
rom[41987] = 12'haaa;
rom[41988] = 12'haaa;
rom[41989] = 12'haaa;
rom[41990] = 12'haaa;
rom[41991] = 12'haaa;
rom[41992] = 12'haaa;
rom[41993] = 12'haaa;
rom[41994] = 12'h999;
rom[41995] = 12'h999;
rom[41996] = 12'haaa;
rom[41997] = 12'haaa;
rom[41998] = 12'haaa;
rom[41999] = 12'haaa;
rom[42000] = 12'h999;
rom[42001] = 12'h999;
rom[42002] = 12'h999;
rom[42003] = 12'h999;
rom[42004] = 12'h999;
rom[42005] = 12'h999;
rom[42006] = 12'h999;
rom[42007] = 12'h999;
rom[42008] = 12'h999;
rom[42009] = 12'h999;
rom[42010] = 12'h999;
rom[42011] = 12'h999;
rom[42012] = 12'h999;
rom[42013] = 12'h999;
rom[42014] = 12'h888;
rom[42015] = 12'h888;
rom[42016] = 12'h888;
rom[42017] = 12'h888;
rom[42018] = 12'h888;
rom[42019] = 12'h888;
rom[42020] = 12'h888;
rom[42021] = 12'h888;
rom[42022] = 12'h888;
rom[42023] = 12'h888;
rom[42024] = 12'h888;
rom[42025] = 12'h888;
rom[42026] = 12'h888;
rom[42027] = 12'h888;
rom[42028] = 12'h888;
rom[42029] = 12'h888;
rom[42030] = 12'h888;
rom[42031] = 12'h888;
rom[42032] = 12'h888;
rom[42033] = 12'h888;
rom[42034] = 12'h888;
rom[42035] = 12'h888;
rom[42036] = 12'h888;
rom[42037] = 12'h888;
rom[42038] = 12'h888;
rom[42039] = 12'h888;
rom[42040] = 12'h999;
rom[42041] = 12'h999;
rom[42042] = 12'h999;
rom[42043] = 12'h999;
rom[42044] = 12'h999;
rom[42045] = 12'h999;
rom[42046] = 12'haaa;
rom[42047] = 12'haaa;
rom[42048] = 12'haaa;
rom[42049] = 12'hbbb;
rom[42050] = 12'hbbb;
rom[42051] = 12'hbbb;
rom[42052] = 12'hbbb;
rom[42053] = 12'hbbb;
rom[42054] = 12'hbbb;
rom[42055] = 12'hbbb;
rom[42056] = 12'hbbb;
rom[42057] = 12'hbbb;
rom[42058] = 12'haaa;
rom[42059] = 12'haaa;
rom[42060] = 12'haaa;
rom[42061] = 12'h999;
rom[42062] = 12'h999;
rom[42063] = 12'h888;
rom[42064] = 12'h888;
rom[42065] = 12'h888;
rom[42066] = 12'h888;
rom[42067] = 12'h888;
rom[42068] = 12'h888;
rom[42069] = 12'h777;
rom[42070] = 12'h777;
rom[42071] = 12'h777;
rom[42072] = 12'h777;
rom[42073] = 12'h666;
rom[42074] = 12'h666;
rom[42075] = 12'h666;
rom[42076] = 12'h666;
rom[42077] = 12'h666;
rom[42078] = 12'h666;
rom[42079] = 12'h666;
rom[42080] = 12'h555;
rom[42081] = 12'h555;
rom[42082] = 12'h555;
rom[42083] = 12'h555;
rom[42084] = 12'h555;
rom[42085] = 12'h666;
rom[42086] = 12'h666;
rom[42087] = 12'h777;
rom[42088] = 12'h777;
rom[42089] = 12'h777;
rom[42090] = 12'h777;
rom[42091] = 12'h666;
rom[42092] = 12'h666;
rom[42093] = 12'h555;
rom[42094] = 12'h555;
rom[42095] = 12'h444;
rom[42096] = 12'h444;
rom[42097] = 12'h444;
rom[42098] = 12'h333;
rom[42099] = 12'h333;
rom[42100] = 12'h333;
rom[42101] = 12'h333;
rom[42102] = 12'h333;
rom[42103] = 12'h333;
rom[42104] = 12'h333;
rom[42105] = 12'h222;
rom[42106] = 12'h222;
rom[42107] = 12'h222;
rom[42108] = 12'h111;
rom[42109] = 12'h111;
rom[42110] = 12'h111;
rom[42111] = 12'h  0;
rom[42112] = 12'h111;
rom[42113] = 12'h  0;
rom[42114] = 12'h  0;
rom[42115] = 12'h  0;
rom[42116] = 12'h  0;
rom[42117] = 12'h  0;
rom[42118] = 12'h  0;
rom[42119] = 12'h  0;
rom[42120] = 12'h  0;
rom[42121] = 12'h  0;
rom[42122] = 12'h  0;
rom[42123] = 12'h  0;
rom[42124] = 12'h  0;
rom[42125] = 12'h  0;
rom[42126] = 12'h  0;
rom[42127] = 12'h  0;
rom[42128] = 12'h  0;
rom[42129] = 12'h  0;
rom[42130] = 12'h  0;
rom[42131] = 12'h  0;
rom[42132] = 12'h  0;
rom[42133] = 12'h  0;
rom[42134] = 12'h  0;
rom[42135] = 12'h  0;
rom[42136] = 12'h  0;
rom[42137] = 12'h  0;
rom[42138] = 12'h  0;
rom[42139] = 12'h  0;
rom[42140] = 12'h  0;
rom[42141] = 12'h  0;
rom[42142] = 12'h  0;
rom[42143] = 12'h  0;
rom[42144] = 12'h  0;
rom[42145] = 12'h  0;
rom[42146] = 12'h  0;
rom[42147] = 12'h  0;
rom[42148] = 12'h  0;
rom[42149] = 12'h  0;
rom[42150] = 12'h  0;
rom[42151] = 12'h  0;
rom[42152] = 12'h  0;
rom[42153] = 12'h  0;
rom[42154] = 12'h  0;
rom[42155] = 12'h  0;
rom[42156] = 12'h  0;
rom[42157] = 12'h  0;
rom[42158] = 12'h  0;
rom[42159] = 12'h  0;
rom[42160] = 12'h  0;
rom[42161] = 12'h  0;
rom[42162] = 12'h  0;
rom[42163] = 12'h  0;
rom[42164] = 12'h  0;
rom[42165] = 12'h  0;
rom[42166] = 12'h  0;
rom[42167] = 12'h111;
rom[42168] = 12'h111;
rom[42169] = 12'h111;
rom[42170] = 12'h111;
rom[42171] = 12'h111;
rom[42172] = 12'h111;
rom[42173] = 12'h222;
rom[42174] = 12'h222;
rom[42175] = 12'h222;
rom[42176] = 12'h222;
rom[42177] = 12'h222;
rom[42178] = 12'h222;
rom[42179] = 12'h222;
rom[42180] = 12'h222;
rom[42181] = 12'h222;
rom[42182] = 12'h222;
rom[42183] = 12'h222;
rom[42184] = 12'h222;
rom[42185] = 12'h222;
rom[42186] = 12'h222;
rom[42187] = 12'h333;
rom[42188] = 12'h333;
rom[42189] = 12'h333;
rom[42190] = 12'h333;
rom[42191] = 12'h333;
rom[42192] = 12'h333;
rom[42193] = 12'h333;
rom[42194] = 12'h333;
rom[42195] = 12'h333;
rom[42196] = 12'h333;
rom[42197] = 12'h333;
rom[42198] = 12'h333;
rom[42199] = 12'h333;
rom[42200] = 12'h444;
rom[42201] = 12'h444;
rom[42202] = 12'h444;
rom[42203] = 12'h444;
rom[42204] = 12'h444;
rom[42205] = 12'h444;
rom[42206] = 12'h444;
rom[42207] = 12'h444;
rom[42208] = 12'h444;
rom[42209] = 12'h444;
rom[42210] = 12'h444;
rom[42211] = 12'h444;
rom[42212] = 12'h444;
rom[42213] = 12'h444;
rom[42214] = 12'h444;
rom[42215] = 12'h444;
rom[42216] = 12'h444;
rom[42217] = 12'h444;
rom[42218] = 12'h444;
rom[42219] = 12'h444;
rom[42220] = 12'h444;
rom[42221] = 12'h444;
rom[42222] = 12'h444;
rom[42223] = 12'h444;
rom[42224] = 12'h444;
rom[42225] = 12'h444;
rom[42226] = 12'h333;
rom[42227] = 12'h333;
rom[42228] = 12'h333;
rom[42229] = 12'h333;
rom[42230] = 12'h333;
rom[42231] = 12'h333;
rom[42232] = 12'h333;
rom[42233] = 12'h333;
rom[42234] = 12'h222;
rom[42235] = 12'h222;
rom[42236] = 12'h222;
rom[42237] = 12'h222;
rom[42238] = 12'h222;
rom[42239] = 12'h222;
rom[42240] = 12'h222;
rom[42241] = 12'h222;
rom[42242] = 12'h222;
rom[42243] = 12'h111;
rom[42244] = 12'h111;
rom[42245] = 12'h111;
rom[42246] = 12'h111;
rom[42247] = 12'h111;
rom[42248] = 12'h111;
rom[42249] = 12'h  0;
rom[42250] = 12'h  0;
rom[42251] = 12'h  0;
rom[42252] = 12'h  0;
rom[42253] = 12'h  0;
rom[42254] = 12'h  0;
rom[42255] = 12'h  0;
rom[42256] = 12'h  0;
rom[42257] = 12'h  0;
rom[42258] = 12'h  0;
rom[42259] = 12'h  0;
rom[42260] = 12'h  0;
rom[42261] = 12'h  0;
rom[42262] = 12'h  0;
rom[42263] = 12'h  0;
rom[42264] = 12'h  0;
rom[42265] = 12'h  0;
rom[42266] = 12'h  0;
rom[42267] = 12'h  0;
rom[42268] = 12'h  0;
rom[42269] = 12'h  0;
rom[42270] = 12'h  0;
rom[42271] = 12'h  0;
rom[42272] = 12'h111;
rom[42273] = 12'h111;
rom[42274] = 12'h111;
rom[42275] = 12'h222;
rom[42276] = 12'h222;
rom[42277] = 12'h222;
rom[42278] = 12'h222;
rom[42279] = 12'h333;
rom[42280] = 12'h444;
rom[42281] = 12'h444;
rom[42282] = 12'h444;
rom[42283] = 12'h555;
rom[42284] = 12'h555;
rom[42285] = 12'h555;
rom[42286] = 12'h666;
rom[42287] = 12'h777;
rom[42288] = 12'h777;
rom[42289] = 12'h888;
rom[42290] = 12'h888;
rom[42291] = 12'h888;
rom[42292] = 12'h999;
rom[42293] = 12'haaa;
rom[42294] = 12'hbbb;
rom[42295] = 12'hddd;
rom[42296] = 12'hedd;
rom[42297] = 12'hfee;
rom[42298] = 12'hb99;
rom[42299] = 12'h632;
rom[42300] = 12'h511;
rom[42301] = 12'h511;
rom[42302] = 12'h510;
rom[42303] = 12'h500;
rom[42304] = 12'h610;
rom[42305] = 12'h610;
rom[42306] = 12'h610;
rom[42307] = 12'h610;
rom[42308] = 12'h710;
rom[42309] = 12'h710;
rom[42310] = 12'h710;
rom[42311] = 12'h710;
rom[42312] = 12'h710;
rom[42313] = 12'h810;
rom[42314] = 12'h810;
rom[42315] = 12'h810;
rom[42316] = 12'h810;
rom[42317] = 12'h810;
rom[42318] = 12'h810;
rom[42319] = 12'h820;
rom[42320] = 12'h920;
rom[42321] = 12'h920;
rom[42322] = 12'h920;
rom[42323] = 12'h920;
rom[42324] = 12'h920;
rom[42325] = 12'h920;
rom[42326] = 12'h920;
rom[42327] = 12'h920;
rom[42328] = 12'ha21;
rom[42329] = 12'ha21;
rom[42330] = 12'ha20;
rom[42331] = 12'ha20;
rom[42332] = 12'ha20;
rom[42333] = 12'ha20;
rom[42334] = 12'ha20;
rom[42335] = 12'ha20;
rom[42336] = 12'ha20;
rom[42337] = 12'h920;
rom[42338] = 12'h920;
rom[42339] = 12'h920;
rom[42340] = 12'h910;
rom[42341] = 12'h920;
rom[42342] = 12'h920;
rom[42343] = 12'h920;
rom[42344] = 12'h920;
rom[42345] = 12'h930;
rom[42346] = 12'h941;
rom[42347] = 12'h941;
rom[42348] = 12'h941;
rom[42349] = 12'h840;
rom[42350] = 12'h830;
rom[42351] = 12'h730;
rom[42352] = 12'h730;
rom[42353] = 12'h620;
rom[42354] = 12'h620;
rom[42355] = 12'h620;
rom[42356] = 12'h620;
rom[42357] = 12'h530;
rom[42358] = 12'h530;
rom[42359] = 12'h530;
rom[42360] = 12'h430;
rom[42361] = 12'h430;
rom[42362] = 12'h431;
rom[42363] = 12'h431;
rom[42364] = 12'h431;
rom[42365] = 12'h431;
rom[42366] = 12'h432;
rom[42367] = 12'h432;
rom[42368] = 12'h432;
rom[42369] = 12'h543;
rom[42370] = 12'h543;
rom[42371] = 12'h544;
rom[42372] = 12'h554;
rom[42373] = 12'h655;
rom[42374] = 12'h665;
rom[42375] = 12'h666;
rom[42376] = 12'h767;
rom[42377] = 12'h777;
rom[42378] = 12'h777;
rom[42379] = 12'h778;
rom[42380] = 12'h888;
rom[42381] = 12'h888;
rom[42382] = 12'h999;
rom[42383] = 12'h999;
rom[42384] = 12'haaa;
rom[42385] = 12'haaa;
rom[42386] = 12'haaa;
rom[42387] = 12'haaa;
rom[42388] = 12'haaa;
rom[42389] = 12'haaa;
rom[42390] = 12'haaa;
rom[42391] = 12'haaa;
rom[42392] = 12'haaa;
rom[42393] = 12'haaa;
rom[42394] = 12'h999;
rom[42395] = 12'h999;
rom[42396] = 12'haaa;
rom[42397] = 12'haaa;
rom[42398] = 12'haaa;
rom[42399] = 12'haaa;
rom[42400] = 12'h999;
rom[42401] = 12'h999;
rom[42402] = 12'h999;
rom[42403] = 12'h999;
rom[42404] = 12'h999;
rom[42405] = 12'h999;
rom[42406] = 12'h999;
rom[42407] = 12'h999;
rom[42408] = 12'h888;
rom[42409] = 12'h888;
rom[42410] = 12'h888;
rom[42411] = 12'h888;
rom[42412] = 12'h888;
rom[42413] = 12'h888;
rom[42414] = 12'h888;
rom[42415] = 12'h888;
rom[42416] = 12'h777;
rom[42417] = 12'h777;
rom[42418] = 12'h777;
rom[42419] = 12'h777;
rom[42420] = 12'h777;
rom[42421] = 12'h777;
rom[42422] = 12'h777;
rom[42423] = 12'h777;
rom[42424] = 12'h777;
rom[42425] = 12'h777;
rom[42426] = 12'h777;
rom[42427] = 12'h777;
rom[42428] = 12'h777;
rom[42429] = 12'h777;
rom[42430] = 12'h777;
rom[42431] = 12'h777;
rom[42432] = 12'h777;
rom[42433] = 12'h777;
rom[42434] = 12'h777;
rom[42435] = 12'h888;
rom[42436] = 12'h888;
rom[42437] = 12'h888;
rom[42438] = 12'h888;
rom[42439] = 12'h888;
rom[42440] = 12'h888;
rom[42441] = 12'h888;
rom[42442] = 12'h888;
rom[42443] = 12'h999;
rom[42444] = 12'h999;
rom[42445] = 12'h999;
rom[42446] = 12'h999;
rom[42447] = 12'h999;
rom[42448] = 12'haaa;
rom[42449] = 12'haaa;
rom[42450] = 12'haaa;
rom[42451] = 12'hbbb;
rom[42452] = 12'hbbb;
rom[42453] = 12'hbbb;
rom[42454] = 12'hbbb;
rom[42455] = 12'hbbb;
rom[42456] = 12'hbbb;
rom[42457] = 12'hbbb;
rom[42458] = 12'hbbb;
rom[42459] = 12'haaa;
rom[42460] = 12'haaa;
rom[42461] = 12'haaa;
rom[42462] = 12'h999;
rom[42463] = 12'h999;
rom[42464] = 12'h999;
rom[42465] = 12'h888;
rom[42466] = 12'h888;
rom[42467] = 12'h888;
rom[42468] = 12'h888;
rom[42469] = 12'h777;
rom[42470] = 12'h777;
rom[42471] = 12'h777;
rom[42472] = 12'h777;
rom[42473] = 12'h777;
rom[42474] = 12'h666;
rom[42475] = 12'h666;
rom[42476] = 12'h666;
rom[42477] = 12'h666;
rom[42478] = 12'h666;
rom[42479] = 12'h666;
rom[42480] = 12'h555;
rom[42481] = 12'h555;
rom[42482] = 12'h555;
rom[42483] = 12'h555;
rom[42484] = 12'h555;
rom[42485] = 12'h666;
rom[42486] = 12'h666;
rom[42487] = 12'h666;
rom[42488] = 12'h777;
rom[42489] = 12'h777;
rom[42490] = 12'h777;
rom[42491] = 12'h777;
rom[42492] = 12'h666;
rom[42493] = 12'h666;
rom[42494] = 12'h555;
rom[42495] = 12'h555;
rom[42496] = 12'h444;
rom[42497] = 12'h444;
rom[42498] = 12'h444;
rom[42499] = 12'h333;
rom[42500] = 12'h333;
rom[42501] = 12'h333;
rom[42502] = 12'h333;
rom[42503] = 12'h333;
rom[42504] = 12'h333;
rom[42505] = 12'h333;
rom[42506] = 12'h222;
rom[42507] = 12'h222;
rom[42508] = 12'h222;
rom[42509] = 12'h111;
rom[42510] = 12'h111;
rom[42511] = 12'h  0;
rom[42512] = 12'h  0;
rom[42513] = 12'h  0;
rom[42514] = 12'h  0;
rom[42515] = 12'h  0;
rom[42516] = 12'h  0;
rom[42517] = 12'h  0;
rom[42518] = 12'h  0;
rom[42519] = 12'h  0;
rom[42520] = 12'h  0;
rom[42521] = 12'h  0;
rom[42522] = 12'h  0;
rom[42523] = 12'h  0;
rom[42524] = 12'h  0;
rom[42525] = 12'h  0;
rom[42526] = 12'h  0;
rom[42527] = 12'h  0;
rom[42528] = 12'h  0;
rom[42529] = 12'h  0;
rom[42530] = 12'h  0;
rom[42531] = 12'h  0;
rom[42532] = 12'h  0;
rom[42533] = 12'h  0;
rom[42534] = 12'h  0;
rom[42535] = 12'h  0;
rom[42536] = 12'h  0;
rom[42537] = 12'h  0;
rom[42538] = 12'h  0;
rom[42539] = 12'h  0;
rom[42540] = 12'h  0;
rom[42541] = 12'h  0;
rom[42542] = 12'h  0;
rom[42543] = 12'h  0;
rom[42544] = 12'h  0;
rom[42545] = 12'h  0;
rom[42546] = 12'h  0;
rom[42547] = 12'h  0;
rom[42548] = 12'h  0;
rom[42549] = 12'h  0;
rom[42550] = 12'h  0;
rom[42551] = 12'h  0;
rom[42552] = 12'h  0;
rom[42553] = 12'h  0;
rom[42554] = 12'h  0;
rom[42555] = 12'h  0;
rom[42556] = 12'h  0;
rom[42557] = 12'h  0;
rom[42558] = 12'h  0;
rom[42559] = 12'h  0;
rom[42560] = 12'h  0;
rom[42561] = 12'h  0;
rom[42562] = 12'h  0;
rom[42563] = 12'h  0;
rom[42564] = 12'h111;
rom[42565] = 12'h111;
rom[42566] = 12'h111;
rom[42567] = 12'h111;
rom[42568] = 12'h111;
rom[42569] = 12'h111;
rom[42570] = 12'h111;
rom[42571] = 12'h222;
rom[42572] = 12'h222;
rom[42573] = 12'h222;
rom[42574] = 12'h222;
rom[42575] = 12'h222;
rom[42576] = 12'h222;
rom[42577] = 12'h222;
rom[42578] = 12'h222;
rom[42579] = 12'h222;
rom[42580] = 12'h222;
rom[42581] = 12'h222;
rom[42582] = 12'h333;
rom[42583] = 12'h333;
rom[42584] = 12'h222;
rom[42585] = 12'h222;
rom[42586] = 12'h222;
rom[42587] = 12'h333;
rom[42588] = 12'h333;
rom[42589] = 12'h333;
rom[42590] = 12'h333;
rom[42591] = 12'h333;
rom[42592] = 12'h333;
rom[42593] = 12'h333;
rom[42594] = 12'h333;
rom[42595] = 12'h333;
rom[42596] = 12'h333;
rom[42597] = 12'h333;
rom[42598] = 12'h333;
rom[42599] = 12'h333;
rom[42600] = 12'h333;
rom[42601] = 12'h333;
rom[42602] = 12'h333;
rom[42603] = 12'h444;
rom[42604] = 12'h444;
rom[42605] = 12'h444;
rom[42606] = 12'h444;
rom[42607] = 12'h444;
rom[42608] = 12'h444;
rom[42609] = 12'h444;
rom[42610] = 12'h444;
rom[42611] = 12'h444;
rom[42612] = 12'h444;
rom[42613] = 12'h444;
rom[42614] = 12'h444;
rom[42615] = 12'h444;
rom[42616] = 12'h444;
rom[42617] = 12'h444;
rom[42618] = 12'h444;
rom[42619] = 12'h444;
rom[42620] = 12'h444;
rom[42621] = 12'h444;
rom[42622] = 12'h444;
rom[42623] = 12'h444;
rom[42624] = 12'h444;
rom[42625] = 12'h333;
rom[42626] = 12'h333;
rom[42627] = 12'h333;
rom[42628] = 12'h333;
rom[42629] = 12'h333;
rom[42630] = 12'h333;
rom[42631] = 12'h333;
rom[42632] = 12'h333;
rom[42633] = 12'h333;
rom[42634] = 12'h222;
rom[42635] = 12'h222;
rom[42636] = 12'h222;
rom[42637] = 12'h222;
rom[42638] = 12'h222;
rom[42639] = 12'h222;
rom[42640] = 12'h222;
rom[42641] = 12'h222;
rom[42642] = 12'h222;
rom[42643] = 12'h111;
rom[42644] = 12'h111;
rom[42645] = 12'h111;
rom[42646] = 12'h111;
rom[42647] = 12'h111;
rom[42648] = 12'h  0;
rom[42649] = 12'h  0;
rom[42650] = 12'h  0;
rom[42651] = 12'h  0;
rom[42652] = 12'h  0;
rom[42653] = 12'h  0;
rom[42654] = 12'h  0;
rom[42655] = 12'h  0;
rom[42656] = 12'h  0;
rom[42657] = 12'h  0;
rom[42658] = 12'h  0;
rom[42659] = 12'h  0;
rom[42660] = 12'h  0;
rom[42661] = 12'h  0;
rom[42662] = 12'h  0;
rom[42663] = 12'h  0;
rom[42664] = 12'h  0;
rom[42665] = 12'h  0;
rom[42666] = 12'h  0;
rom[42667] = 12'h  0;
rom[42668] = 12'h  0;
rom[42669] = 12'h  0;
rom[42670] = 12'h111;
rom[42671] = 12'h111;
rom[42672] = 12'h111;
rom[42673] = 12'h111;
rom[42674] = 12'h111;
rom[42675] = 12'h222;
rom[42676] = 12'h222;
rom[42677] = 12'h222;
rom[42678] = 12'h333;
rom[42679] = 12'h444;
rom[42680] = 12'h444;
rom[42681] = 12'h444;
rom[42682] = 12'h555;
rom[42683] = 12'h555;
rom[42684] = 12'h555;
rom[42685] = 12'h666;
rom[42686] = 12'h666;
rom[42687] = 12'h777;
rom[42688] = 12'h777;
rom[42689] = 12'h888;
rom[42690] = 12'h888;
rom[42691] = 12'h899;
rom[42692] = 12'h9a9;
rom[42693] = 12'haaa;
rom[42694] = 12'hbbb;
rom[42695] = 12'hddd;
rom[42696] = 12'hfee;
rom[42697] = 12'hecc;
rom[42698] = 12'h976;
rom[42699] = 12'h421;
rom[42700] = 12'h410;
rom[42701] = 12'h511;
rom[42702] = 12'h510;
rom[42703] = 12'h500;
rom[42704] = 12'h610;
rom[42705] = 12'h610;
rom[42706] = 12'h610;
rom[42707] = 12'h610;
rom[42708] = 12'h610;
rom[42709] = 12'h610;
rom[42710] = 12'h610;
rom[42711] = 12'h710;
rom[42712] = 12'h710;
rom[42713] = 12'h710;
rom[42714] = 12'h710;
rom[42715] = 12'h710;
rom[42716] = 12'h710;
rom[42717] = 12'h710;
rom[42718] = 12'h710;
rom[42719] = 12'h810;
rom[42720] = 12'h810;
rom[42721] = 12'h810;
rom[42722] = 12'h810;
rom[42723] = 12'h810;
rom[42724] = 12'h810;
rom[42725] = 12'h820;
rom[42726] = 12'h920;
rom[42727] = 12'h920;
rom[42728] = 12'h910;
rom[42729] = 12'h910;
rom[42730] = 12'h910;
rom[42731] = 12'h910;
rom[42732] = 12'h910;
rom[42733] = 12'h910;
rom[42734] = 12'h910;
rom[42735] = 12'h810;
rom[42736] = 12'h810;
rom[42737] = 12'h810;
rom[42738] = 12'h810;
rom[42739] = 12'h810;
rom[42740] = 12'h810;
rom[42741] = 12'h810;
rom[42742] = 12'h810;
rom[42743] = 12'h820;
rom[42744] = 12'h820;
rom[42745] = 12'h830;
rom[42746] = 12'h930;
rom[42747] = 12'h840;
rom[42748] = 12'h830;
rom[42749] = 12'h830;
rom[42750] = 12'h730;
rom[42751] = 12'h730;
rom[42752] = 12'h720;
rom[42753] = 12'h620;
rom[42754] = 12'h620;
rom[42755] = 12'h620;
rom[42756] = 12'h520;
rom[42757] = 12'h530;
rom[42758] = 12'h530;
rom[42759] = 12'h530;
rom[42760] = 12'h430;
rom[42761] = 12'h431;
rom[42762] = 12'h431;
rom[42763] = 12'h431;
rom[42764] = 12'h431;
rom[42765] = 12'h432;
rom[42766] = 12'h432;
rom[42767] = 12'h432;
rom[42768] = 12'h432;
rom[42769] = 12'h543;
rom[42770] = 12'h543;
rom[42771] = 12'h554;
rom[42772] = 12'h655;
rom[42773] = 12'h665;
rom[42774] = 12'h666;
rom[42775] = 12'h666;
rom[42776] = 12'h677;
rom[42777] = 12'h777;
rom[42778] = 12'h777;
rom[42779] = 12'h788;
rom[42780] = 12'h888;
rom[42781] = 12'h999;
rom[42782] = 12'h999;
rom[42783] = 12'haaa;
rom[42784] = 12'haaa;
rom[42785] = 12'haaa;
rom[42786] = 12'haaa;
rom[42787] = 12'haaa;
rom[42788] = 12'haaa;
rom[42789] = 12'haaa;
rom[42790] = 12'haaa;
rom[42791] = 12'haaa;
rom[42792] = 12'haaa;
rom[42793] = 12'h999;
rom[42794] = 12'h999;
rom[42795] = 12'h999;
rom[42796] = 12'haaa;
rom[42797] = 12'haaa;
rom[42798] = 12'haaa;
rom[42799] = 12'haaa;
rom[42800] = 12'h999;
rom[42801] = 12'h999;
rom[42802] = 12'h999;
rom[42803] = 12'h888;
rom[42804] = 12'h888;
rom[42805] = 12'h888;
rom[42806] = 12'h888;
rom[42807] = 12'h888;
rom[42808] = 12'h777;
rom[42809] = 12'h777;
rom[42810] = 12'h777;
rom[42811] = 12'h777;
rom[42812] = 12'h777;
rom[42813] = 12'h777;
rom[42814] = 12'h777;
rom[42815] = 12'h777;
rom[42816] = 12'h777;
rom[42817] = 12'h777;
rom[42818] = 12'h777;
rom[42819] = 12'h777;
rom[42820] = 12'h777;
rom[42821] = 12'h777;
rom[42822] = 12'h777;
rom[42823] = 12'h777;
rom[42824] = 12'h777;
rom[42825] = 12'h777;
rom[42826] = 12'h777;
rom[42827] = 12'h777;
rom[42828] = 12'h777;
rom[42829] = 12'h777;
rom[42830] = 12'h777;
rom[42831] = 12'h777;
rom[42832] = 12'h777;
rom[42833] = 12'h777;
rom[42834] = 12'h777;
rom[42835] = 12'h888;
rom[42836] = 12'h888;
rom[42837] = 12'h888;
rom[42838] = 12'h888;
rom[42839] = 12'h888;
rom[42840] = 12'h888;
rom[42841] = 12'h888;
rom[42842] = 12'h888;
rom[42843] = 12'h888;
rom[42844] = 12'h888;
rom[42845] = 12'h888;
rom[42846] = 12'h999;
rom[42847] = 12'h999;
rom[42848] = 12'h999;
rom[42849] = 12'h999;
rom[42850] = 12'haaa;
rom[42851] = 12'haaa;
rom[42852] = 12'haaa;
rom[42853] = 12'haaa;
rom[42854] = 12'hbbb;
rom[42855] = 12'hbbb;
rom[42856] = 12'hbbb;
rom[42857] = 12'hbbb;
rom[42858] = 12'hbbb;
rom[42859] = 12'hbbb;
rom[42860] = 12'hbbb;
rom[42861] = 12'haaa;
rom[42862] = 12'h999;
rom[42863] = 12'h999;
rom[42864] = 12'h999;
rom[42865] = 12'h888;
rom[42866] = 12'h888;
rom[42867] = 12'h888;
rom[42868] = 12'h777;
rom[42869] = 12'h777;
rom[42870] = 12'h777;
rom[42871] = 12'h777;
rom[42872] = 12'h777;
rom[42873] = 12'h777;
rom[42874] = 12'h666;
rom[42875] = 12'h666;
rom[42876] = 12'h666;
rom[42877] = 12'h666;
rom[42878] = 12'h666;
rom[42879] = 12'h666;
rom[42880] = 12'h666;
rom[42881] = 12'h666;
rom[42882] = 12'h555;
rom[42883] = 12'h555;
rom[42884] = 12'h555;
rom[42885] = 12'h555;
rom[42886] = 12'h666;
rom[42887] = 12'h666;
rom[42888] = 12'h666;
rom[42889] = 12'h666;
rom[42890] = 12'h777;
rom[42891] = 12'h777;
rom[42892] = 12'h777;
rom[42893] = 12'h666;
rom[42894] = 12'h555;
rom[42895] = 12'h555;
rom[42896] = 12'h444;
rom[42897] = 12'h444;
rom[42898] = 12'h444;
rom[42899] = 12'h333;
rom[42900] = 12'h333;
rom[42901] = 12'h333;
rom[42902] = 12'h333;
rom[42903] = 12'h333;
rom[42904] = 12'h333;
rom[42905] = 12'h333;
rom[42906] = 12'h333;
rom[42907] = 12'h222;
rom[42908] = 12'h222;
rom[42909] = 12'h111;
rom[42910] = 12'h111;
rom[42911] = 12'h111;
rom[42912] = 12'h  0;
rom[42913] = 12'h  0;
rom[42914] = 12'h  0;
rom[42915] = 12'h  0;
rom[42916] = 12'h  0;
rom[42917] = 12'h  0;
rom[42918] = 12'h  0;
rom[42919] = 12'h  0;
rom[42920] = 12'h  0;
rom[42921] = 12'h  0;
rom[42922] = 12'h  0;
rom[42923] = 12'h  0;
rom[42924] = 12'h  0;
rom[42925] = 12'h  0;
rom[42926] = 12'h  0;
rom[42927] = 12'h  0;
rom[42928] = 12'h  0;
rom[42929] = 12'h  0;
rom[42930] = 12'h  0;
rom[42931] = 12'h  0;
rom[42932] = 12'h  0;
rom[42933] = 12'h  0;
rom[42934] = 12'h  0;
rom[42935] = 12'h  0;
rom[42936] = 12'h  0;
rom[42937] = 12'h  0;
rom[42938] = 12'h  0;
rom[42939] = 12'h  0;
rom[42940] = 12'h  0;
rom[42941] = 12'h  0;
rom[42942] = 12'h  0;
rom[42943] = 12'h  0;
rom[42944] = 12'h  0;
rom[42945] = 12'h  0;
rom[42946] = 12'h  0;
rom[42947] = 12'h  0;
rom[42948] = 12'h  0;
rom[42949] = 12'h  0;
rom[42950] = 12'h  0;
rom[42951] = 12'h  0;
rom[42952] = 12'h  0;
rom[42953] = 12'h  0;
rom[42954] = 12'h  0;
rom[42955] = 12'h  0;
rom[42956] = 12'h  0;
rom[42957] = 12'h  0;
rom[42958] = 12'h  0;
rom[42959] = 12'h  0;
rom[42960] = 12'h  0;
rom[42961] = 12'h  0;
rom[42962] = 12'h111;
rom[42963] = 12'h111;
rom[42964] = 12'h111;
rom[42965] = 12'h111;
rom[42966] = 12'h111;
rom[42967] = 12'h111;
rom[42968] = 12'h111;
rom[42969] = 12'h111;
rom[42970] = 12'h222;
rom[42971] = 12'h222;
rom[42972] = 12'h222;
rom[42973] = 12'h222;
rom[42974] = 12'h222;
rom[42975] = 12'h222;
rom[42976] = 12'h222;
rom[42977] = 12'h222;
rom[42978] = 12'h222;
rom[42979] = 12'h222;
rom[42980] = 12'h222;
rom[42981] = 12'h222;
rom[42982] = 12'h333;
rom[42983] = 12'h333;
rom[42984] = 12'h222;
rom[42985] = 12'h222;
rom[42986] = 12'h222;
rom[42987] = 12'h222;
rom[42988] = 12'h333;
rom[42989] = 12'h333;
rom[42990] = 12'h333;
rom[42991] = 12'h333;
rom[42992] = 12'h333;
rom[42993] = 12'h333;
rom[42994] = 12'h333;
rom[42995] = 12'h333;
rom[42996] = 12'h333;
rom[42997] = 12'h333;
rom[42998] = 12'h333;
rom[42999] = 12'h333;
rom[43000] = 12'h333;
rom[43001] = 12'h333;
rom[43002] = 12'h333;
rom[43003] = 12'h333;
rom[43004] = 12'h333;
rom[43005] = 12'h333;
rom[43006] = 12'h333;
rom[43007] = 12'h333;
rom[43008] = 12'h444;
rom[43009] = 12'h444;
rom[43010] = 12'h444;
rom[43011] = 12'h444;
rom[43012] = 12'h444;
rom[43013] = 12'h444;
rom[43014] = 12'h444;
rom[43015] = 12'h444;
rom[43016] = 12'h444;
rom[43017] = 12'h444;
rom[43018] = 12'h444;
rom[43019] = 12'h444;
rom[43020] = 12'h444;
rom[43021] = 12'h444;
rom[43022] = 12'h444;
rom[43023] = 12'h444;
rom[43024] = 12'h444;
rom[43025] = 12'h333;
rom[43026] = 12'h333;
rom[43027] = 12'h333;
rom[43028] = 12'h333;
rom[43029] = 12'h333;
rom[43030] = 12'h333;
rom[43031] = 12'h333;
rom[43032] = 12'h333;
rom[43033] = 12'h333;
rom[43034] = 12'h222;
rom[43035] = 12'h222;
rom[43036] = 12'h222;
rom[43037] = 12'h222;
rom[43038] = 12'h222;
rom[43039] = 12'h222;
rom[43040] = 12'h222;
rom[43041] = 12'h222;
rom[43042] = 12'h111;
rom[43043] = 12'h111;
rom[43044] = 12'h111;
rom[43045] = 12'h111;
rom[43046] = 12'h111;
rom[43047] = 12'h111;
rom[43048] = 12'h  0;
rom[43049] = 12'h  0;
rom[43050] = 12'h  0;
rom[43051] = 12'h  0;
rom[43052] = 12'h  0;
rom[43053] = 12'h  0;
rom[43054] = 12'h  0;
rom[43055] = 12'h  0;
rom[43056] = 12'h  0;
rom[43057] = 12'h  0;
rom[43058] = 12'h  0;
rom[43059] = 12'h  0;
rom[43060] = 12'h  0;
rom[43061] = 12'h  0;
rom[43062] = 12'h  0;
rom[43063] = 12'h  0;
rom[43064] = 12'h  0;
rom[43065] = 12'h  0;
rom[43066] = 12'h  0;
rom[43067] = 12'h  0;
rom[43068] = 12'h  0;
rom[43069] = 12'h  0;
rom[43070] = 12'h111;
rom[43071] = 12'h111;
rom[43072] = 12'h111;
rom[43073] = 12'h111;
rom[43074] = 12'h222;
rom[43075] = 12'h222;
rom[43076] = 12'h222;
rom[43077] = 12'h222;
rom[43078] = 12'h333;
rom[43079] = 12'h444;
rom[43080] = 12'h444;
rom[43081] = 12'h555;
rom[43082] = 12'h555;
rom[43083] = 12'h555;
rom[43084] = 12'h555;
rom[43085] = 12'h666;
rom[43086] = 12'h777;
rom[43087] = 12'h777;
rom[43088] = 12'h777;
rom[43089] = 12'h888;
rom[43090] = 12'h888;
rom[43091] = 12'h999;
rom[43092] = 12'h9aa;
rom[43093] = 12'haaa;
rom[43094] = 12'hbbb;
rom[43095] = 12'hddd;
rom[43096] = 12'hfee;
rom[43097] = 12'hcba;
rom[43098] = 12'h654;
rom[43099] = 12'h311;
rom[43100] = 12'h410;
rom[43101] = 12'h511;
rom[43102] = 12'h510;
rom[43103] = 12'h500;
rom[43104] = 12'h510;
rom[43105] = 12'h510;
rom[43106] = 12'h500;
rom[43107] = 12'h500;
rom[43108] = 12'h500;
rom[43109] = 12'h500;
rom[43110] = 12'h600;
rom[43111] = 12'h600;
rom[43112] = 12'h600;
rom[43113] = 12'h600;
rom[43114] = 12'h600;
rom[43115] = 12'h600;
rom[43116] = 12'h600;
rom[43117] = 12'h710;
rom[43118] = 12'h710;
rom[43119] = 12'h710;
rom[43120] = 12'h710;
rom[43121] = 12'h710;
rom[43122] = 12'h710;
rom[43123] = 12'h710;
rom[43124] = 12'h710;
rom[43125] = 12'h710;
rom[43126] = 12'h810;
rom[43127] = 12'h810;
rom[43128] = 12'h810;
rom[43129] = 12'h710;
rom[43130] = 12'h710;
rom[43131] = 12'h810;
rom[43132] = 12'h710;
rom[43133] = 12'h700;
rom[43134] = 12'h700;
rom[43135] = 12'h700;
rom[43136] = 12'h710;
rom[43137] = 12'h710;
rom[43138] = 12'h710;
rom[43139] = 12'h710;
rom[43140] = 12'h710;
rom[43141] = 12'h710;
rom[43142] = 12'h710;
rom[43143] = 12'h710;
rom[43144] = 12'h820;
rom[43145] = 12'h820;
rom[43146] = 12'h830;
rom[43147] = 12'h830;
rom[43148] = 12'h730;
rom[43149] = 12'h730;
rom[43150] = 12'h720;
rom[43151] = 12'h720;
rom[43152] = 12'h620;
rom[43153] = 12'h620;
rom[43154] = 12'h620;
rom[43155] = 12'h520;
rom[43156] = 12'h520;
rom[43157] = 12'h520;
rom[43158] = 12'h530;
rom[43159] = 12'h530;
rom[43160] = 12'h431;
rom[43161] = 12'h431;
rom[43162] = 12'h431;
rom[43163] = 12'h432;
rom[43164] = 12'h432;
rom[43165] = 12'h432;
rom[43166] = 12'h532;
rom[43167] = 12'h543;
rom[43168] = 12'h543;
rom[43169] = 12'h543;
rom[43170] = 12'h554;
rom[43171] = 12'h654;
rom[43172] = 12'h665;
rom[43173] = 12'h666;
rom[43174] = 12'h766;
rom[43175] = 12'h777;
rom[43176] = 12'h677;
rom[43177] = 12'h777;
rom[43178] = 12'h778;
rom[43179] = 12'h888;
rom[43180] = 12'h889;
rom[43181] = 12'h999;
rom[43182] = 12'haaa;
rom[43183] = 12'haaa;
rom[43184] = 12'hbab;
rom[43185] = 12'hbbb;
rom[43186] = 12'hbbb;
rom[43187] = 12'hbbb;
rom[43188] = 12'haaa;
rom[43189] = 12'haaa;
rom[43190] = 12'haaa;
rom[43191] = 12'haaa;
rom[43192] = 12'haaa;
rom[43193] = 12'h999;
rom[43194] = 12'h999;
rom[43195] = 12'h999;
rom[43196] = 12'haaa;
rom[43197] = 12'haaa;
rom[43198] = 12'haaa;
rom[43199] = 12'haaa;
rom[43200] = 12'h888;
rom[43201] = 12'h888;
rom[43202] = 12'h888;
rom[43203] = 12'h888;
rom[43204] = 12'h777;
rom[43205] = 12'h777;
rom[43206] = 12'h777;
rom[43207] = 12'h777;
rom[43208] = 12'h888;
rom[43209] = 12'h777;
rom[43210] = 12'h777;
rom[43211] = 12'h777;
rom[43212] = 12'h777;
rom[43213] = 12'h777;
rom[43214] = 12'h777;
rom[43215] = 12'h777;
rom[43216] = 12'h777;
rom[43217] = 12'h777;
rom[43218] = 12'h666;
rom[43219] = 12'h666;
rom[43220] = 12'h666;
rom[43221] = 12'h777;
rom[43222] = 12'h777;
rom[43223] = 12'h777;
rom[43224] = 12'h777;
rom[43225] = 12'h777;
rom[43226] = 12'h777;
rom[43227] = 12'h777;
rom[43228] = 12'h777;
rom[43229] = 12'h777;
rom[43230] = 12'h777;
rom[43231] = 12'h777;
rom[43232] = 12'h777;
rom[43233] = 12'h777;
rom[43234] = 12'h777;
rom[43235] = 12'h888;
rom[43236] = 12'h888;
rom[43237] = 12'h888;
rom[43238] = 12'h888;
rom[43239] = 12'h888;
rom[43240] = 12'h888;
rom[43241] = 12'h888;
rom[43242] = 12'h888;
rom[43243] = 12'h888;
rom[43244] = 12'h888;
rom[43245] = 12'h888;
rom[43246] = 12'h888;
rom[43247] = 12'h999;
rom[43248] = 12'h999;
rom[43249] = 12'h999;
rom[43250] = 12'h999;
rom[43251] = 12'h999;
rom[43252] = 12'h999;
rom[43253] = 12'haaa;
rom[43254] = 12'haaa;
rom[43255] = 12'hbbb;
rom[43256] = 12'hbbb;
rom[43257] = 12'hbbb;
rom[43258] = 12'hbbb;
rom[43259] = 12'hbbb;
rom[43260] = 12'hbbb;
rom[43261] = 12'haaa;
rom[43262] = 12'haaa;
rom[43263] = 12'h999;
rom[43264] = 12'h999;
rom[43265] = 12'h999;
rom[43266] = 12'h888;
rom[43267] = 12'h888;
rom[43268] = 12'h777;
rom[43269] = 12'h777;
rom[43270] = 12'h777;
rom[43271] = 12'h777;
rom[43272] = 12'h777;
rom[43273] = 12'h777;
rom[43274] = 12'h666;
rom[43275] = 12'h666;
rom[43276] = 12'h666;
rom[43277] = 12'h666;
rom[43278] = 12'h666;
rom[43279] = 12'h666;
rom[43280] = 12'h666;
rom[43281] = 12'h666;
rom[43282] = 12'h666;
rom[43283] = 12'h666;
rom[43284] = 12'h555;
rom[43285] = 12'h555;
rom[43286] = 12'h666;
rom[43287] = 12'h666;
rom[43288] = 12'h666;
rom[43289] = 12'h666;
rom[43290] = 12'h777;
rom[43291] = 12'h777;
rom[43292] = 12'h777;
rom[43293] = 12'h666;
rom[43294] = 12'h555;
rom[43295] = 12'h555;
rom[43296] = 12'h444;
rom[43297] = 12'h444;
rom[43298] = 12'h444;
rom[43299] = 12'h333;
rom[43300] = 12'h333;
rom[43301] = 12'h333;
rom[43302] = 12'h333;
rom[43303] = 12'h333;
rom[43304] = 12'h333;
rom[43305] = 12'h333;
rom[43306] = 12'h333;
rom[43307] = 12'h333;
rom[43308] = 12'h222;
rom[43309] = 12'h222;
rom[43310] = 12'h222;
rom[43311] = 12'h111;
rom[43312] = 12'h111;
rom[43313] = 12'h111;
rom[43314] = 12'h  0;
rom[43315] = 12'h  0;
rom[43316] = 12'h  0;
rom[43317] = 12'h  0;
rom[43318] = 12'h  0;
rom[43319] = 12'h  0;
rom[43320] = 12'h  0;
rom[43321] = 12'h  0;
rom[43322] = 12'h  0;
rom[43323] = 12'h  0;
rom[43324] = 12'h  0;
rom[43325] = 12'h  0;
rom[43326] = 12'h  0;
rom[43327] = 12'h  0;
rom[43328] = 12'h  0;
rom[43329] = 12'h  0;
rom[43330] = 12'h  0;
rom[43331] = 12'h  0;
rom[43332] = 12'h  0;
rom[43333] = 12'h  0;
rom[43334] = 12'h  0;
rom[43335] = 12'h  0;
rom[43336] = 12'h  0;
rom[43337] = 12'h  0;
rom[43338] = 12'h  0;
rom[43339] = 12'h  0;
rom[43340] = 12'h  0;
rom[43341] = 12'h  0;
rom[43342] = 12'h  0;
rom[43343] = 12'h  0;
rom[43344] = 12'h  0;
rom[43345] = 12'h  0;
rom[43346] = 12'h  0;
rom[43347] = 12'h  0;
rom[43348] = 12'h  0;
rom[43349] = 12'h  0;
rom[43350] = 12'h  0;
rom[43351] = 12'h  0;
rom[43352] = 12'h  0;
rom[43353] = 12'h111;
rom[43354] = 12'h111;
rom[43355] = 12'h111;
rom[43356] = 12'h111;
rom[43357] = 12'h111;
rom[43358] = 12'h111;
rom[43359] = 12'h111;
rom[43360] = 12'h111;
rom[43361] = 12'h111;
rom[43362] = 12'h111;
rom[43363] = 12'h111;
rom[43364] = 12'h111;
rom[43365] = 12'h111;
rom[43366] = 12'h222;
rom[43367] = 12'h222;
rom[43368] = 12'h222;
rom[43369] = 12'h222;
rom[43370] = 12'h222;
rom[43371] = 12'h222;
rom[43372] = 12'h222;
rom[43373] = 12'h222;
rom[43374] = 12'h222;
rom[43375] = 12'h222;
rom[43376] = 12'h222;
rom[43377] = 12'h222;
rom[43378] = 12'h222;
rom[43379] = 12'h222;
rom[43380] = 12'h222;
rom[43381] = 12'h222;
rom[43382] = 12'h222;
rom[43383] = 12'h222;
rom[43384] = 12'h222;
rom[43385] = 12'h222;
rom[43386] = 12'h222;
rom[43387] = 12'h222;
rom[43388] = 12'h222;
rom[43389] = 12'h333;
rom[43390] = 12'h333;
rom[43391] = 12'h333;
rom[43392] = 12'h333;
rom[43393] = 12'h333;
rom[43394] = 12'h333;
rom[43395] = 12'h333;
rom[43396] = 12'h333;
rom[43397] = 12'h333;
rom[43398] = 12'h333;
rom[43399] = 12'h333;
rom[43400] = 12'h333;
rom[43401] = 12'h333;
rom[43402] = 12'h333;
rom[43403] = 12'h333;
rom[43404] = 12'h333;
rom[43405] = 12'h333;
rom[43406] = 12'h333;
rom[43407] = 12'h333;
rom[43408] = 12'h333;
rom[43409] = 12'h333;
rom[43410] = 12'h333;
rom[43411] = 12'h333;
rom[43412] = 12'h333;
rom[43413] = 12'h444;
rom[43414] = 12'h444;
rom[43415] = 12'h444;
rom[43416] = 12'h444;
rom[43417] = 12'h444;
rom[43418] = 12'h444;
rom[43419] = 12'h444;
rom[43420] = 12'h444;
rom[43421] = 12'h444;
rom[43422] = 12'h444;
rom[43423] = 12'h444;
rom[43424] = 12'h444;
rom[43425] = 12'h333;
rom[43426] = 12'h333;
rom[43427] = 12'h333;
rom[43428] = 12'h333;
rom[43429] = 12'h333;
rom[43430] = 12'h333;
rom[43431] = 12'h333;
rom[43432] = 12'h333;
rom[43433] = 12'h333;
rom[43434] = 12'h222;
rom[43435] = 12'h222;
rom[43436] = 12'h222;
rom[43437] = 12'h222;
rom[43438] = 12'h222;
rom[43439] = 12'h222;
rom[43440] = 12'h111;
rom[43441] = 12'h111;
rom[43442] = 12'h111;
rom[43443] = 12'h111;
rom[43444] = 12'h111;
rom[43445] = 12'h111;
rom[43446] = 12'h111;
rom[43447] = 12'h111;
rom[43448] = 12'h  0;
rom[43449] = 12'h  0;
rom[43450] = 12'h  0;
rom[43451] = 12'h  0;
rom[43452] = 12'h  0;
rom[43453] = 12'h  0;
rom[43454] = 12'h  0;
rom[43455] = 12'h  0;
rom[43456] = 12'h  0;
rom[43457] = 12'h  0;
rom[43458] = 12'h  0;
rom[43459] = 12'h  0;
rom[43460] = 12'h  0;
rom[43461] = 12'h  0;
rom[43462] = 12'h  0;
rom[43463] = 12'h  0;
rom[43464] = 12'h  0;
rom[43465] = 12'h  0;
rom[43466] = 12'h  0;
rom[43467] = 12'h  0;
rom[43468] = 12'h  0;
rom[43469] = 12'h  0;
rom[43470] = 12'h111;
rom[43471] = 12'h111;
rom[43472] = 12'h111;
rom[43473] = 12'h111;
rom[43474] = 12'h222;
rom[43475] = 12'h222;
rom[43476] = 12'h222;
rom[43477] = 12'h222;
rom[43478] = 12'h333;
rom[43479] = 12'h444;
rom[43480] = 12'h444;
rom[43481] = 12'h555;
rom[43482] = 12'h555;
rom[43483] = 12'h555;
rom[43484] = 12'h555;
rom[43485] = 12'h666;
rom[43486] = 12'h777;
rom[43487] = 12'h777;
rom[43488] = 12'h777;
rom[43489] = 12'h888;
rom[43490] = 12'h888;
rom[43491] = 12'h999;
rom[43492] = 12'haaa;
rom[43493] = 12'habb;
rom[43494] = 12'hccc;
rom[43495] = 12'hedd;
rom[43496] = 12'heee;
rom[43497] = 12'ha99;
rom[43498] = 12'h533;
rom[43499] = 12'h310;
rom[43500] = 12'h411;
rom[43501] = 12'h511;
rom[43502] = 12'h410;
rom[43503] = 12'h500;
rom[43504] = 12'h500;
rom[43505] = 12'h400;
rom[43506] = 12'h400;
rom[43507] = 12'h400;
rom[43508] = 12'h400;
rom[43509] = 12'h400;
rom[43510] = 12'h500;
rom[43511] = 12'h500;
rom[43512] = 12'h500;
rom[43513] = 12'h500;
rom[43514] = 12'h500;
rom[43515] = 12'h500;
rom[43516] = 12'h600;
rom[43517] = 12'h600;
rom[43518] = 12'h600;
rom[43519] = 12'h600;
rom[43520] = 12'h600;
rom[43521] = 12'h600;
rom[43522] = 12'h600;
rom[43523] = 12'h600;
rom[43524] = 12'h600;
rom[43525] = 12'h600;
rom[43526] = 12'h600;
rom[43527] = 12'h600;
rom[43528] = 12'h600;
rom[43529] = 12'h600;
rom[43530] = 12'h600;
rom[43531] = 12'h600;
rom[43532] = 12'h600;
rom[43533] = 12'h600;
rom[43534] = 12'h600;
rom[43535] = 12'h600;
rom[43536] = 12'h600;
rom[43537] = 12'h600;
rom[43538] = 12'h600;
rom[43539] = 12'h600;
rom[43540] = 12'h600;
rom[43541] = 12'h610;
rom[43542] = 12'h610;
rom[43543] = 12'h610;
rom[43544] = 12'h720;
rom[43545] = 12'h720;
rom[43546] = 12'h720;
rom[43547] = 12'h730;
rom[43548] = 12'h720;
rom[43549] = 12'h720;
rom[43550] = 12'h720;
rom[43551] = 12'h720;
rom[43552] = 12'h620;
rom[43553] = 12'h620;
rom[43554] = 12'h620;
rom[43555] = 12'h520;
rom[43556] = 12'h520;
rom[43557] = 12'h520;
rom[43558] = 12'h530;
rom[43559] = 12'h531;
rom[43560] = 12'h531;
rom[43561] = 12'h431;
rom[43562] = 12'h432;
rom[43563] = 12'h432;
rom[43564] = 12'h432;
rom[43565] = 12'h432;
rom[43566] = 12'h543;
rom[43567] = 12'h543;
rom[43568] = 12'h543;
rom[43569] = 12'h654;
rom[43570] = 12'h654;
rom[43571] = 12'h665;
rom[43572] = 12'h665;
rom[43573] = 12'h666;
rom[43574] = 12'h766;
rom[43575] = 12'h777;
rom[43576] = 12'h677;
rom[43577] = 12'h777;
rom[43578] = 12'h788;
rom[43579] = 12'h888;
rom[43580] = 12'h899;
rom[43581] = 12'h99a;
rom[43582] = 12'haaa;
rom[43583] = 12'haaa;
rom[43584] = 12'hbbb;
rom[43585] = 12'hbbb;
rom[43586] = 12'hbbb;
rom[43587] = 12'hbbb;
rom[43588] = 12'haaa;
rom[43589] = 12'haaa;
rom[43590] = 12'haaa;
rom[43591] = 12'haaa;
rom[43592] = 12'haaa;
rom[43593] = 12'h999;
rom[43594] = 12'h999;
rom[43595] = 12'h999;
rom[43596] = 12'haaa;
rom[43597] = 12'haaa;
rom[43598] = 12'haaa;
rom[43599] = 12'haaa;
rom[43600] = 12'h888;
rom[43601] = 12'h888;
rom[43602] = 12'h777;
rom[43603] = 12'h777;
rom[43604] = 12'h777;
rom[43605] = 12'h777;
rom[43606] = 12'h777;
rom[43607] = 12'h888;
rom[43608] = 12'h888;
rom[43609] = 12'h888;
rom[43610] = 12'h777;
rom[43611] = 12'h777;
rom[43612] = 12'h777;
rom[43613] = 12'h777;
rom[43614] = 12'h777;
rom[43615] = 12'h777;
rom[43616] = 12'h666;
rom[43617] = 12'h666;
rom[43618] = 12'h666;
rom[43619] = 12'h666;
rom[43620] = 12'h666;
rom[43621] = 12'h777;
rom[43622] = 12'h777;
rom[43623] = 12'h777;
rom[43624] = 12'h777;
rom[43625] = 12'h777;
rom[43626] = 12'h777;
rom[43627] = 12'h777;
rom[43628] = 12'h777;
rom[43629] = 12'h777;
rom[43630] = 12'h777;
rom[43631] = 12'h777;
rom[43632] = 12'h777;
rom[43633] = 12'h777;
rom[43634] = 12'h777;
rom[43635] = 12'h777;
rom[43636] = 12'h888;
rom[43637] = 12'h888;
rom[43638] = 12'h888;
rom[43639] = 12'h777;
rom[43640] = 12'h888;
rom[43641] = 12'h888;
rom[43642] = 12'h888;
rom[43643] = 12'h888;
rom[43644] = 12'h888;
rom[43645] = 12'h888;
rom[43646] = 12'h888;
rom[43647] = 12'h888;
rom[43648] = 12'h999;
rom[43649] = 12'h999;
rom[43650] = 12'h999;
rom[43651] = 12'h999;
rom[43652] = 12'h999;
rom[43653] = 12'h999;
rom[43654] = 12'haaa;
rom[43655] = 12'haaa;
rom[43656] = 12'haaa;
rom[43657] = 12'haaa;
rom[43658] = 12'hbbb;
rom[43659] = 12'hbbb;
rom[43660] = 12'hbbb;
rom[43661] = 12'hbbb;
rom[43662] = 12'haaa;
rom[43663] = 12'haaa;
rom[43664] = 12'h999;
rom[43665] = 12'h999;
rom[43666] = 12'h999;
rom[43667] = 12'h888;
rom[43668] = 12'h888;
rom[43669] = 12'h888;
rom[43670] = 12'h888;
rom[43671] = 12'h888;
rom[43672] = 12'h777;
rom[43673] = 12'h777;
rom[43674] = 12'h777;
rom[43675] = 12'h666;
rom[43676] = 12'h666;
rom[43677] = 12'h666;
rom[43678] = 12'h666;
rom[43679] = 12'h666;
rom[43680] = 12'h666;
rom[43681] = 12'h666;
rom[43682] = 12'h666;
rom[43683] = 12'h666;
rom[43684] = 12'h555;
rom[43685] = 12'h555;
rom[43686] = 12'h555;
rom[43687] = 12'h555;
rom[43688] = 12'h666;
rom[43689] = 12'h666;
rom[43690] = 12'h666;
rom[43691] = 12'h777;
rom[43692] = 12'h777;
rom[43693] = 12'h666;
rom[43694] = 12'h666;
rom[43695] = 12'h555;
rom[43696] = 12'h555;
rom[43697] = 12'h444;
rom[43698] = 12'h444;
rom[43699] = 12'h444;
rom[43700] = 12'h333;
rom[43701] = 12'h333;
rom[43702] = 12'h333;
rom[43703] = 12'h333;
rom[43704] = 12'h333;
rom[43705] = 12'h333;
rom[43706] = 12'h333;
rom[43707] = 12'h333;
rom[43708] = 12'h222;
rom[43709] = 12'h222;
rom[43710] = 12'h222;
rom[43711] = 12'h222;
rom[43712] = 12'h222;
rom[43713] = 12'h111;
rom[43714] = 12'h111;
rom[43715] = 12'h  0;
rom[43716] = 12'h  0;
rom[43717] = 12'h  0;
rom[43718] = 12'h  0;
rom[43719] = 12'h  0;
rom[43720] = 12'h  0;
rom[43721] = 12'h  0;
rom[43722] = 12'h  0;
rom[43723] = 12'h  0;
rom[43724] = 12'h  0;
rom[43725] = 12'h  0;
rom[43726] = 12'h  0;
rom[43727] = 12'h  0;
rom[43728] = 12'h  0;
rom[43729] = 12'h  0;
rom[43730] = 12'h  0;
rom[43731] = 12'h  0;
rom[43732] = 12'h  0;
rom[43733] = 12'h  0;
rom[43734] = 12'h  0;
rom[43735] = 12'h  0;
rom[43736] = 12'h  0;
rom[43737] = 12'h  0;
rom[43738] = 12'h  0;
rom[43739] = 12'h  0;
rom[43740] = 12'h  0;
rom[43741] = 12'h  0;
rom[43742] = 12'h  0;
rom[43743] = 12'h  0;
rom[43744] = 12'h111;
rom[43745] = 12'h111;
rom[43746] = 12'h111;
rom[43747] = 12'h111;
rom[43748] = 12'h111;
rom[43749] = 12'h111;
rom[43750] = 12'h111;
rom[43751] = 12'h111;
rom[43752] = 12'h111;
rom[43753] = 12'h111;
rom[43754] = 12'h111;
rom[43755] = 12'h111;
rom[43756] = 12'h111;
rom[43757] = 12'h111;
rom[43758] = 12'h111;
rom[43759] = 12'h111;
rom[43760] = 12'h111;
rom[43761] = 12'h111;
rom[43762] = 12'h111;
rom[43763] = 12'h111;
rom[43764] = 12'h222;
rom[43765] = 12'h222;
rom[43766] = 12'h222;
rom[43767] = 12'h222;
rom[43768] = 12'h222;
rom[43769] = 12'h222;
rom[43770] = 12'h222;
rom[43771] = 12'h222;
rom[43772] = 12'h222;
rom[43773] = 12'h222;
rom[43774] = 12'h222;
rom[43775] = 12'h222;
rom[43776] = 12'h222;
rom[43777] = 12'h222;
rom[43778] = 12'h222;
rom[43779] = 12'h222;
rom[43780] = 12'h222;
rom[43781] = 12'h222;
rom[43782] = 12'h222;
rom[43783] = 12'h222;
rom[43784] = 12'h222;
rom[43785] = 12'h222;
rom[43786] = 12'h222;
rom[43787] = 12'h222;
rom[43788] = 12'h222;
rom[43789] = 12'h222;
rom[43790] = 12'h333;
rom[43791] = 12'h333;
rom[43792] = 12'h333;
rom[43793] = 12'h333;
rom[43794] = 12'h333;
rom[43795] = 12'h333;
rom[43796] = 12'h333;
rom[43797] = 12'h333;
rom[43798] = 12'h333;
rom[43799] = 12'h333;
rom[43800] = 12'h333;
rom[43801] = 12'h333;
rom[43802] = 12'h333;
rom[43803] = 12'h333;
rom[43804] = 12'h222;
rom[43805] = 12'h222;
rom[43806] = 12'h222;
rom[43807] = 12'h222;
rom[43808] = 12'h333;
rom[43809] = 12'h333;
rom[43810] = 12'h333;
rom[43811] = 12'h333;
rom[43812] = 12'h333;
rom[43813] = 12'h333;
rom[43814] = 12'h333;
rom[43815] = 12'h333;
rom[43816] = 12'h333;
rom[43817] = 12'h333;
rom[43818] = 12'h333;
rom[43819] = 12'h333;
rom[43820] = 12'h333;
rom[43821] = 12'h333;
rom[43822] = 12'h333;
rom[43823] = 12'h333;
rom[43824] = 12'h333;
rom[43825] = 12'h333;
rom[43826] = 12'h333;
rom[43827] = 12'h333;
rom[43828] = 12'h333;
rom[43829] = 12'h333;
rom[43830] = 12'h333;
rom[43831] = 12'h333;
rom[43832] = 12'h333;
rom[43833] = 12'h222;
rom[43834] = 12'h222;
rom[43835] = 12'h222;
rom[43836] = 12'h222;
rom[43837] = 12'h222;
rom[43838] = 12'h222;
rom[43839] = 12'h222;
rom[43840] = 12'h111;
rom[43841] = 12'h111;
rom[43842] = 12'h111;
rom[43843] = 12'h111;
rom[43844] = 12'h111;
rom[43845] = 12'h111;
rom[43846] = 12'h111;
rom[43847] = 12'h111;
rom[43848] = 12'h  0;
rom[43849] = 12'h  0;
rom[43850] = 12'h  0;
rom[43851] = 12'h  0;
rom[43852] = 12'h  0;
rom[43853] = 12'h  0;
rom[43854] = 12'h  0;
rom[43855] = 12'h  0;
rom[43856] = 12'h  0;
rom[43857] = 12'h  0;
rom[43858] = 12'h  0;
rom[43859] = 12'h  0;
rom[43860] = 12'h  0;
rom[43861] = 12'h  0;
rom[43862] = 12'h  0;
rom[43863] = 12'h  0;
rom[43864] = 12'h  0;
rom[43865] = 12'h  0;
rom[43866] = 12'h  0;
rom[43867] = 12'h  0;
rom[43868] = 12'h  0;
rom[43869] = 12'h  0;
rom[43870] = 12'h111;
rom[43871] = 12'h111;
rom[43872] = 12'h111;
rom[43873] = 12'h111;
rom[43874] = 12'h222;
rom[43875] = 12'h222;
rom[43876] = 12'h222;
rom[43877] = 12'h222;
rom[43878] = 12'h333;
rom[43879] = 12'h444;
rom[43880] = 12'h444;
rom[43881] = 12'h555;
rom[43882] = 12'h555;
rom[43883] = 12'h555;
rom[43884] = 12'h666;
rom[43885] = 12'h666;
rom[43886] = 12'h666;
rom[43887] = 12'h777;
rom[43888] = 12'h777;
rom[43889] = 12'h888;
rom[43890] = 12'h888;
rom[43891] = 12'h999;
rom[43892] = 12'haaa;
rom[43893] = 12'hbbb;
rom[43894] = 12'hccc;
rom[43895] = 12'hddd;
rom[43896] = 12'hddd;
rom[43897] = 12'h887;
rom[43898] = 12'h422;
rom[43899] = 12'h311;
rom[43900] = 12'h411;
rom[43901] = 12'h410;
rom[43902] = 12'h410;
rom[43903] = 12'h400;
rom[43904] = 12'h400;
rom[43905] = 12'h400;
rom[43906] = 12'h400;
rom[43907] = 12'h400;
rom[43908] = 12'h400;
rom[43909] = 12'h400;
rom[43910] = 12'h400;
rom[43911] = 12'h400;
rom[43912] = 12'h400;
rom[43913] = 12'h400;
rom[43914] = 12'h500;
rom[43915] = 12'h500;
rom[43916] = 12'h500;
rom[43917] = 12'h500;
rom[43918] = 12'h500;
rom[43919] = 12'h500;
rom[43920] = 12'h500;
rom[43921] = 12'h500;
rom[43922] = 12'h500;
rom[43923] = 12'h500;
rom[43924] = 12'h500;
rom[43925] = 12'h500;
rom[43926] = 12'h600;
rom[43927] = 12'h600;
rom[43928] = 12'h600;
rom[43929] = 12'h500;
rom[43930] = 12'h500;
rom[43931] = 12'h500;
rom[43932] = 12'h500;
rom[43933] = 12'h500;
rom[43934] = 12'h500;
rom[43935] = 12'h500;
rom[43936] = 12'h500;
rom[43937] = 12'h500;
rom[43938] = 12'h500;
rom[43939] = 12'h500;
rom[43940] = 12'h500;
rom[43941] = 12'h510;
rom[43942] = 12'h610;
rom[43943] = 12'h610;
rom[43944] = 12'h620;
rom[43945] = 12'h620;
rom[43946] = 12'h720;
rom[43947] = 12'h720;
rom[43948] = 12'h720;
rom[43949] = 12'h720;
rom[43950] = 12'h720;
rom[43951] = 12'h720;
rom[43952] = 12'h620;
rom[43953] = 12'h620;
rom[43954] = 12'h620;
rom[43955] = 12'h520;
rom[43956] = 12'h520;
rom[43957] = 12'h520;
rom[43958] = 12'h530;
rom[43959] = 12'h531;
rom[43960] = 12'h531;
rom[43961] = 12'h531;
rom[43962] = 12'h532;
rom[43963] = 12'h532;
rom[43964] = 12'h543;
rom[43965] = 12'h543;
rom[43966] = 12'h544;
rom[43967] = 12'h644;
rom[43968] = 12'h654;
rom[43969] = 12'h654;
rom[43970] = 12'h665;
rom[43971] = 12'h765;
rom[43972] = 12'h766;
rom[43973] = 12'h766;
rom[43974] = 12'h777;
rom[43975] = 12'h777;
rom[43976] = 12'h777;
rom[43977] = 12'h778;
rom[43978] = 12'h888;
rom[43979] = 12'h889;
rom[43980] = 12'h999;
rom[43981] = 12'h9aa;
rom[43982] = 12'haab;
rom[43983] = 12'habb;
rom[43984] = 12'hbbb;
rom[43985] = 12'hbbb;
rom[43986] = 12'hbbb;
rom[43987] = 12'hbbb;
rom[43988] = 12'haaa;
rom[43989] = 12'haaa;
rom[43990] = 12'haaa;
rom[43991] = 12'haaa;
rom[43992] = 12'h999;
rom[43993] = 12'h999;
rom[43994] = 12'h999;
rom[43995] = 12'h999;
rom[43996] = 12'haaa;
rom[43997] = 12'haaa;
rom[43998] = 12'haaa;
rom[43999] = 12'haaa;
rom[44000] = 12'h888;
rom[44001] = 12'h888;
rom[44002] = 12'h888;
rom[44003] = 12'h777;
rom[44004] = 12'h777;
rom[44005] = 12'h888;
rom[44006] = 12'h888;
rom[44007] = 12'h888;
rom[44008] = 12'h888;
rom[44009] = 12'h777;
rom[44010] = 12'h777;
rom[44011] = 12'h777;
rom[44012] = 12'h777;
rom[44013] = 12'h777;
rom[44014] = 12'h666;
rom[44015] = 12'h666;
rom[44016] = 12'h666;
rom[44017] = 12'h666;
rom[44018] = 12'h666;
rom[44019] = 12'h777;
rom[44020] = 12'h777;
rom[44021] = 12'h777;
rom[44022] = 12'h777;
rom[44023] = 12'h777;
rom[44024] = 12'h777;
rom[44025] = 12'h777;
rom[44026] = 12'h777;
rom[44027] = 12'h777;
rom[44028] = 12'h777;
rom[44029] = 12'h777;
rom[44030] = 12'h777;
rom[44031] = 12'h777;
rom[44032] = 12'h777;
rom[44033] = 12'h777;
rom[44034] = 12'h777;
rom[44035] = 12'h777;
rom[44036] = 12'h777;
rom[44037] = 12'h777;
rom[44038] = 12'h777;
rom[44039] = 12'h777;
rom[44040] = 12'h888;
rom[44041] = 12'h888;
rom[44042] = 12'h888;
rom[44043] = 12'h888;
rom[44044] = 12'h888;
rom[44045] = 12'h888;
rom[44046] = 12'h888;
rom[44047] = 12'h888;
rom[44048] = 12'h888;
rom[44049] = 12'h888;
rom[44050] = 12'h999;
rom[44051] = 12'h999;
rom[44052] = 12'h999;
rom[44053] = 12'h999;
rom[44054] = 12'h999;
rom[44055] = 12'haaa;
rom[44056] = 12'haaa;
rom[44057] = 12'haaa;
rom[44058] = 12'haaa;
rom[44059] = 12'hbbb;
rom[44060] = 12'hbbb;
rom[44061] = 12'haaa;
rom[44062] = 12'haaa;
rom[44063] = 12'haaa;
rom[44064] = 12'haaa;
rom[44065] = 12'h999;
rom[44066] = 12'h999;
rom[44067] = 12'h888;
rom[44068] = 12'h888;
rom[44069] = 12'h888;
rom[44070] = 12'h888;
rom[44071] = 12'h888;
rom[44072] = 12'h777;
rom[44073] = 12'h777;
rom[44074] = 12'h777;
rom[44075] = 12'h666;
rom[44076] = 12'h666;
rom[44077] = 12'h666;
rom[44078] = 12'h666;
rom[44079] = 12'h666;
rom[44080] = 12'h666;
rom[44081] = 12'h666;
rom[44082] = 12'h666;
rom[44083] = 12'h555;
rom[44084] = 12'h555;
rom[44085] = 12'h555;
rom[44086] = 12'h555;
rom[44087] = 12'h555;
rom[44088] = 12'h555;
rom[44089] = 12'h666;
rom[44090] = 12'h666;
rom[44091] = 12'h777;
rom[44092] = 12'h777;
rom[44093] = 12'h666;
rom[44094] = 12'h666;
rom[44095] = 12'h666;
rom[44096] = 12'h555;
rom[44097] = 12'h555;
rom[44098] = 12'h444;
rom[44099] = 12'h444;
rom[44100] = 12'h444;
rom[44101] = 12'h333;
rom[44102] = 12'h333;
rom[44103] = 12'h333;
rom[44104] = 12'h333;
rom[44105] = 12'h333;
rom[44106] = 12'h333;
rom[44107] = 12'h333;
rom[44108] = 12'h222;
rom[44109] = 12'h222;
rom[44110] = 12'h222;
rom[44111] = 12'h111;
rom[44112] = 12'h222;
rom[44113] = 12'h111;
rom[44114] = 12'h111;
rom[44115] = 12'h111;
rom[44116] = 12'h  0;
rom[44117] = 12'h  0;
rom[44118] = 12'h  0;
rom[44119] = 12'h  0;
rom[44120] = 12'h  0;
rom[44121] = 12'h  0;
rom[44122] = 12'h  0;
rom[44123] = 12'h  0;
rom[44124] = 12'h  0;
rom[44125] = 12'h  0;
rom[44126] = 12'h  0;
rom[44127] = 12'h  0;
rom[44128] = 12'h  0;
rom[44129] = 12'h  0;
rom[44130] = 12'h  0;
rom[44131] = 12'h  0;
rom[44132] = 12'h  0;
rom[44133] = 12'h  0;
rom[44134] = 12'h  0;
rom[44135] = 12'h  0;
rom[44136] = 12'h  0;
rom[44137] = 12'h  0;
rom[44138] = 12'h  0;
rom[44139] = 12'h  0;
rom[44140] = 12'h  0;
rom[44141] = 12'h  0;
rom[44142] = 12'h  0;
rom[44143] = 12'h111;
rom[44144] = 12'h111;
rom[44145] = 12'h111;
rom[44146] = 12'h111;
rom[44147] = 12'h111;
rom[44148] = 12'h111;
rom[44149] = 12'h111;
rom[44150] = 12'h111;
rom[44151] = 12'h111;
rom[44152] = 12'h111;
rom[44153] = 12'h111;
rom[44154] = 12'h111;
rom[44155] = 12'h111;
rom[44156] = 12'h111;
rom[44157] = 12'h111;
rom[44158] = 12'h111;
rom[44159] = 12'h111;
rom[44160] = 12'h111;
rom[44161] = 12'h111;
rom[44162] = 12'h222;
rom[44163] = 12'h222;
rom[44164] = 12'h222;
rom[44165] = 12'h222;
rom[44166] = 12'h222;
rom[44167] = 12'h222;
rom[44168] = 12'h222;
rom[44169] = 12'h222;
rom[44170] = 12'h222;
rom[44171] = 12'h222;
rom[44172] = 12'h222;
rom[44173] = 12'h222;
rom[44174] = 12'h222;
rom[44175] = 12'h222;
rom[44176] = 12'h222;
rom[44177] = 12'h222;
rom[44178] = 12'h222;
rom[44179] = 12'h222;
rom[44180] = 12'h222;
rom[44181] = 12'h222;
rom[44182] = 12'h222;
rom[44183] = 12'h222;
rom[44184] = 12'h222;
rom[44185] = 12'h222;
rom[44186] = 12'h222;
rom[44187] = 12'h222;
rom[44188] = 12'h222;
rom[44189] = 12'h222;
rom[44190] = 12'h333;
rom[44191] = 12'h333;
rom[44192] = 12'h333;
rom[44193] = 12'h333;
rom[44194] = 12'h333;
rom[44195] = 12'h333;
rom[44196] = 12'h333;
rom[44197] = 12'h333;
rom[44198] = 12'h333;
rom[44199] = 12'h222;
rom[44200] = 12'h222;
rom[44201] = 12'h222;
rom[44202] = 12'h222;
rom[44203] = 12'h222;
rom[44204] = 12'h222;
rom[44205] = 12'h222;
rom[44206] = 12'h222;
rom[44207] = 12'h222;
rom[44208] = 12'h222;
rom[44209] = 12'h222;
rom[44210] = 12'h222;
rom[44211] = 12'h333;
rom[44212] = 12'h333;
rom[44213] = 12'h333;
rom[44214] = 12'h333;
rom[44215] = 12'h333;
rom[44216] = 12'h333;
rom[44217] = 12'h333;
rom[44218] = 12'h333;
rom[44219] = 12'h333;
rom[44220] = 12'h333;
rom[44221] = 12'h333;
rom[44222] = 12'h333;
rom[44223] = 12'h333;
rom[44224] = 12'h333;
rom[44225] = 12'h333;
rom[44226] = 12'h333;
rom[44227] = 12'h333;
rom[44228] = 12'h333;
rom[44229] = 12'h333;
rom[44230] = 12'h333;
rom[44231] = 12'h333;
rom[44232] = 12'h333;
rom[44233] = 12'h222;
rom[44234] = 12'h222;
rom[44235] = 12'h222;
rom[44236] = 12'h222;
rom[44237] = 12'h222;
rom[44238] = 12'h222;
rom[44239] = 12'h111;
rom[44240] = 12'h111;
rom[44241] = 12'h111;
rom[44242] = 12'h111;
rom[44243] = 12'h111;
rom[44244] = 12'h111;
rom[44245] = 12'h111;
rom[44246] = 12'h111;
rom[44247] = 12'h111;
rom[44248] = 12'h111;
rom[44249] = 12'h  0;
rom[44250] = 12'h  0;
rom[44251] = 12'h  0;
rom[44252] = 12'h  0;
rom[44253] = 12'h  0;
rom[44254] = 12'h  0;
rom[44255] = 12'h  0;
rom[44256] = 12'h  0;
rom[44257] = 12'h  0;
rom[44258] = 12'h  0;
rom[44259] = 12'h  0;
rom[44260] = 12'h  0;
rom[44261] = 12'h  0;
rom[44262] = 12'h  0;
rom[44263] = 12'h  0;
rom[44264] = 12'h  0;
rom[44265] = 12'h  0;
rom[44266] = 12'h  0;
rom[44267] = 12'h  0;
rom[44268] = 12'h  0;
rom[44269] = 12'h  0;
rom[44270] = 12'h  0;
rom[44271] = 12'h111;
rom[44272] = 12'h111;
rom[44273] = 12'h111;
rom[44274] = 12'h222;
rom[44275] = 12'h222;
rom[44276] = 12'h222;
rom[44277] = 12'h333;
rom[44278] = 12'h333;
rom[44279] = 12'h444;
rom[44280] = 12'h444;
rom[44281] = 12'h555;
rom[44282] = 12'h555;
rom[44283] = 12'h555;
rom[44284] = 12'h666;
rom[44285] = 12'h666;
rom[44286] = 12'h666;
rom[44287] = 12'h777;
rom[44288] = 12'h777;
rom[44289] = 12'h888;
rom[44290] = 12'h888;
rom[44291] = 12'h999;
rom[44292] = 12'haaa;
rom[44293] = 12'hbcb;
rom[44294] = 12'hccc;
rom[44295] = 12'hddd;
rom[44296] = 12'hccc;
rom[44297] = 12'h776;
rom[44298] = 12'h322;
rom[44299] = 12'h310;
rom[44300] = 12'h410;
rom[44301] = 12'h410;
rom[44302] = 12'h400;
rom[44303] = 12'h400;
rom[44304] = 12'h300;
rom[44305] = 12'h300;
rom[44306] = 12'h300;
rom[44307] = 12'h300;
rom[44308] = 12'h300;
rom[44309] = 12'h300;
rom[44310] = 12'h300;
rom[44311] = 12'h300;
rom[44312] = 12'h400;
rom[44313] = 12'h400;
rom[44314] = 12'h400;
rom[44315] = 12'h400;
rom[44316] = 12'h400;
rom[44317] = 12'h500;
rom[44318] = 12'h500;
rom[44319] = 12'h500;
rom[44320] = 12'h500;
rom[44321] = 12'h500;
rom[44322] = 12'h500;
rom[44323] = 12'h500;
rom[44324] = 12'h500;
rom[44325] = 12'h500;
rom[44326] = 12'h500;
rom[44327] = 12'h500;
rom[44328] = 12'h500;
rom[44329] = 12'h500;
rom[44330] = 12'h500;
rom[44331] = 12'h500;
rom[44332] = 12'h400;
rom[44333] = 12'h400;
rom[44334] = 12'h400;
rom[44335] = 12'h400;
rom[44336] = 12'h400;
rom[44337] = 12'h500;
rom[44338] = 12'h400;
rom[44339] = 12'h500;
rom[44340] = 12'h500;
rom[44341] = 12'h500;
rom[44342] = 12'h510;
rom[44343] = 12'h510;
rom[44344] = 12'h610;
rom[44345] = 12'h620;
rom[44346] = 12'h620;
rom[44347] = 12'h620;
rom[44348] = 12'h620;
rom[44349] = 12'h620;
rom[44350] = 12'h720;
rom[44351] = 12'h620;
rom[44352] = 12'h620;
rom[44353] = 12'h620;
rom[44354] = 12'h620;
rom[44355] = 12'h520;
rom[44356] = 12'h520;
rom[44357] = 12'h520;
rom[44358] = 12'h530;
rom[44359] = 12'h531;
rom[44360] = 12'h531;
rom[44361] = 12'h532;
rom[44362] = 12'h542;
rom[44363] = 12'h542;
rom[44364] = 12'h543;
rom[44365] = 12'h544;
rom[44366] = 12'h644;
rom[44367] = 12'h655;
rom[44368] = 12'h655;
rom[44369] = 12'h665;
rom[44370] = 12'h765;
rom[44371] = 12'h766;
rom[44372] = 12'h766;
rom[44373] = 12'h776;
rom[44374] = 12'h777;
rom[44375] = 12'h777;
rom[44376] = 12'h777;
rom[44377] = 12'h788;
rom[44378] = 12'h889;
rom[44379] = 12'h999;
rom[44380] = 12'h9aa;
rom[44381] = 12'haaa;
rom[44382] = 12'habb;
rom[44383] = 12'hbbb;
rom[44384] = 12'hbbb;
rom[44385] = 12'hbbb;
rom[44386] = 12'hbbb;
rom[44387] = 12'hbbb;
rom[44388] = 12'haaa;
rom[44389] = 12'haaa;
rom[44390] = 12'haaa;
rom[44391] = 12'haaa;
rom[44392] = 12'h999;
rom[44393] = 12'h999;
rom[44394] = 12'h999;
rom[44395] = 12'h999;
rom[44396] = 12'haaa;
rom[44397] = 12'haaa;
rom[44398] = 12'haaa;
rom[44399] = 12'haaa;
rom[44400] = 12'h888;
rom[44401] = 12'h888;
rom[44402] = 12'h888;
rom[44403] = 12'h888;
rom[44404] = 12'h777;
rom[44405] = 12'h777;
rom[44406] = 12'h777;
rom[44407] = 12'h777;
rom[44408] = 12'h777;
rom[44409] = 12'h777;
rom[44410] = 12'h777;
rom[44411] = 12'h777;
rom[44412] = 12'h777;
rom[44413] = 12'h666;
rom[44414] = 12'h666;
rom[44415] = 12'h666;
rom[44416] = 12'h666;
rom[44417] = 12'h666;
rom[44418] = 12'h777;
rom[44419] = 12'h777;
rom[44420] = 12'h777;
rom[44421] = 12'h777;
rom[44422] = 12'h777;
rom[44423] = 12'h777;
rom[44424] = 12'h777;
rom[44425] = 12'h777;
rom[44426] = 12'h777;
rom[44427] = 12'h777;
rom[44428] = 12'h777;
rom[44429] = 12'h777;
rom[44430] = 12'h777;
rom[44431] = 12'h777;
rom[44432] = 12'h777;
rom[44433] = 12'h777;
rom[44434] = 12'h777;
rom[44435] = 12'h777;
rom[44436] = 12'h777;
rom[44437] = 12'h888;
rom[44438] = 12'h777;
rom[44439] = 12'h777;
rom[44440] = 12'h888;
rom[44441] = 12'h888;
rom[44442] = 12'h888;
rom[44443] = 12'h888;
rom[44444] = 12'h888;
rom[44445] = 12'h888;
rom[44446] = 12'h888;
rom[44447] = 12'h888;
rom[44448] = 12'h888;
rom[44449] = 12'h888;
rom[44450] = 12'h888;
rom[44451] = 12'h888;
rom[44452] = 12'h888;
rom[44453] = 12'h999;
rom[44454] = 12'h999;
rom[44455] = 12'h999;
rom[44456] = 12'haaa;
rom[44457] = 12'haaa;
rom[44458] = 12'haaa;
rom[44459] = 12'haaa;
rom[44460] = 12'hbbb;
rom[44461] = 12'haaa;
rom[44462] = 12'haaa;
rom[44463] = 12'haaa;
rom[44464] = 12'haaa;
rom[44465] = 12'h999;
rom[44466] = 12'h999;
rom[44467] = 12'h888;
rom[44468] = 12'h888;
rom[44469] = 12'h888;
rom[44470] = 12'h888;
rom[44471] = 12'h777;
rom[44472] = 12'h777;
rom[44473] = 12'h777;
rom[44474] = 12'h777;
rom[44475] = 12'h666;
rom[44476] = 12'h666;
rom[44477] = 12'h666;
rom[44478] = 12'h666;
rom[44479] = 12'h666;
rom[44480] = 12'h555;
rom[44481] = 12'h555;
rom[44482] = 12'h555;
rom[44483] = 12'h555;
rom[44484] = 12'h555;
rom[44485] = 12'h555;
rom[44486] = 12'h555;
rom[44487] = 12'h555;
rom[44488] = 12'h555;
rom[44489] = 12'h555;
rom[44490] = 12'h666;
rom[44491] = 12'h666;
rom[44492] = 12'h777;
rom[44493] = 12'h666;
rom[44494] = 12'h666;
rom[44495] = 12'h666;
rom[44496] = 12'h555;
rom[44497] = 12'h555;
rom[44498] = 12'h555;
rom[44499] = 12'h444;
rom[44500] = 12'h444;
rom[44501] = 12'h444;
rom[44502] = 12'h333;
rom[44503] = 12'h333;
rom[44504] = 12'h222;
rom[44505] = 12'h333;
rom[44506] = 12'h333;
rom[44507] = 12'h333;
rom[44508] = 12'h333;
rom[44509] = 12'h222;
rom[44510] = 12'h111;
rom[44511] = 12'h111;
rom[44512] = 12'h111;
rom[44513] = 12'h111;
rom[44514] = 12'h111;
rom[44515] = 12'h111;
rom[44516] = 12'h111;
rom[44517] = 12'h111;
rom[44518] = 12'h  0;
rom[44519] = 12'h  0;
rom[44520] = 12'h  0;
rom[44521] = 12'h  0;
rom[44522] = 12'h  0;
rom[44523] = 12'h  0;
rom[44524] = 12'h  0;
rom[44525] = 12'h  0;
rom[44526] = 12'h  0;
rom[44527] = 12'h  0;
rom[44528] = 12'h  0;
rom[44529] = 12'h  0;
rom[44530] = 12'h  0;
rom[44531] = 12'h  0;
rom[44532] = 12'h  0;
rom[44533] = 12'h  0;
rom[44534] = 12'h  0;
rom[44535] = 12'h  0;
rom[44536] = 12'h  0;
rom[44537] = 12'h  0;
rom[44538] = 12'h  0;
rom[44539] = 12'h  0;
rom[44540] = 12'h  0;
rom[44541] = 12'h111;
rom[44542] = 12'h111;
rom[44543] = 12'h111;
rom[44544] = 12'h111;
rom[44545] = 12'h111;
rom[44546] = 12'h111;
rom[44547] = 12'h111;
rom[44548] = 12'h111;
rom[44549] = 12'h111;
rom[44550] = 12'h111;
rom[44551] = 12'h111;
rom[44552] = 12'h111;
rom[44553] = 12'h111;
rom[44554] = 12'h111;
rom[44555] = 12'h111;
rom[44556] = 12'h111;
rom[44557] = 12'h111;
rom[44558] = 12'h111;
rom[44559] = 12'h111;
rom[44560] = 12'h111;
rom[44561] = 12'h111;
rom[44562] = 12'h111;
rom[44563] = 12'h111;
rom[44564] = 12'h222;
rom[44565] = 12'h222;
rom[44566] = 12'h222;
rom[44567] = 12'h222;
rom[44568] = 12'h222;
rom[44569] = 12'h222;
rom[44570] = 12'h222;
rom[44571] = 12'h222;
rom[44572] = 12'h111;
rom[44573] = 12'h222;
rom[44574] = 12'h222;
rom[44575] = 12'h222;
rom[44576] = 12'h222;
rom[44577] = 12'h222;
rom[44578] = 12'h222;
rom[44579] = 12'h222;
rom[44580] = 12'h222;
rom[44581] = 12'h222;
rom[44582] = 12'h222;
rom[44583] = 12'h222;
rom[44584] = 12'h222;
rom[44585] = 12'h222;
rom[44586] = 12'h222;
rom[44587] = 12'h222;
rom[44588] = 12'h222;
rom[44589] = 12'h222;
rom[44590] = 12'h333;
rom[44591] = 12'h333;
rom[44592] = 12'h333;
rom[44593] = 12'h333;
rom[44594] = 12'h333;
rom[44595] = 12'h333;
rom[44596] = 12'h222;
rom[44597] = 12'h222;
rom[44598] = 12'h222;
rom[44599] = 12'h222;
rom[44600] = 12'h222;
rom[44601] = 12'h222;
rom[44602] = 12'h222;
rom[44603] = 12'h222;
rom[44604] = 12'h222;
rom[44605] = 12'h222;
rom[44606] = 12'h222;
rom[44607] = 12'h222;
rom[44608] = 12'h222;
rom[44609] = 12'h222;
rom[44610] = 12'h222;
rom[44611] = 12'h222;
rom[44612] = 12'h333;
rom[44613] = 12'h333;
rom[44614] = 12'h333;
rom[44615] = 12'h333;
rom[44616] = 12'h333;
rom[44617] = 12'h333;
rom[44618] = 12'h333;
rom[44619] = 12'h333;
rom[44620] = 12'h333;
rom[44621] = 12'h333;
rom[44622] = 12'h333;
rom[44623] = 12'h333;
rom[44624] = 12'h333;
rom[44625] = 12'h333;
rom[44626] = 12'h333;
rom[44627] = 12'h333;
rom[44628] = 12'h333;
rom[44629] = 12'h333;
rom[44630] = 12'h333;
rom[44631] = 12'h222;
rom[44632] = 12'h222;
rom[44633] = 12'h222;
rom[44634] = 12'h222;
rom[44635] = 12'h222;
rom[44636] = 12'h222;
rom[44637] = 12'h222;
rom[44638] = 12'h111;
rom[44639] = 12'h111;
rom[44640] = 12'h111;
rom[44641] = 12'h111;
rom[44642] = 12'h111;
rom[44643] = 12'h111;
rom[44644] = 12'h111;
rom[44645] = 12'h111;
rom[44646] = 12'h111;
rom[44647] = 12'h111;
rom[44648] = 12'h111;
rom[44649] = 12'h111;
rom[44650] = 12'h  0;
rom[44651] = 12'h  0;
rom[44652] = 12'h  0;
rom[44653] = 12'h  0;
rom[44654] = 12'h  0;
rom[44655] = 12'h  0;
rom[44656] = 12'h  0;
rom[44657] = 12'h  0;
rom[44658] = 12'h  0;
rom[44659] = 12'h  0;
rom[44660] = 12'h  0;
rom[44661] = 12'h  0;
rom[44662] = 12'h  0;
rom[44663] = 12'h  0;
rom[44664] = 12'h  0;
rom[44665] = 12'h  0;
rom[44666] = 12'h  0;
rom[44667] = 12'h  0;
rom[44668] = 12'h  0;
rom[44669] = 12'h  0;
rom[44670] = 12'h  0;
rom[44671] = 12'h  0;
rom[44672] = 12'h111;
rom[44673] = 12'h111;
rom[44674] = 12'h222;
rom[44675] = 12'h222;
rom[44676] = 12'h333;
rom[44677] = 12'h333;
rom[44678] = 12'h444;
rom[44679] = 12'h444;
rom[44680] = 12'h444;
rom[44681] = 12'h555;
rom[44682] = 12'h555;
rom[44683] = 12'h666;
rom[44684] = 12'h666;
rom[44685] = 12'h666;
rom[44686] = 12'h666;
rom[44687] = 12'h777;
rom[44688] = 12'h777;
rom[44689] = 12'h888;
rom[44690] = 12'h888;
rom[44691] = 12'h899;
rom[44692] = 12'haaa;
rom[44693] = 12'hbcc;
rom[44694] = 12'hccc;
rom[44695] = 12'hddd;
rom[44696] = 12'hbbb;
rom[44697] = 12'h766;
rom[44698] = 12'h321;
rom[44699] = 12'h210;
rom[44700] = 12'h300;
rom[44701] = 12'h300;
rom[44702] = 12'h300;
rom[44703] = 12'h300;
rom[44704] = 12'h300;
rom[44705] = 12'h300;
rom[44706] = 12'h300;
rom[44707] = 12'h300;
rom[44708] = 12'h300;
rom[44709] = 12'h300;
rom[44710] = 12'h300;
rom[44711] = 12'h300;
rom[44712] = 12'h300;
rom[44713] = 12'h300;
rom[44714] = 12'h300;
rom[44715] = 12'h400;
rom[44716] = 12'h400;
rom[44717] = 12'h400;
rom[44718] = 12'h400;
rom[44719] = 12'h400;
rom[44720] = 12'h400;
rom[44721] = 12'h400;
rom[44722] = 12'h400;
rom[44723] = 12'h400;
rom[44724] = 12'h400;
rom[44725] = 12'h400;
rom[44726] = 12'h400;
rom[44727] = 12'h400;
rom[44728] = 12'h400;
rom[44729] = 12'h400;
rom[44730] = 12'h400;
rom[44731] = 12'h400;
rom[44732] = 12'h400;
rom[44733] = 12'h400;
rom[44734] = 12'h400;
rom[44735] = 12'h400;
rom[44736] = 12'h400;
rom[44737] = 12'h400;
rom[44738] = 12'h400;
rom[44739] = 12'h400;
rom[44740] = 12'h400;
rom[44741] = 12'h500;
rom[44742] = 12'h510;
rom[44743] = 12'h510;
rom[44744] = 12'h510;
rom[44745] = 12'h610;
rom[44746] = 12'h620;
rom[44747] = 12'h620;
rom[44748] = 12'h620;
rom[44749] = 12'h620;
rom[44750] = 12'h620;
rom[44751] = 12'h620;
rom[44752] = 12'h620;
rom[44753] = 12'h520;
rom[44754] = 12'h520;
rom[44755] = 12'h520;
rom[44756] = 12'h520;
rom[44757] = 12'h520;
rom[44758] = 12'h531;
rom[44759] = 12'h531;
rom[44760] = 12'h532;
rom[44761] = 12'h532;
rom[44762] = 12'h542;
rom[44763] = 12'h543;
rom[44764] = 12'h543;
rom[44765] = 12'h544;
rom[44766] = 12'h654;
rom[44767] = 12'h655;
rom[44768] = 12'h655;
rom[44769] = 12'h665;
rom[44770] = 12'h765;
rom[44771] = 12'h766;
rom[44772] = 12'h776;
rom[44773] = 12'h777;
rom[44774] = 12'h777;
rom[44775] = 12'h777;
rom[44776] = 12'h788;
rom[44777] = 12'h888;
rom[44778] = 12'h899;
rom[44779] = 12'h99a;
rom[44780] = 12'haaa;
rom[44781] = 12'haab;
rom[44782] = 12'hbbb;
rom[44783] = 12'hbbc;
rom[44784] = 12'hbbb;
rom[44785] = 12'hbbb;
rom[44786] = 12'hbbb;
rom[44787] = 12'hbbb;
rom[44788] = 12'haaa;
rom[44789] = 12'haaa;
rom[44790] = 12'haaa;
rom[44791] = 12'haaa;
rom[44792] = 12'h999;
rom[44793] = 12'h999;
rom[44794] = 12'h999;
rom[44795] = 12'h999;
rom[44796] = 12'haaa;
rom[44797] = 12'haaa;
rom[44798] = 12'haaa;
rom[44799] = 12'haaa;
rom[44800] = 12'h888;
rom[44801] = 12'h888;
rom[44802] = 12'h888;
rom[44803] = 12'h888;
rom[44804] = 12'h888;
rom[44805] = 12'h888;
rom[44806] = 12'h888;
rom[44807] = 12'h888;
rom[44808] = 12'h777;
rom[44809] = 12'h777;
rom[44810] = 12'h777;
rom[44811] = 12'h777;
rom[44812] = 12'h777;
rom[44813] = 12'h777;
rom[44814] = 12'h777;
rom[44815] = 12'h777;
rom[44816] = 12'h777;
rom[44817] = 12'h777;
rom[44818] = 12'h777;
rom[44819] = 12'h777;
rom[44820] = 12'h777;
rom[44821] = 12'h777;
rom[44822] = 12'h777;
rom[44823] = 12'h777;
rom[44824] = 12'h777;
rom[44825] = 12'h777;
rom[44826] = 12'h777;
rom[44827] = 12'h777;
rom[44828] = 12'h777;
rom[44829] = 12'h777;
rom[44830] = 12'h777;
rom[44831] = 12'h666;
rom[44832] = 12'h777;
rom[44833] = 12'h777;
rom[44834] = 12'h777;
rom[44835] = 12'h777;
rom[44836] = 12'h777;
rom[44837] = 12'h777;
rom[44838] = 12'h777;
rom[44839] = 12'h777;
rom[44840] = 12'h777;
rom[44841] = 12'h888;
rom[44842] = 12'h888;
rom[44843] = 12'h888;
rom[44844] = 12'h888;
rom[44845] = 12'h888;
rom[44846] = 12'h888;
rom[44847] = 12'h888;
rom[44848] = 12'h888;
rom[44849] = 12'h888;
rom[44850] = 12'h888;
rom[44851] = 12'h888;
rom[44852] = 12'h888;
rom[44853] = 12'h999;
rom[44854] = 12'h999;
rom[44855] = 12'h999;
rom[44856] = 12'h999;
rom[44857] = 12'h999;
rom[44858] = 12'h999;
rom[44859] = 12'haaa;
rom[44860] = 12'haaa;
rom[44861] = 12'haaa;
rom[44862] = 12'haaa;
rom[44863] = 12'haaa;
rom[44864] = 12'haaa;
rom[44865] = 12'haaa;
rom[44866] = 12'h999;
rom[44867] = 12'h888;
rom[44868] = 12'h888;
rom[44869] = 12'h888;
rom[44870] = 12'h777;
rom[44871] = 12'h777;
rom[44872] = 12'h777;
rom[44873] = 12'h777;
rom[44874] = 12'h777;
rom[44875] = 12'h777;
rom[44876] = 12'h777;
rom[44877] = 12'h666;
rom[44878] = 12'h666;
rom[44879] = 12'h666;
rom[44880] = 12'h666;
rom[44881] = 12'h555;
rom[44882] = 12'h555;
rom[44883] = 12'h555;
rom[44884] = 12'h555;
rom[44885] = 12'h555;
rom[44886] = 12'h555;
rom[44887] = 12'h555;
rom[44888] = 12'h555;
rom[44889] = 12'h555;
rom[44890] = 12'h666;
rom[44891] = 12'h666;
rom[44892] = 12'h666;
rom[44893] = 12'h777;
rom[44894] = 12'h666;
rom[44895] = 12'h666;
rom[44896] = 12'h666;
rom[44897] = 12'h666;
rom[44898] = 12'h555;
rom[44899] = 12'h555;
rom[44900] = 12'h444;
rom[44901] = 12'h444;
rom[44902] = 12'h444;
rom[44903] = 12'h333;
rom[44904] = 12'h222;
rom[44905] = 12'h222;
rom[44906] = 12'h333;
rom[44907] = 12'h333;
rom[44908] = 12'h333;
rom[44909] = 12'h222;
rom[44910] = 12'h111;
rom[44911] = 12'h111;
rom[44912] = 12'h111;
rom[44913] = 12'h111;
rom[44914] = 12'h111;
rom[44915] = 12'h111;
rom[44916] = 12'h111;
rom[44917] = 12'h111;
rom[44918] = 12'h111;
rom[44919] = 12'h  0;
rom[44920] = 12'h  0;
rom[44921] = 12'h  0;
rom[44922] = 12'h  0;
rom[44923] = 12'h  0;
rom[44924] = 12'h  0;
rom[44925] = 12'h  0;
rom[44926] = 12'h  0;
rom[44927] = 12'h  0;
rom[44928] = 12'h  0;
rom[44929] = 12'h  0;
rom[44930] = 12'h  0;
rom[44931] = 12'h  0;
rom[44932] = 12'h  0;
rom[44933] = 12'h  0;
rom[44934] = 12'h  0;
rom[44935] = 12'h  0;
rom[44936] = 12'h  0;
rom[44937] = 12'h  0;
rom[44938] = 12'h  0;
rom[44939] = 12'h  0;
rom[44940] = 12'h  0;
rom[44941] = 12'h  0;
rom[44942] = 12'h  0;
rom[44943] = 12'h  0;
rom[44944] = 12'h111;
rom[44945] = 12'h111;
rom[44946] = 12'h111;
rom[44947] = 12'h111;
rom[44948] = 12'h111;
rom[44949] = 12'h111;
rom[44950] = 12'h111;
rom[44951] = 12'h111;
rom[44952] = 12'h111;
rom[44953] = 12'h111;
rom[44954] = 12'h111;
rom[44955] = 12'h111;
rom[44956] = 12'h111;
rom[44957] = 12'h111;
rom[44958] = 12'h111;
rom[44959] = 12'h111;
rom[44960] = 12'h111;
rom[44961] = 12'h111;
rom[44962] = 12'h111;
rom[44963] = 12'h111;
rom[44964] = 12'h222;
rom[44965] = 12'h222;
rom[44966] = 12'h111;
rom[44967] = 12'h111;
rom[44968] = 12'h222;
rom[44969] = 12'h222;
rom[44970] = 12'h222;
rom[44971] = 12'h222;
rom[44972] = 12'h222;
rom[44973] = 12'h222;
rom[44974] = 12'h222;
rom[44975] = 12'h222;
rom[44976] = 12'h222;
rom[44977] = 12'h222;
rom[44978] = 12'h111;
rom[44979] = 12'h111;
rom[44980] = 12'h111;
rom[44981] = 12'h222;
rom[44982] = 12'h222;
rom[44983] = 12'h222;
rom[44984] = 12'h222;
rom[44985] = 12'h222;
rom[44986] = 12'h222;
rom[44987] = 12'h222;
rom[44988] = 12'h222;
rom[44989] = 12'h222;
rom[44990] = 12'h222;
rom[44991] = 12'h222;
rom[44992] = 12'h222;
rom[44993] = 12'h222;
rom[44994] = 12'h222;
rom[44995] = 12'h222;
rom[44996] = 12'h222;
rom[44997] = 12'h222;
rom[44998] = 12'h222;
rom[44999] = 12'h222;
rom[45000] = 12'h222;
rom[45001] = 12'h222;
rom[45002] = 12'h222;
rom[45003] = 12'h111;
rom[45004] = 12'h111;
rom[45005] = 12'h222;
rom[45006] = 12'h222;
rom[45007] = 12'h222;
rom[45008] = 12'h222;
rom[45009] = 12'h222;
rom[45010] = 12'h222;
rom[45011] = 12'h222;
rom[45012] = 12'h222;
rom[45013] = 12'h222;
rom[45014] = 12'h222;
rom[45015] = 12'h333;
rom[45016] = 12'h333;
rom[45017] = 12'h333;
rom[45018] = 12'h333;
rom[45019] = 12'h333;
rom[45020] = 12'h333;
rom[45021] = 12'h333;
rom[45022] = 12'h333;
rom[45023] = 12'h333;
rom[45024] = 12'h333;
rom[45025] = 12'h333;
rom[45026] = 12'h333;
rom[45027] = 12'h333;
rom[45028] = 12'h333;
rom[45029] = 12'h222;
rom[45030] = 12'h333;
rom[45031] = 12'h333;
rom[45032] = 12'h222;
rom[45033] = 12'h222;
rom[45034] = 12'h222;
rom[45035] = 12'h222;
rom[45036] = 12'h222;
rom[45037] = 12'h111;
rom[45038] = 12'h111;
rom[45039] = 12'h111;
rom[45040] = 12'h111;
rom[45041] = 12'h111;
rom[45042] = 12'h111;
rom[45043] = 12'h111;
rom[45044] = 12'h111;
rom[45045] = 12'h111;
rom[45046] = 12'h111;
rom[45047] = 12'h111;
rom[45048] = 12'h  0;
rom[45049] = 12'h  0;
rom[45050] = 12'h  0;
rom[45051] = 12'h  0;
rom[45052] = 12'h  0;
rom[45053] = 12'h  0;
rom[45054] = 12'h  0;
rom[45055] = 12'h  0;
rom[45056] = 12'h  0;
rom[45057] = 12'h  0;
rom[45058] = 12'h  0;
rom[45059] = 12'h  0;
rom[45060] = 12'h  0;
rom[45061] = 12'h  0;
rom[45062] = 12'h  0;
rom[45063] = 12'h  0;
rom[45064] = 12'h  0;
rom[45065] = 12'h  0;
rom[45066] = 12'h  0;
rom[45067] = 12'h  0;
rom[45068] = 12'h  0;
rom[45069] = 12'h  0;
rom[45070] = 12'h  0;
rom[45071] = 12'h  0;
rom[45072] = 12'h111;
rom[45073] = 12'h111;
rom[45074] = 12'h222;
rom[45075] = 12'h222;
rom[45076] = 12'h333;
rom[45077] = 12'h444;
rom[45078] = 12'h444;
rom[45079] = 12'h555;
rom[45080] = 12'h555;
rom[45081] = 12'h555;
rom[45082] = 12'h555;
rom[45083] = 12'h666;
rom[45084] = 12'h666;
rom[45085] = 12'h666;
rom[45086] = 12'h666;
rom[45087] = 12'h777;
rom[45088] = 12'h888;
rom[45089] = 12'h888;
rom[45090] = 12'h888;
rom[45091] = 12'h999;
rom[45092] = 12'haaa;
rom[45093] = 12'hbbb;
rom[45094] = 12'hccc;
rom[45095] = 12'hddd;
rom[45096] = 12'hbaa;
rom[45097] = 12'h665;
rom[45098] = 12'h211;
rom[45099] = 12'h100;
rom[45100] = 12'h211;
rom[45101] = 12'h200;
rom[45102] = 12'h200;
rom[45103] = 12'h200;
rom[45104] = 12'h200;
rom[45105] = 12'h200;
rom[45106] = 12'h200;
rom[45107] = 12'h200;
rom[45108] = 12'h200;
rom[45109] = 12'h200;
rom[45110] = 12'h200;
rom[45111] = 12'h200;
rom[45112] = 12'h200;
rom[45113] = 12'h300;
rom[45114] = 12'h300;
rom[45115] = 12'h300;
rom[45116] = 12'h300;
rom[45117] = 12'h300;
rom[45118] = 12'h300;
rom[45119] = 12'h300;
rom[45120] = 12'h300;
rom[45121] = 12'h300;
rom[45122] = 12'h300;
rom[45123] = 12'h300;
rom[45124] = 12'h400;
rom[45125] = 12'h400;
rom[45126] = 12'h400;
rom[45127] = 12'h400;
rom[45128] = 12'h400;
rom[45129] = 12'h400;
rom[45130] = 12'h400;
rom[45131] = 12'h400;
rom[45132] = 12'h400;
rom[45133] = 12'h400;
rom[45134] = 12'h400;
rom[45135] = 12'h400;
rom[45136] = 12'h300;
rom[45137] = 12'h300;
rom[45138] = 12'h300;
rom[45139] = 12'h400;
rom[45140] = 12'h400;
rom[45141] = 12'h400;
rom[45142] = 12'h510;
rom[45143] = 12'h510;
rom[45144] = 12'h510;
rom[45145] = 12'h510;
rom[45146] = 12'h510;
rom[45147] = 12'h510;
rom[45148] = 12'h510;
rom[45149] = 12'h520;
rom[45150] = 12'h520;
rom[45151] = 12'h520;
rom[45152] = 12'h520;
rom[45153] = 12'h520;
rom[45154] = 12'h520;
rom[45155] = 12'h520;
rom[45156] = 12'h420;
rom[45157] = 12'h421;
rom[45158] = 12'h532;
rom[45159] = 12'h532;
rom[45160] = 12'h533;
rom[45161] = 12'h543;
rom[45162] = 12'h543;
rom[45163] = 12'h544;
rom[45164] = 12'h544;
rom[45165] = 12'h554;
rom[45166] = 12'h554;
rom[45167] = 12'h654;
rom[45168] = 12'h655;
rom[45169] = 12'h665;
rom[45170] = 12'h766;
rom[45171] = 12'h776;
rom[45172] = 12'h777;
rom[45173] = 12'h777;
rom[45174] = 12'h877;
rom[45175] = 12'h878;
rom[45176] = 12'h888;
rom[45177] = 12'h989;
rom[45178] = 12'h999;
rom[45179] = 12'haaa;
rom[45180] = 12'hbab;
rom[45181] = 12'hbbb;
rom[45182] = 12'hbbb;
rom[45183] = 12'hbbb;
rom[45184] = 12'hbbb;
rom[45185] = 12'hbbb;
rom[45186] = 12'hbbb;
rom[45187] = 12'hbbb;
rom[45188] = 12'haaa;
rom[45189] = 12'haaa;
rom[45190] = 12'haaa;
rom[45191] = 12'haaa;
rom[45192] = 12'h999;
rom[45193] = 12'h999;
rom[45194] = 12'h999;
rom[45195] = 12'h999;
rom[45196] = 12'haaa;
rom[45197] = 12'haaa;
rom[45198] = 12'haaa;
rom[45199] = 12'haaa;
rom[45200] = 12'h888;
rom[45201] = 12'h888;
rom[45202] = 12'h888;
rom[45203] = 12'h888;
rom[45204] = 12'h888;
rom[45205] = 12'h888;
rom[45206] = 12'h888;
rom[45207] = 12'h888;
rom[45208] = 12'h888;
rom[45209] = 12'h888;
rom[45210] = 12'h888;
rom[45211] = 12'h888;
rom[45212] = 12'h888;
rom[45213] = 12'h888;
rom[45214] = 12'h777;
rom[45215] = 12'h777;
rom[45216] = 12'h777;
rom[45217] = 12'h777;
rom[45218] = 12'h777;
rom[45219] = 12'h777;
rom[45220] = 12'h777;
rom[45221] = 12'h666;
rom[45222] = 12'h666;
rom[45223] = 12'h666;
rom[45224] = 12'h777;
rom[45225] = 12'h777;
rom[45226] = 12'h777;
rom[45227] = 12'h777;
rom[45228] = 12'h777;
rom[45229] = 12'h777;
rom[45230] = 12'h777;
rom[45231] = 12'h666;
rom[45232] = 12'h777;
rom[45233] = 12'h777;
rom[45234] = 12'h777;
rom[45235] = 12'h777;
rom[45236] = 12'h777;
rom[45237] = 12'h777;
rom[45238] = 12'h777;
rom[45239] = 12'h777;
rom[45240] = 12'h777;
rom[45241] = 12'h777;
rom[45242] = 12'h777;
rom[45243] = 12'h777;
rom[45244] = 12'h777;
rom[45245] = 12'h777;
rom[45246] = 12'h777;
rom[45247] = 12'h777;
rom[45248] = 12'h888;
rom[45249] = 12'h888;
rom[45250] = 12'h888;
rom[45251] = 12'h888;
rom[45252] = 12'h888;
rom[45253] = 12'h888;
rom[45254] = 12'h999;
rom[45255] = 12'h999;
rom[45256] = 12'h999;
rom[45257] = 12'h999;
rom[45258] = 12'h999;
rom[45259] = 12'h999;
rom[45260] = 12'haaa;
rom[45261] = 12'haaa;
rom[45262] = 12'haaa;
rom[45263] = 12'haaa;
rom[45264] = 12'haaa;
rom[45265] = 12'haaa;
rom[45266] = 12'h999;
rom[45267] = 12'h999;
rom[45268] = 12'h888;
rom[45269] = 12'h888;
rom[45270] = 12'h777;
rom[45271] = 12'h777;
rom[45272] = 12'h777;
rom[45273] = 12'h777;
rom[45274] = 12'h777;
rom[45275] = 12'h777;
rom[45276] = 12'h777;
rom[45277] = 12'h666;
rom[45278] = 12'h666;
rom[45279] = 12'h666;
rom[45280] = 12'h666;
rom[45281] = 12'h666;
rom[45282] = 12'h555;
rom[45283] = 12'h555;
rom[45284] = 12'h555;
rom[45285] = 12'h555;
rom[45286] = 12'h555;
rom[45287] = 12'h555;
rom[45288] = 12'h555;
rom[45289] = 12'h555;
rom[45290] = 12'h666;
rom[45291] = 12'h666;
rom[45292] = 12'h666;
rom[45293] = 12'h666;
rom[45294] = 12'h666;
rom[45295] = 12'h666;
rom[45296] = 12'h666;
rom[45297] = 12'h555;
rom[45298] = 12'h555;
rom[45299] = 12'h555;
rom[45300] = 12'h555;
rom[45301] = 12'h444;
rom[45302] = 12'h444;
rom[45303] = 12'h333;
rom[45304] = 12'h333;
rom[45305] = 12'h333;
rom[45306] = 12'h333;
rom[45307] = 12'h333;
rom[45308] = 12'h333;
rom[45309] = 12'h222;
rom[45310] = 12'h222;
rom[45311] = 12'h111;
rom[45312] = 12'h111;
rom[45313] = 12'h111;
rom[45314] = 12'h  0;
rom[45315] = 12'h  0;
rom[45316] = 12'h  0;
rom[45317] = 12'h  0;
rom[45318] = 12'h  0;
rom[45319] = 12'h  0;
rom[45320] = 12'h  0;
rom[45321] = 12'h  0;
rom[45322] = 12'h  0;
rom[45323] = 12'h  0;
rom[45324] = 12'h  0;
rom[45325] = 12'h  0;
rom[45326] = 12'h  0;
rom[45327] = 12'h  0;
rom[45328] = 12'h  0;
rom[45329] = 12'h  0;
rom[45330] = 12'h  0;
rom[45331] = 12'h  0;
rom[45332] = 12'h  0;
rom[45333] = 12'h  0;
rom[45334] = 12'h  0;
rom[45335] = 12'h  0;
rom[45336] = 12'h  0;
rom[45337] = 12'h  0;
rom[45338] = 12'h  0;
rom[45339] = 12'h  0;
rom[45340] = 12'h  0;
rom[45341] = 12'h  0;
rom[45342] = 12'h  0;
rom[45343] = 12'h  0;
rom[45344] = 12'h111;
rom[45345] = 12'h111;
rom[45346] = 12'h111;
rom[45347] = 12'h111;
rom[45348] = 12'h111;
rom[45349] = 12'h111;
rom[45350] = 12'h111;
rom[45351] = 12'h111;
rom[45352] = 12'h111;
rom[45353] = 12'h111;
rom[45354] = 12'h111;
rom[45355] = 12'h111;
rom[45356] = 12'h111;
rom[45357] = 12'h111;
rom[45358] = 12'h111;
rom[45359] = 12'h111;
rom[45360] = 12'h111;
rom[45361] = 12'h111;
rom[45362] = 12'h111;
rom[45363] = 12'h111;
rom[45364] = 12'h222;
rom[45365] = 12'h111;
rom[45366] = 12'h111;
rom[45367] = 12'h111;
rom[45368] = 12'h222;
rom[45369] = 12'h222;
rom[45370] = 12'h222;
rom[45371] = 12'h222;
rom[45372] = 12'h111;
rom[45373] = 12'h111;
rom[45374] = 12'h111;
rom[45375] = 12'h111;
rom[45376] = 12'h222;
rom[45377] = 12'h111;
rom[45378] = 12'h111;
rom[45379] = 12'h111;
rom[45380] = 12'h111;
rom[45381] = 12'h222;
rom[45382] = 12'h222;
rom[45383] = 12'h222;
rom[45384] = 12'h222;
rom[45385] = 12'h222;
rom[45386] = 12'h222;
rom[45387] = 12'h222;
rom[45388] = 12'h222;
rom[45389] = 12'h222;
rom[45390] = 12'h222;
rom[45391] = 12'h222;
rom[45392] = 12'h222;
rom[45393] = 12'h222;
rom[45394] = 12'h222;
rom[45395] = 12'h222;
rom[45396] = 12'h222;
rom[45397] = 12'h111;
rom[45398] = 12'h111;
rom[45399] = 12'h111;
rom[45400] = 12'h111;
rom[45401] = 12'h111;
rom[45402] = 12'h111;
rom[45403] = 12'h111;
rom[45404] = 12'h111;
rom[45405] = 12'h111;
rom[45406] = 12'h111;
rom[45407] = 12'h111;
rom[45408] = 12'h111;
rom[45409] = 12'h222;
rom[45410] = 12'h222;
rom[45411] = 12'h222;
rom[45412] = 12'h222;
rom[45413] = 12'h222;
rom[45414] = 12'h222;
rom[45415] = 12'h222;
rom[45416] = 12'h333;
rom[45417] = 12'h333;
rom[45418] = 12'h333;
rom[45419] = 12'h333;
rom[45420] = 12'h333;
rom[45421] = 12'h333;
rom[45422] = 12'h333;
rom[45423] = 12'h333;
rom[45424] = 12'h333;
rom[45425] = 12'h333;
rom[45426] = 12'h333;
rom[45427] = 12'h333;
rom[45428] = 12'h222;
rom[45429] = 12'h222;
rom[45430] = 12'h222;
rom[45431] = 12'h222;
rom[45432] = 12'h222;
rom[45433] = 12'h222;
rom[45434] = 12'h222;
rom[45435] = 12'h111;
rom[45436] = 12'h111;
rom[45437] = 12'h111;
rom[45438] = 12'h111;
rom[45439] = 12'h111;
rom[45440] = 12'h111;
rom[45441] = 12'h111;
rom[45442] = 12'h111;
rom[45443] = 12'h111;
rom[45444] = 12'h111;
rom[45445] = 12'h  0;
rom[45446] = 12'h  0;
rom[45447] = 12'h  0;
rom[45448] = 12'h  0;
rom[45449] = 12'h  0;
rom[45450] = 12'h  0;
rom[45451] = 12'h  0;
rom[45452] = 12'h  0;
rom[45453] = 12'h  0;
rom[45454] = 12'h  0;
rom[45455] = 12'h  0;
rom[45456] = 12'h  0;
rom[45457] = 12'h  0;
rom[45458] = 12'h  0;
rom[45459] = 12'h  0;
rom[45460] = 12'h  0;
rom[45461] = 12'h  0;
rom[45462] = 12'h  0;
rom[45463] = 12'h  0;
rom[45464] = 12'h  0;
rom[45465] = 12'h  0;
rom[45466] = 12'h  0;
rom[45467] = 12'h  0;
rom[45468] = 12'h  0;
rom[45469] = 12'h  0;
rom[45470] = 12'h111;
rom[45471] = 12'h111;
rom[45472] = 12'h111;
rom[45473] = 12'h111;
rom[45474] = 12'h222;
rom[45475] = 12'h222;
rom[45476] = 12'h333;
rom[45477] = 12'h444;
rom[45478] = 12'h444;
rom[45479] = 12'h555;
rom[45480] = 12'h555;
rom[45481] = 12'h555;
rom[45482] = 12'h555;
rom[45483] = 12'h666;
rom[45484] = 12'h666;
rom[45485] = 12'h666;
rom[45486] = 12'h666;
rom[45487] = 12'h777;
rom[45488] = 12'h787;
rom[45489] = 12'h888;
rom[45490] = 12'h888;
rom[45491] = 12'h999;
rom[45492] = 12'haaa;
rom[45493] = 12'hbbb;
rom[45494] = 12'hccc;
rom[45495] = 12'hccc;
rom[45496] = 12'haaa;
rom[45497] = 12'h665;
rom[45498] = 12'h222;
rom[45499] = 12'h100;
rom[45500] = 12'h211;
rom[45501] = 12'h100;
rom[45502] = 12'h100;
rom[45503] = 12'h100;
rom[45504] = 12'h100;
rom[45505] = 12'h100;
rom[45506] = 12'h100;
rom[45507] = 12'h100;
rom[45508] = 12'h100;
rom[45509] = 12'h200;
rom[45510] = 12'h200;
rom[45511] = 12'h200;
rom[45512] = 12'h200;
rom[45513] = 12'h200;
rom[45514] = 12'h200;
rom[45515] = 12'h200;
rom[45516] = 12'h200;
rom[45517] = 12'h200;
rom[45518] = 12'h200;
rom[45519] = 12'h200;
rom[45520] = 12'h300;
rom[45521] = 12'h300;
rom[45522] = 12'h300;
rom[45523] = 12'h300;
rom[45524] = 12'h300;
rom[45525] = 12'h300;
rom[45526] = 12'h300;
rom[45527] = 12'h300;
rom[45528] = 12'h300;
rom[45529] = 12'h300;
rom[45530] = 12'h300;
rom[45531] = 12'h300;
rom[45532] = 12'h300;
rom[45533] = 12'h300;
rom[45534] = 12'h300;
rom[45535] = 12'h300;
rom[45536] = 12'h300;
rom[45537] = 12'h300;
rom[45538] = 12'h300;
rom[45539] = 12'h300;
rom[45540] = 12'h400;
rom[45541] = 12'h400;
rom[45542] = 12'h500;
rom[45543] = 12'h510;
rom[45544] = 12'h510;
rom[45545] = 12'h510;
rom[45546] = 12'h510;
rom[45547] = 12'h510;
rom[45548] = 12'h510;
rom[45549] = 12'h510;
rom[45550] = 12'h510;
rom[45551] = 12'h520;
rom[45552] = 12'h520;
rom[45553] = 12'h520;
rom[45554] = 12'h520;
rom[45555] = 12'h521;
rom[45556] = 12'h421;
rom[45557] = 12'h422;
rom[45558] = 12'h532;
rom[45559] = 12'h533;
rom[45560] = 12'h533;
rom[45561] = 12'h544;
rom[45562] = 12'h544;
rom[45563] = 12'h544;
rom[45564] = 12'h554;
rom[45565] = 12'h554;
rom[45566] = 12'h654;
rom[45567] = 12'h655;
rom[45568] = 12'h665;
rom[45569] = 12'h666;
rom[45570] = 12'h776;
rom[45571] = 12'h777;
rom[45572] = 12'h777;
rom[45573] = 12'h877;
rom[45574] = 12'h888;
rom[45575] = 12'h888;
rom[45576] = 12'h988;
rom[45577] = 12'h999;
rom[45578] = 12'ha9a;
rom[45579] = 12'hbaa;
rom[45580] = 12'hbbb;
rom[45581] = 12'hbbb;
rom[45582] = 12'hcbc;
rom[45583] = 12'hcbb;
rom[45584] = 12'hbbb;
rom[45585] = 12'hbbb;
rom[45586] = 12'hbbb;
rom[45587] = 12'hbbb;
rom[45588] = 12'haaa;
rom[45589] = 12'haaa;
rom[45590] = 12'haaa;
rom[45591] = 12'haaa;
rom[45592] = 12'h999;
rom[45593] = 12'h999;
rom[45594] = 12'h999;
rom[45595] = 12'h999;
rom[45596] = 12'haaa;
rom[45597] = 12'haaa;
rom[45598] = 12'haaa;
rom[45599] = 12'haaa;
rom[45600] = 12'h999;
rom[45601] = 12'h999;
rom[45602] = 12'h999;
rom[45603] = 12'h999;
rom[45604] = 12'h999;
rom[45605] = 12'h999;
rom[45606] = 12'h999;
rom[45607] = 12'h999;
rom[45608] = 12'h999;
rom[45609] = 12'h999;
rom[45610] = 12'h888;
rom[45611] = 12'h888;
rom[45612] = 12'h888;
rom[45613] = 12'h888;
rom[45614] = 12'h777;
rom[45615] = 12'h777;
rom[45616] = 12'h777;
rom[45617] = 12'h777;
rom[45618] = 12'h777;
rom[45619] = 12'h666;
rom[45620] = 12'h666;
rom[45621] = 12'h666;
rom[45622] = 12'h666;
rom[45623] = 12'h666;
rom[45624] = 12'h666;
rom[45625] = 12'h777;
rom[45626] = 12'h777;
rom[45627] = 12'h777;
rom[45628] = 12'h777;
rom[45629] = 12'h777;
rom[45630] = 12'h777;
rom[45631] = 12'h777;
rom[45632] = 12'h777;
rom[45633] = 12'h777;
rom[45634] = 12'h777;
rom[45635] = 12'h888;
rom[45636] = 12'h888;
rom[45637] = 12'h777;
rom[45638] = 12'h777;
rom[45639] = 12'h777;
rom[45640] = 12'h777;
rom[45641] = 12'h777;
rom[45642] = 12'h777;
rom[45643] = 12'h777;
rom[45644] = 12'h777;
rom[45645] = 12'h777;
rom[45646] = 12'h777;
rom[45647] = 12'h777;
rom[45648] = 12'h777;
rom[45649] = 12'h888;
rom[45650] = 12'h888;
rom[45651] = 12'h888;
rom[45652] = 12'h888;
rom[45653] = 12'h888;
rom[45654] = 12'h999;
rom[45655] = 12'h999;
rom[45656] = 12'h999;
rom[45657] = 12'h999;
rom[45658] = 12'h999;
rom[45659] = 12'h999;
rom[45660] = 12'h999;
rom[45661] = 12'haaa;
rom[45662] = 12'haaa;
rom[45663] = 12'haaa;
rom[45664] = 12'haaa;
rom[45665] = 12'haaa;
rom[45666] = 12'haaa;
rom[45667] = 12'h999;
rom[45668] = 12'h999;
rom[45669] = 12'h888;
rom[45670] = 12'h777;
rom[45671] = 12'h777;
rom[45672] = 12'h777;
rom[45673] = 12'h777;
rom[45674] = 12'h666;
rom[45675] = 12'h777;
rom[45676] = 12'h777;
rom[45677] = 12'h666;
rom[45678] = 12'h666;
rom[45679] = 12'h666;
rom[45680] = 12'h666;
rom[45681] = 12'h666;
rom[45682] = 12'h555;
rom[45683] = 12'h555;
rom[45684] = 12'h555;
rom[45685] = 12'h555;
rom[45686] = 12'h555;
rom[45687] = 12'h555;
rom[45688] = 12'h555;
rom[45689] = 12'h555;
rom[45690] = 12'h555;
rom[45691] = 12'h666;
rom[45692] = 12'h666;
rom[45693] = 12'h666;
rom[45694] = 12'h666;
rom[45695] = 12'h666;
rom[45696] = 12'h666;
rom[45697] = 12'h555;
rom[45698] = 12'h555;
rom[45699] = 12'h555;
rom[45700] = 12'h555;
rom[45701] = 12'h555;
rom[45702] = 12'h444;
rom[45703] = 12'h444;
rom[45704] = 12'h333;
rom[45705] = 12'h333;
rom[45706] = 12'h333;
rom[45707] = 12'h333;
rom[45708] = 12'h333;
rom[45709] = 12'h333;
rom[45710] = 12'h222;
rom[45711] = 12'h222;
rom[45712] = 12'h111;
rom[45713] = 12'h111;
rom[45714] = 12'h  0;
rom[45715] = 12'h  0;
rom[45716] = 12'h  0;
rom[45717] = 12'h  0;
rom[45718] = 12'h  0;
rom[45719] = 12'h  0;
rom[45720] = 12'h  0;
rom[45721] = 12'h  0;
rom[45722] = 12'h  0;
rom[45723] = 12'h  0;
rom[45724] = 12'h  0;
rom[45725] = 12'h  0;
rom[45726] = 12'h  0;
rom[45727] = 12'h  0;
rom[45728] = 12'h  0;
rom[45729] = 12'h  0;
rom[45730] = 12'h  0;
rom[45731] = 12'h  0;
rom[45732] = 12'h  0;
rom[45733] = 12'h  0;
rom[45734] = 12'h  0;
rom[45735] = 12'h  0;
rom[45736] = 12'h  0;
rom[45737] = 12'h  0;
rom[45738] = 12'h  0;
rom[45739] = 12'h  0;
rom[45740] = 12'h  0;
rom[45741] = 12'h  0;
rom[45742] = 12'h  0;
rom[45743] = 12'h  0;
rom[45744] = 12'h  0;
rom[45745] = 12'h  0;
rom[45746] = 12'h111;
rom[45747] = 12'h111;
rom[45748] = 12'h111;
rom[45749] = 12'h111;
rom[45750] = 12'h111;
rom[45751] = 12'h111;
rom[45752] = 12'h111;
rom[45753] = 12'h111;
rom[45754] = 12'h111;
rom[45755] = 12'h111;
rom[45756] = 12'h111;
rom[45757] = 12'h111;
rom[45758] = 12'h111;
rom[45759] = 12'h111;
rom[45760] = 12'h111;
rom[45761] = 12'h111;
rom[45762] = 12'h111;
rom[45763] = 12'h111;
rom[45764] = 12'h111;
rom[45765] = 12'h111;
rom[45766] = 12'h111;
rom[45767] = 12'h111;
rom[45768] = 12'h222;
rom[45769] = 12'h222;
rom[45770] = 12'h222;
rom[45771] = 12'h222;
rom[45772] = 12'h111;
rom[45773] = 12'h111;
rom[45774] = 12'h111;
rom[45775] = 12'h111;
rom[45776] = 12'h111;
rom[45777] = 12'h111;
rom[45778] = 12'h111;
rom[45779] = 12'h111;
rom[45780] = 12'h222;
rom[45781] = 12'h222;
rom[45782] = 12'h222;
rom[45783] = 12'h222;
rom[45784] = 12'h222;
rom[45785] = 12'h222;
rom[45786] = 12'h222;
rom[45787] = 12'h222;
rom[45788] = 12'h222;
rom[45789] = 12'h222;
rom[45790] = 12'h222;
rom[45791] = 12'h222;
rom[45792] = 12'h222;
rom[45793] = 12'h222;
rom[45794] = 12'h222;
rom[45795] = 12'h111;
rom[45796] = 12'h111;
rom[45797] = 12'h111;
rom[45798] = 12'h111;
rom[45799] = 12'h111;
rom[45800] = 12'h111;
rom[45801] = 12'h111;
rom[45802] = 12'h111;
rom[45803] = 12'h111;
rom[45804] = 12'h111;
rom[45805] = 12'h111;
rom[45806] = 12'h111;
rom[45807] = 12'h111;
rom[45808] = 12'h111;
rom[45809] = 12'h111;
rom[45810] = 12'h222;
rom[45811] = 12'h222;
rom[45812] = 12'h222;
rom[45813] = 12'h222;
rom[45814] = 12'h222;
rom[45815] = 12'h222;
rom[45816] = 12'h222;
rom[45817] = 12'h222;
rom[45818] = 12'h333;
rom[45819] = 12'h333;
rom[45820] = 12'h333;
rom[45821] = 12'h333;
rom[45822] = 12'h333;
rom[45823] = 12'h333;
rom[45824] = 12'h333;
rom[45825] = 12'h333;
rom[45826] = 12'h222;
rom[45827] = 12'h222;
rom[45828] = 12'h222;
rom[45829] = 12'h222;
rom[45830] = 12'h222;
rom[45831] = 12'h222;
rom[45832] = 12'h222;
rom[45833] = 12'h222;
rom[45834] = 12'h111;
rom[45835] = 12'h111;
rom[45836] = 12'h111;
rom[45837] = 12'h111;
rom[45838] = 12'h111;
rom[45839] = 12'h111;
rom[45840] = 12'h111;
rom[45841] = 12'h111;
rom[45842] = 12'h111;
rom[45843] = 12'h  0;
rom[45844] = 12'h  0;
rom[45845] = 12'h  0;
rom[45846] = 12'h  0;
rom[45847] = 12'h  0;
rom[45848] = 12'h  0;
rom[45849] = 12'h  0;
rom[45850] = 12'h  0;
rom[45851] = 12'h  0;
rom[45852] = 12'h  0;
rom[45853] = 12'h  0;
rom[45854] = 12'h  0;
rom[45855] = 12'h  0;
rom[45856] = 12'h  0;
rom[45857] = 12'h  0;
rom[45858] = 12'h  0;
rom[45859] = 12'h  0;
rom[45860] = 12'h  0;
rom[45861] = 12'h  0;
rom[45862] = 12'h  0;
rom[45863] = 12'h  0;
rom[45864] = 12'h  0;
rom[45865] = 12'h  0;
rom[45866] = 12'h  0;
rom[45867] = 12'h  0;
rom[45868] = 12'h111;
rom[45869] = 12'h111;
rom[45870] = 12'h111;
rom[45871] = 12'h111;
rom[45872] = 12'h111;
rom[45873] = 12'h222;
rom[45874] = 12'h222;
rom[45875] = 12'h222;
rom[45876] = 12'h333;
rom[45877] = 12'h444;
rom[45878] = 12'h555;
rom[45879] = 12'h555;
rom[45880] = 12'h555;
rom[45881] = 12'h555;
rom[45882] = 12'h555;
rom[45883] = 12'h555;
rom[45884] = 12'h666;
rom[45885] = 12'h666;
rom[45886] = 12'h666;
rom[45887] = 12'h777;
rom[45888] = 12'h777;
rom[45889] = 12'h888;
rom[45890] = 12'h898;
rom[45891] = 12'h999;
rom[45892] = 12'haaa;
rom[45893] = 12'hbbb;
rom[45894] = 12'hbbb;
rom[45895] = 12'hbbb;
rom[45896] = 12'h999;
rom[45897] = 12'h655;
rom[45898] = 12'h222;
rom[45899] = 12'h111;
rom[45900] = 12'h100;
rom[45901] = 12'h100;
rom[45902] = 12'h100;
rom[45903] = 12'h100;
rom[45904] = 12'h100;
rom[45905] = 12'h100;
rom[45906] = 12'h100;
rom[45907] = 12'h100;
rom[45908] = 12'h100;
rom[45909] = 12'h100;
rom[45910] = 12'h100;
rom[45911] = 12'h100;
rom[45912] = 12'h100;
rom[45913] = 12'h200;
rom[45914] = 12'h200;
rom[45915] = 12'h200;
rom[45916] = 12'h200;
rom[45917] = 12'h200;
rom[45918] = 12'h200;
rom[45919] = 12'h200;
rom[45920] = 12'h200;
rom[45921] = 12'h200;
rom[45922] = 12'h200;
rom[45923] = 12'h200;
rom[45924] = 12'h200;
rom[45925] = 12'h200;
rom[45926] = 12'h200;
rom[45927] = 12'h200;
rom[45928] = 12'h200;
rom[45929] = 12'h200;
rom[45930] = 12'h300;
rom[45931] = 12'h300;
rom[45932] = 12'h300;
rom[45933] = 12'h300;
rom[45934] = 12'h300;
rom[45935] = 12'h300;
rom[45936] = 12'h300;
rom[45937] = 12'h300;
rom[45938] = 12'h300;
rom[45939] = 12'h300;
rom[45940] = 12'h400;
rom[45941] = 12'h400;
rom[45942] = 12'h500;
rom[45943] = 12'h500;
rom[45944] = 12'h510;
rom[45945] = 12'h510;
rom[45946] = 12'h510;
rom[45947] = 12'h510;
rom[45948] = 12'h510;
rom[45949] = 12'h510;
rom[45950] = 12'h510;
rom[45951] = 12'h520;
rom[45952] = 12'h520;
rom[45953] = 12'h520;
rom[45954] = 12'h520;
rom[45955] = 12'h521;
rom[45956] = 12'h421;
rom[45957] = 12'h432;
rom[45958] = 12'h533;
rom[45959] = 12'h533;
rom[45960] = 12'h544;
rom[45961] = 12'h544;
rom[45962] = 12'h544;
rom[45963] = 12'h555;
rom[45964] = 12'h655;
rom[45965] = 12'h655;
rom[45966] = 12'h665;
rom[45967] = 12'h665;
rom[45968] = 12'h766;
rom[45969] = 12'h776;
rom[45970] = 12'h777;
rom[45971] = 12'h877;
rom[45972] = 12'h887;
rom[45973] = 12'h888;
rom[45974] = 12'h888;
rom[45975] = 12'h888;
rom[45976] = 12'h999;
rom[45977] = 12'ha99;
rom[45978] = 12'haaa;
rom[45979] = 12'hbbb;
rom[45980] = 12'hcbc;
rom[45981] = 12'hcbc;
rom[45982] = 12'hcbc;
rom[45983] = 12'hcbc;
rom[45984] = 12'hbbb;
rom[45985] = 12'hbbb;
rom[45986] = 12'hbbb;
rom[45987] = 12'hbbb;
rom[45988] = 12'haaa;
rom[45989] = 12'haaa;
rom[45990] = 12'haaa;
rom[45991] = 12'haaa;
rom[45992] = 12'h999;
rom[45993] = 12'h999;
rom[45994] = 12'h999;
rom[45995] = 12'haaa;
rom[45996] = 12'haaa;
rom[45997] = 12'haaa;
rom[45998] = 12'haaa;
rom[45999] = 12'haaa;
rom[46000] = 12'haaa;
rom[46001] = 12'haaa;
rom[46002] = 12'haaa;
rom[46003] = 12'h999;
rom[46004] = 12'h999;
rom[46005] = 12'h999;
rom[46006] = 12'h999;
rom[46007] = 12'h999;
rom[46008] = 12'h888;
rom[46009] = 12'h888;
rom[46010] = 12'h888;
rom[46011] = 12'h777;
rom[46012] = 12'h777;
rom[46013] = 12'h777;
rom[46014] = 12'h777;
rom[46015] = 12'h666;
rom[46016] = 12'h777;
rom[46017] = 12'h666;
rom[46018] = 12'h666;
rom[46019] = 12'h666;
rom[46020] = 12'h666;
rom[46021] = 12'h666;
rom[46022] = 12'h666;
rom[46023] = 12'h666;
rom[46024] = 12'h666;
rom[46025] = 12'h777;
rom[46026] = 12'h777;
rom[46027] = 12'h777;
rom[46028] = 12'h777;
rom[46029] = 12'h777;
rom[46030] = 12'h777;
rom[46031] = 12'h777;
rom[46032] = 12'h777;
rom[46033] = 12'h777;
rom[46034] = 12'h777;
rom[46035] = 12'h888;
rom[46036] = 12'h888;
rom[46037] = 12'h777;
rom[46038] = 12'h777;
rom[46039] = 12'h777;
rom[46040] = 12'h777;
rom[46041] = 12'h777;
rom[46042] = 12'h777;
rom[46043] = 12'h777;
rom[46044] = 12'h777;
rom[46045] = 12'h888;
rom[46046] = 12'h888;
rom[46047] = 12'h888;
rom[46048] = 12'h777;
rom[46049] = 12'h888;
rom[46050] = 12'h888;
rom[46051] = 12'h888;
rom[46052] = 12'h888;
rom[46053] = 12'h888;
rom[46054] = 12'h888;
rom[46055] = 12'h999;
rom[46056] = 12'h999;
rom[46057] = 12'h999;
rom[46058] = 12'h999;
rom[46059] = 12'h999;
rom[46060] = 12'h999;
rom[46061] = 12'haaa;
rom[46062] = 12'haaa;
rom[46063] = 12'haaa;
rom[46064] = 12'haaa;
rom[46065] = 12'haaa;
rom[46066] = 12'haaa;
rom[46067] = 12'haaa;
rom[46068] = 12'h999;
rom[46069] = 12'h888;
rom[46070] = 12'h888;
rom[46071] = 12'h777;
rom[46072] = 12'h777;
rom[46073] = 12'h777;
rom[46074] = 12'h777;
rom[46075] = 12'h777;
rom[46076] = 12'h777;
rom[46077] = 12'h666;
rom[46078] = 12'h666;
rom[46079] = 12'h666;
rom[46080] = 12'h666;
rom[46081] = 12'h666;
rom[46082] = 12'h666;
rom[46083] = 12'h555;
rom[46084] = 12'h555;
rom[46085] = 12'h555;
rom[46086] = 12'h555;
rom[46087] = 12'h555;
rom[46088] = 12'h555;
rom[46089] = 12'h555;
rom[46090] = 12'h555;
rom[46091] = 12'h555;
rom[46092] = 12'h666;
rom[46093] = 12'h666;
rom[46094] = 12'h666;
rom[46095] = 12'h666;
rom[46096] = 12'h666;
rom[46097] = 12'h666;
rom[46098] = 12'h555;
rom[46099] = 12'h555;
rom[46100] = 12'h555;
rom[46101] = 12'h555;
rom[46102] = 12'h444;
rom[46103] = 12'h444;
rom[46104] = 12'h444;
rom[46105] = 12'h333;
rom[46106] = 12'h333;
rom[46107] = 12'h333;
rom[46108] = 12'h333;
rom[46109] = 12'h333;
rom[46110] = 12'h333;
rom[46111] = 12'h222;
rom[46112] = 12'h111;
rom[46113] = 12'h111;
rom[46114] = 12'h111;
rom[46115] = 12'h  0;
rom[46116] = 12'h  0;
rom[46117] = 12'h  0;
rom[46118] = 12'h  0;
rom[46119] = 12'h  0;
rom[46120] = 12'h  0;
rom[46121] = 12'h  0;
rom[46122] = 12'h  0;
rom[46123] = 12'h  0;
rom[46124] = 12'h  0;
rom[46125] = 12'h  0;
rom[46126] = 12'h  0;
rom[46127] = 12'h  0;
rom[46128] = 12'h  0;
rom[46129] = 12'h  0;
rom[46130] = 12'h  0;
rom[46131] = 12'h  0;
rom[46132] = 12'h  0;
rom[46133] = 12'h  0;
rom[46134] = 12'h  0;
rom[46135] = 12'h  0;
rom[46136] = 12'h  0;
rom[46137] = 12'h  0;
rom[46138] = 12'h  0;
rom[46139] = 12'h  0;
rom[46140] = 12'h  0;
rom[46141] = 12'h  0;
rom[46142] = 12'h  0;
rom[46143] = 12'h  0;
rom[46144] = 12'h  0;
rom[46145] = 12'h  0;
rom[46146] = 12'h  0;
rom[46147] = 12'h111;
rom[46148] = 12'h111;
rom[46149] = 12'h111;
rom[46150] = 12'h111;
rom[46151] = 12'h111;
rom[46152] = 12'h111;
rom[46153] = 12'h111;
rom[46154] = 12'h111;
rom[46155] = 12'h111;
rom[46156] = 12'h111;
rom[46157] = 12'h111;
rom[46158] = 12'h111;
rom[46159] = 12'h111;
rom[46160] = 12'h111;
rom[46161] = 12'h111;
rom[46162] = 12'h111;
rom[46163] = 12'h111;
rom[46164] = 12'h111;
rom[46165] = 12'h111;
rom[46166] = 12'h111;
rom[46167] = 12'h111;
rom[46168] = 12'h222;
rom[46169] = 12'h222;
rom[46170] = 12'h222;
rom[46171] = 12'h111;
rom[46172] = 12'h111;
rom[46173] = 12'h111;
rom[46174] = 12'h111;
rom[46175] = 12'h111;
rom[46176] = 12'h111;
rom[46177] = 12'h111;
rom[46178] = 12'h111;
rom[46179] = 12'h222;
rom[46180] = 12'h222;
rom[46181] = 12'h222;
rom[46182] = 12'h222;
rom[46183] = 12'h222;
rom[46184] = 12'h222;
rom[46185] = 12'h222;
rom[46186] = 12'h222;
rom[46187] = 12'h222;
rom[46188] = 12'h222;
rom[46189] = 12'h222;
rom[46190] = 12'h222;
rom[46191] = 12'h222;
rom[46192] = 12'h111;
rom[46193] = 12'h111;
rom[46194] = 12'h111;
rom[46195] = 12'h111;
rom[46196] = 12'h111;
rom[46197] = 12'h111;
rom[46198] = 12'h111;
rom[46199] = 12'h111;
rom[46200] = 12'h111;
rom[46201] = 12'h111;
rom[46202] = 12'h111;
rom[46203] = 12'h111;
rom[46204] = 12'h111;
rom[46205] = 12'h111;
rom[46206] = 12'h111;
rom[46207] = 12'h111;
rom[46208] = 12'h111;
rom[46209] = 12'h111;
rom[46210] = 12'h222;
rom[46211] = 12'h222;
rom[46212] = 12'h222;
rom[46213] = 12'h222;
rom[46214] = 12'h222;
rom[46215] = 12'h222;
rom[46216] = 12'h222;
rom[46217] = 12'h222;
rom[46218] = 12'h222;
rom[46219] = 12'h333;
rom[46220] = 12'h333;
rom[46221] = 12'h333;
rom[46222] = 12'h333;
rom[46223] = 12'h333;
rom[46224] = 12'h333;
rom[46225] = 12'h222;
rom[46226] = 12'h222;
rom[46227] = 12'h222;
rom[46228] = 12'h222;
rom[46229] = 12'h222;
rom[46230] = 12'h222;
rom[46231] = 12'h222;
rom[46232] = 12'h222;
rom[46233] = 12'h222;
rom[46234] = 12'h111;
rom[46235] = 12'h111;
rom[46236] = 12'h111;
rom[46237] = 12'h111;
rom[46238] = 12'h111;
rom[46239] = 12'h111;
rom[46240] = 12'h111;
rom[46241] = 12'h111;
rom[46242] = 12'h  0;
rom[46243] = 12'h  0;
rom[46244] = 12'h  0;
rom[46245] = 12'h  0;
rom[46246] = 12'h  0;
rom[46247] = 12'h  0;
rom[46248] = 12'h  0;
rom[46249] = 12'h  0;
rom[46250] = 12'h  0;
rom[46251] = 12'h  0;
rom[46252] = 12'h  0;
rom[46253] = 12'h  0;
rom[46254] = 12'h  0;
rom[46255] = 12'h  0;
rom[46256] = 12'h  0;
rom[46257] = 12'h  0;
rom[46258] = 12'h  0;
rom[46259] = 12'h  0;
rom[46260] = 12'h  0;
rom[46261] = 12'h  0;
rom[46262] = 12'h  0;
rom[46263] = 12'h  0;
rom[46264] = 12'h  0;
rom[46265] = 12'h  0;
rom[46266] = 12'h  0;
rom[46267] = 12'h111;
rom[46268] = 12'h111;
rom[46269] = 12'h111;
rom[46270] = 12'h111;
rom[46271] = 12'h111;
rom[46272] = 12'h222;
rom[46273] = 12'h222;
rom[46274] = 12'h222;
rom[46275] = 12'h222;
rom[46276] = 12'h333;
rom[46277] = 12'h444;
rom[46278] = 12'h555;
rom[46279] = 12'h555;
rom[46280] = 12'h555;
rom[46281] = 12'h555;
rom[46282] = 12'h555;
rom[46283] = 12'h555;
rom[46284] = 12'h555;
rom[46285] = 12'h555;
rom[46286] = 12'h666;
rom[46287] = 12'h777;
rom[46288] = 12'h777;
rom[46289] = 12'h788;
rom[46290] = 12'h899;
rom[46291] = 12'h9aa;
rom[46292] = 12'haaa;
rom[46293] = 12'habb;
rom[46294] = 12'hbbb;
rom[46295] = 12'hbbb;
rom[46296] = 12'h988;
rom[46297] = 12'h655;
rom[46298] = 12'h322;
rom[46299] = 12'h211;
rom[46300] = 12'h100;
rom[46301] = 12'h100;
rom[46302] = 12'h100;
rom[46303] = 12'h100;
rom[46304] = 12'h100;
rom[46305] = 12'h100;
rom[46306] = 12'h100;
rom[46307] = 12'h100;
rom[46308] = 12'h100;
rom[46309] = 12'h100;
rom[46310] = 12'h100;
rom[46311] = 12'h100;
rom[46312] = 12'h100;
rom[46313] = 12'h100;
rom[46314] = 12'h100;
rom[46315] = 12'h100;
rom[46316] = 12'h200;
rom[46317] = 12'h200;
rom[46318] = 12'h200;
rom[46319] = 12'h200;
rom[46320] = 12'h200;
rom[46321] = 12'h200;
rom[46322] = 12'h200;
rom[46323] = 12'h200;
rom[46324] = 12'h200;
rom[46325] = 12'h200;
rom[46326] = 12'h200;
rom[46327] = 12'h200;
rom[46328] = 12'h200;
rom[46329] = 12'h200;
rom[46330] = 12'h200;
rom[46331] = 12'h200;
rom[46332] = 12'h200;
rom[46333] = 12'h200;
rom[46334] = 12'h200;
rom[46335] = 12'h200;
rom[46336] = 12'h200;
rom[46337] = 12'h200;
rom[46338] = 12'h300;
rom[46339] = 12'h300;
rom[46340] = 12'h300;
rom[46341] = 12'h400;
rom[46342] = 12'h400;
rom[46343] = 12'h400;
rom[46344] = 12'h510;
rom[46345] = 12'h510;
rom[46346] = 12'h510;
rom[46347] = 12'h510;
rom[46348] = 12'h510;
rom[46349] = 12'h510;
rom[46350] = 12'h520;
rom[46351] = 12'h520;
rom[46352] = 12'h420;
rom[46353] = 12'h520;
rom[46354] = 12'h521;
rom[46355] = 12'h521;
rom[46356] = 12'h532;
rom[46357] = 12'h533;
rom[46358] = 12'h533;
rom[46359] = 12'h544;
rom[46360] = 12'h544;
rom[46361] = 12'h545;
rom[46362] = 12'h655;
rom[46363] = 12'h655;
rom[46364] = 12'h655;
rom[46365] = 12'h665;
rom[46366] = 12'h766;
rom[46367] = 12'h776;
rom[46368] = 12'h777;
rom[46369] = 12'h777;
rom[46370] = 12'h877;
rom[46371] = 12'h877;
rom[46372] = 12'h888;
rom[46373] = 12'h888;
rom[46374] = 12'h988;
rom[46375] = 12'h988;
rom[46376] = 12'h999;
rom[46377] = 12'haaa;
rom[46378] = 12'hbab;
rom[46379] = 12'hcbb;
rom[46380] = 12'hccc;
rom[46381] = 12'hccc;
rom[46382] = 12'hcbc;
rom[46383] = 12'hcbc;
rom[46384] = 12'hbbb;
rom[46385] = 12'hbbb;
rom[46386] = 12'hbbb;
rom[46387] = 12'hbbb;
rom[46388] = 12'haaa;
rom[46389] = 12'haaa;
rom[46390] = 12'haaa;
rom[46391] = 12'haaa;
rom[46392] = 12'h999;
rom[46393] = 12'h999;
rom[46394] = 12'h999;
rom[46395] = 12'haaa;
rom[46396] = 12'haaa;
rom[46397] = 12'haaa;
rom[46398] = 12'haaa;
rom[46399] = 12'hbbb;
rom[46400] = 12'haaa;
rom[46401] = 12'haaa;
rom[46402] = 12'haaa;
rom[46403] = 12'h999;
rom[46404] = 12'h999;
rom[46405] = 12'h999;
rom[46406] = 12'h888;
rom[46407] = 12'h888;
rom[46408] = 12'h777;
rom[46409] = 12'h777;
rom[46410] = 12'h777;
rom[46411] = 12'h666;
rom[46412] = 12'h666;
rom[46413] = 12'h666;
rom[46414] = 12'h666;
rom[46415] = 12'h666;
rom[46416] = 12'h666;
rom[46417] = 12'h666;
rom[46418] = 12'h666;
rom[46419] = 12'h666;
rom[46420] = 12'h666;
rom[46421] = 12'h666;
rom[46422] = 12'h666;
rom[46423] = 12'h666;
rom[46424] = 12'h777;
rom[46425] = 12'h777;
rom[46426] = 12'h777;
rom[46427] = 12'h777;
rom[46428] = 12'h777;
rom[46429] = 12'h777;
rom[46430] = 12'h777;
rom[46431] = 12'h777;
rom[46432] = 12'h777;
rom[46433] = 12'h777;
rom[46434] = 12'h777;
rom[46435] = 12'h777;
rom[46436] = 12'h777;
rom[46437] = 12'h777;
rom[46438] = 12'h777;
rom[46439] = 12'h777;
rom[46440] = 12'h777;
rom[46441] = 12'h777;
rom[46442] = 12'h777;
rom[46443] = 12'h777;
rom[46444] = 12'h777;
rom[46445] = 12'h888;
rom[46446] = 12'h888;
rom[46447] = 12'h888;
rom[46448] = 12'h777;
rom[46449] = 12'h777;
rom[46450] = 12'h888;
rom[46451] = 12'h888;
rom[46452] = 12'h888;
rom[46453] = 12'h888;
rom[46454] = 12'h888;
rom[46455] = 12'h888;
rom[46456] = 12'h999;
rom[46457] = 12'h999;
rom[46458] = 12'h999;
rom[46459] = 12'h999;
rom[46460] = 12'h999;
rom[46461] = 12'haaa;
rom[46462] = 12'haaa;
rom[46463] = 12'haaa;
rom[46464] = 12'haaa;
rom[46465] = 12'haaa;
rom[46466] = 12'haaa;
rom[46467] = 12'haaa;
rom[46468] = 12'haaa;
rom[46469] = 12'h999;
rom[46470] = 12'h888;
rom[46471] = 12'h888;
rom[46472] = 12'h777;
rom[46473] = 12'h777;
rom[46474] = 12'h777;
rom[46475] = 12'h777;
rom[46476] = 12'h777;
rom[46477] = 12'h666;
rom[46478] = 12'h666;
rom[46479] = 12'h666;
rom[46480] = 12'h666;
rom[46481] = 12'h666;
rom[46482] = 12'h666;
rom[46483] = 12'h666;
rom[46484] = 12'h666;
rom[46485] = 12'h666;
rom[46486] = 12'h555;
rom[46487] = 12'h555;
rom[46488] = 12'h555;
rom[46489] = 12'h555;
rom[46490] = 12'h555;
rom[46491] = 12'h555;
rom[46492] = 12'h555;
rom[46493] = 12'h666;
rom[46494] = 12'h666;
rom[46495] = 12'h666;
rom[46496] = 12'h777;
rom[46497] = 12'h666;
rom[46498] = 12'h666;
rom[46499] = 12'h555;
rom[46500] = 12'h555;
rom[46501] = 12'h444;
rom[46502] = 12'h444;
rom[46503] = 12'h444;
rom[46504] = 12'h444;
rom[46505] = 12'h333;
rom[46506] = 12'h333;
rom[46507] = 12'h333;
rom[46508] = 12'h333;
rom[46509] = 12'h333;
rom[46510] = 12'h333;
rom[46511] = 12'h222;
rom[46512] = 12'h111;
rom[46513] = 12'h111;
rom[46514] = 12'h111;
rom[46515] = 12'h111;
rom[46516] = 12'h  0;
rom[46517] = 12'h  0;
rom[46518] = 12'h  0;
rom[46519] = 12'h  0;
rom[46520] = 12'h  0;
rom[46521] = 12'h  0;
rom[46522] = 12'h  0;
rom[46523] = 12'h  0;
rom[46524] = 12'h  0;
rom[46525] = 12'h  0;
rom[46526] = 12'h  0;
rom[46527] = 12'h  0;
rom[46528] = 12'h  0;
rom[46529] = 12'h  0;
rom[46530] = 12'h  0;
rom[46531] = 12'h  0;
rom[46532] = 12'h  0;
rom[46533] = 12'h  0;
rom[46534] = 12'h  0;
rom[46535] = 12'h  0;
rom[46536] = 12'h  0;
rom[46537] = 12'h  0;
rom[46538] = 12'h  0;
rom[46539] = 12'h  0;
rom[46540] = 12'h  0;
rom[46541] = 12'h  0;
rom[46542] = 12'h  0;
rom[46543] = 12'h  0;
rom[46544] = 12'h  0;
rom[46545] = 12'h  0;
rom[46546] = 12'h  0;
rom[46547] = 12'h111;
rom[46548] = 12'h111;
rom[46549] = 12'h111;
rom[46550] = 12'h111;
rom[46551] = 12'h111;
rom[46552] = 12'h111;
rom[46553] = 12'h111;
rom[46554] = 12'h111;
rom[46555] = 12'h111;
rom[46556] = 12'h111;
rom[46557] = 12'h111;
rom[46558] = 12'h111;
rom[46559] = 12'h111;
rom[46560] = 12'h111;
rom[46561] = 12'h111;
rom[46562] = 12'h111;
rom[46563] = 12'h111;
rom[46564] = 12'h111;
rom[46565] = 12'h111;
rom[46566] = 12'h111;
rom[46567] = 12'h111;
rom[46568] = 12'h222;
rom[46569] = 12'h111;
rom[46570] = 12'h111;
rom[46571] = 12'h111;
rom[46572] = 12'h111;
rom[46573] = 12'h111;
rom[46574] = 12'h111;
rom[46575] = 12'h111;
rom[46576] = 12'h111;
rom[46577] = 12'h111;
rom[46578] = 12'h222;
rom[46579] = 12'h222;
rom[46580] = 12'h222;
rom[46581] = 12'h222;
rom[46582] = 12'h222;
rom[46583] = 12'h222;
rom[46584] = 12'h222;
rom[46585] = 12'h222;
rom[46586] = 12'h222;
rom[46587] = 12'h222;
rom[46588] = 12'h222;
rom[46589] = 12'h222;
rom[46590] = 12'h222;
rom[46591] = 12'h111;
rom[46592] = 12'h111;
rom[46593] = 12'h111;
rom[46594] = 12'h111;
rom[46595] = 12'h111;
rom[46596] = 12'h111;
rom[46597] = 12'h111;
rom[46598] = 12'h111;
rom[46599] = 12'h111;
rom[46600] = 12'h111;
rom[46601] = 12'h111;
rom[46602] = 12'h111;
rom[46603] = 12'h111;
rom[46604] = 12'h111;
rom[46605] = 12'h111;
rom[46606] = 12'h111;
rom[46607] = 12'h111;
rom[46608] = 12'h111;
rom[46609] = 12'h111;
rom[46610] = 12'h222;
rom[46611] = 12'h222;
rom[46612] = 12'h222;
rom[46613] = 12'h222;
rom[46614] = 12'h222;
rom[46615] = 12'h222;
rom[46616] = 12'h222;
rom[46617] = 12'h222;
rom[46618] = 12'h222;
rom[46619] = 12'h222;
rom[46620] = 12'h333;
rom[46621] = 12'h333;
rom[46622] = 12'h333;
rom[46623] = 12'h333;
rom[46624] = 12'h333;
rom[46625] = 12'h222;
rom[46626] = 12'h222;
rom[46627] = 12'h222;
rom[46628] = 12'h333;
rom[46629] = 12'h222;
rom[46630] = 12'h222;
rom[46631] = 12'h222;
rom[46632] = 12'h222;
rom[46633] = 12'h222;
rom[46634] = 12'h111;
rom[46635] = 12'h111;
rom[46636] = 12'h111;
rom[46637] = 12'h111;
rom[46638] = 12'h111;
rom[46639] = 12'h111;
rom[46640] = 12'h111;
rom[46641] = 12'h111;
rom[46642] = 12'h  0;
rom[46643] = 12'h  0;
rom[46644] = 12'h  0;
rom[46645] = 12'h  0;
rom[46646] = 12'h  0;
rom[46647] = 12'h  0;
rom[46648] = 12'h  0;
rom[46649] = 12'h  0;
rom[46650] = 12'h  0;
rom[46651] = 12'h  0;
rom[46652] = 12'h  0;
rom[46653] = 12'h  0;
rom[46654] = 12'h  0;
rom[46655] = 12'h  0;
rom[46656] = 12'h  0;
rom[46657] = 12'h  0;
rom[46658] = 12'h  0;
rom[46659] = 12'h  0;
rom[46660] = 12'h  0;
rom[46661] = 12'h  0;
rom[46662] = 12'h  0;
rom[46663] = 12'h  0;
rom[46664] = 12'h  0;
rom[46665] = 12'h  0;
rom[46666] = 12'h  0;
rom[46667] = 12'h111;
rom[46668] = 12'h111;
rom[46669] = 12'h111;
rom[46670] = 12'h111;
rom[46671] = 12'h111;
rom[46672] = 12'h222;
rom[46673] = 12'h222;
rom[46674] = 12'h222;
rom[46675] = 12'h222;
rom[46676] = 12'h333;
rom[46677] = 12'h444;
rom[46678] = 12'h555;
rom[46679] = 12'h555;
rom[46680] = 12'h555;
rom[46681] = 12'h555;
rom[46682] = 12'h555;
rom[46683] = 12'h555;
rom[46684] = 12'h555;
rom[46685] = 12'h555;
rom[46686] = 12'h666;
rom[46687] = 12'h777;
rom[46688] = 12'h777;
rom[46689] = 12'h787;
rom[46690] = 12'h999;
rom[46691] = 12'haaa;
rom[46692] = 12'haaa;
rom[46693] = 12'haaa;
rom[46694] = 12'haba;
rom[46695] = 12'haba;
rom[46696] = 12'h888;
rom[46697] = 12'h655;
rom[46698] = 12'h333;
rom[46699] = 12'h211;
rom[46700] = 12'h101;
rom[46701] = 12'h100;
rom[46702] = 12'h100;
rom[46703] = 12'h100;
rom[46704] = 12'h  0;
rom[46705] = 12'h  0;
rom[46706] = 12'h  0;
rom[46707] = 12'h  0;
rom[46708] = 12'h  0;
rom[46709] = 12'h  0;
rom[46710] = 12'h100;
rom[46711] = 12'h100;
rom[46712] = 12'h100;
rom[46713] = 12'h100;
rom[46714] = 12'h100;
rom[46715] = 12'h100;
rom[46716] = 12'h100;
rom[46717] = 12'h100;
rom[46718] = 12'h100;
rom[46719] = 12'h200;
rom[46720] = 12'h200;
rom[46721] = 12'h200;
rom[46722] = 12'h200;
rom[46723] = 12'h200;
rom[46724] = 12'h200;
rom[46725] = 12'h200;
rom[46726] = 12'h200;
rom[46727] = 12'h200;
rom[46728] = 12'h200;
rom[46729] = 12'h200;
rom[46730] = 12'h200;
rom[46731] = 12'h200;
rom[46732] = 12'h200;
rom[46733] = 12'h200;
rom[46734] = 12'h200;
rom[46735] = 12'h200;
rom[46736] = 12'h200;
rom[46737] = 12'h200;
rom[46738] = 12'h200;
rom[46739] = 12'h300;
rom[46740] = 12'h300;
rom[46741] = 12'h300;
rom[46742] = 12'h400;
rom[46743] = 12'h400;
rom[46744] = 12'h410;
rom[46745] = 12'h410;
rom[46746] = 12'h410;
rom[46747] = 12'h410;
rom[46748] = 12'h410;
rom[46749] = 12'h420;
rom[46750] = 12'h520;
rom[46751] = 12'h420;
rom[46752] = 12'h420;
rom[46753] = 12'h421;
rom[46754] = 12'h521;
rom[46755] = 12'h532;
rom[46756] = 12'h532;
rom[46757] = 12'h533;
rom[46758] = 12'h544;
rom[46759] = 12'h544;
rom[46760] = 12'h545;
rom[46761] = 12'h555;
rom[46762] = 12'h655;
rom[46763] = 12'h655;
rom[46764] = 12'h666;
rom[46765] = 12'h666;
rom[46766] = 12'h776;
rom[46767] = 12'h777;
rom[46768] = 12'h777;
rom[46769] = 12'h777;
rom[46770] = 12'h877;
rom[46771] = 12'h887;
rom[46772] = 12'h888;
rom[46773] = 12'h888;
rom[46774] = 12'h988;
rom[46775] = 12'h999;
rom[46776] = 12'haaa;
rom[46777] = 12'haaa;
rom[46778] = 12'hbbb;
rom[46779] = 12'hccc;
rom[46780] = 12'hccc;
rom[46781] = 12'hccc;
rom[46782] = 12'hccc;
rom[46783] = 12'hcbc;
rom[46784] = 12'hbbb;
rom[46785] = 12'hbbb;
rom[46786] = 12'hbbb;
rom[46787] = 12'hbbb;
rom[46788] = 12'haaa;
rom[46789] = 12'haaa;
rom[46790] = 12'haaa;
rom[46791] = 12'haaa;
rom[46792] = 12'haaa;
rom[46793] = 12'haaa;
rom[46794] = 12'haaa;
rom[46795] = 12'haaa;
rom[46796] = 12'haaa;
rom[46797] = 12'haaa;
rom[46798] = 12'haaa;
rom[46799] = 12'hbbb;
rom[46800] = 12'haaa;
rom[46801] = 12'h999;
rom[46802] = 12'h999;
rom[46803] = 12'h999;
rom[46804] = 12'h888;
rom[46805] = 12'h888;
rom[46806] = 12'h888;
rom[46807] = 12'h777;
rom[46808] = 12'h777;
rom[46809] = 12'h777;
rom[46810] = 12'h666;
rom[46811] = 12'h666;
rom[46812] = 12'h666;
rom[46813] = 12'h666;
rom[46814] = 12'h666;
rom[46815] = 12'h666;
rom[46816] = 12'h666;
rom[46817] = 12'h666;
rom[46818] = 12'h666;
rom[46819] = 12'h666;
rom[46820] = 12'h666;
rom[46821] = 12'h666;
rom[46822] = 12'h666;
rom[46823] = 12'h666;
rom[46824] = 12'h777;
rom[46825] = 12'h777;
rom[46826] = 12'h777;
rom[46827] = 12'h777;
rom[46828] = 12'h777;
rom[46829] = 12'h777;
rom[46830] = 12'h777;
rom[46831] = 12'h777;
rom[46832] = 12'h777;
rom[46833] = 12'h777;
rom[46834] = 12'h777;
rom[46835] = 12'h777;
rom[46836] = 12'h777;
rom[46837] = 12'h777;
rom[46838] = 12'h777;
rom[46839] = 12'h777;
rom[46840] = 12'h777;
rom[46841] = 12'h777;
rom[46842] = 12'h777;
rom[46843] = 12'h777;
rom[46844] = 12'h777;
rom[46845] = 12'h777;
rom[46846] = 12'h777;
rom[46847] = 12'h777;
rom[46848] = 12'h777;
rom[46849] = 12'h777;
rom[46850] = 12'h888;
rom[46851] = 12'h888;
rom[46852] = 12'h888;
rom[46853] = 12'h888;
rom[46854] = 12'h888;
rom[46855] = 12'h888;
rom[46856] = 12'h999;
rom[46857] = 12'h999;
rom[46858] = 12'h999;
rom[46859] = 12'h999;
rom[46860] = 12'h999;
rom[46861] = 12'h999;
rom[46862] = 12'haaa;
rom[46863] = 12'haaa;
rom[46864] = 12'haaa;
rom[46865] = 12'haaa;
rom[46866] = 12'haaa;
rom[46867] = 12'haaa;
rom[46868] = 12'haaa;
rom[46869] = 12'h999;
rom[46870] = 12'h999;
rom[46871] = 12'h888;
rom[46872] = 12'h888;
rom[46873] = 12'h777;
rom[46874] = 12'h777;
rom[46875] = 12'h777;
rom[46876] = 12'h777;
rom[46877] = 12'h666;
rom[46878] = 12'h666;
rom[46879] = 12'h666;
rom[46880] = 12'h666;
rom[46881] = 12'h666;
rom[46882] = 12'h666;
rom[46883] = 12'h666;
rom[46884] = 12'h666;
rom[46885] = 12'h666;
rom[46886] = 12'h666;
rom[46887] = 12'h555;
rom[46888] = 12'h555;
rom[46889] = 12'h555;
rom[46890] = 12'h555;
rom[46891] = 12'h555;
rom[46892] = 12'h555;
rom[46893] = 12'h666;
rom[46894] = 12'h666;
rom[46895] = 12'h666;
rom[46896] = 12'h777;
rom[46897] = 12'h666;
rom[46898] = 12'h666;
rom[46899] = 12'h555;
rom[46900] = 12'h555;
rom[46901] = 12'h444;
rom[46902] = 12'h444;
rom[46903] = 12'h444;
rom[46904] = 12'h444;
rom[46905] = 12'h444;
rom[46906] = 12'h333;
rom[46907] = 12'h333;
rom[46908] = 12'h333;
rom[46909] = 12'h333;
rom[46910] = 12'h333;
rom[46911] = 12'h333;
rom[46912] = 12'h222;
rom[46913] = 12'h111;
rom[46914] = 12'h111;
rom[46915] = 12'h111;
rom[46916] = 12'h111;
rom[46917] = 12'h111;
rom[46918] = 12'h  0;
rom[46919] = 12'h  0;
rom[46920] = 12'h  0;
rom[46921] = 12'h  0;
rom[46922] = 12'h  0;
rom[46923] = 12'h  0;
rom[46924] = 12'h  0;
rom[46925] = 12'h  0;
rom[46926] = 12'h  0;
rom[46927] = 12'h  0;
rom[46928] = 12'h  0;
rom[46929] = 12'h  0;
rom[46930] = 12'h  0;
rom[46931] = 12'h  0;
rom[46932] = 12'h  0;
rom[46933] = 12'h  0;
rom[46934] = 12'h  0;
rom[46935] = 12'h  0;
rom[46936] = 12'h  0;
rom[46937] = 12'h  0;
rom[46938] = 12'h  0;
rom[46939] = 12'h  0;
rom[46940] = 12'h  0;
rom[46941] = 12'h  0;
rom[46942] = 12'h  0;
rom[46943] = 12'h  0;
rom[46944] = 12'h  0;
rom[46945] = 12'h  0;
rom[46946] = 12'h  0;
rom[46947] = 12'h  0;
rom[46948] = 12'h111;
rom[46949] = 12'h111;
rom[46950] = 12'h111;
rom[46951] = 12'h111;
rom[46952] = 12'h111;
rom[46953] = 12'h111;
rom[46954] = 12'h111;
rom[46955] = 12'h111;
rom[46956] = 12'h111;
rom[46957] = 12'h111;
rom[46958] = 12'h111;
rom[46959] = 12'h111;
rom[46960] = 12'h111;
rom[46961] = 12'h111;
rom[46962] = 12'h111;
rom[46963] = 12'h111;
rom[46964] = 12'h111;
rom[46965] = 12'h111;
rom[46966] = 12'h111;
rom[46967] = 12'h111;
rom[46968] = 12'h111;
rom[46969] = 12'h111;
rom[46970] = 12'h111;
rom[46971] = 12'h111;
rom[46972] = 12'h111;
rom[46973] = 12'h111;
rom[46974] = 12'h111;
rom[46975] = 12'h111;
rom[46976] = 12'h222;
rom[46977] = 12'h222;
rom[46978] = 12'h222;
rom[46979] = 12'h222;
rom[46980] = 12'h222;
rom[46981] = 12'h222;
rom[46982] = 12'h222;
rom[46983] = 12'h222;
rom[46984] = 12'h222;
rom[46985] = 12'h222;
rom[46986] = 12'h222;
rom[46987] = 12'h222;
rom[46988] = 12'h222;
rom[46989] = 12'h111;
rom[46990] = 12'h111;
rom[46991] = 12'h111;
rom[46992] = 12'h111;
rom[46993] = 12'h111;
rom[46994] = 12'h111;
rom[46995] = 12'h111;
rom[46996] = 12'h111;
rom[46997] = 12'h111;
rom[46998] = 12'h111;
rom[46999] = 12'h111;
rom[47000] = 12'h111;
rom[47001] = 12'h111;
rom[47002] = 12'h111;
rom[47003] = 12'h  0;
rom[47004] = 12'h  0;
rom[47005] = 12'h111;
rom[47006] = 12'h111;
rom[47007] = 12'h111;
rom[47008] = 12'h111;
rom[47009] = 12'h111;
rom[47010] = 12'h111;
rom[47011] = 12'h222;
rom[47012] = 12'h222;
rom[47013] = 12'h222;
rom[47014] = 12'h222;
rom[47015] = 12'h222;
rom[47016] = 12'h222;
rom[47017] = 12'h222;
rom[47018] = 12'h222;
rom[47019] = 12'h222;
rom[47020] = 12'h222;
rom[47021] = 12'h333;
rom[47022] = 12'h222;
rom[47023] = 12'h222;
rom[47024] = 12'h333;
rom[47025] = 12'h222;
rom[47026] = 12'h222;
rom[47027] = 12'h222;
rom[47028] = 12'h333;
rom[47029] = 12'h333;
rom[47030] = 12'h222;
rom[47031] = 12'h222;
rom[47032] = 12'h222;
rom[47033] = 12'h222;
rom[47034] = 12'h111;
rom[47035] = 12'h111;
rom[47036] = 12'h111;
rom[47037] = 12'h111;
rom[47038] = 12'h111;
rom[47039] = 12'h111;
rom[47040] = 12'h  0;
rom[47041] = 12'h  0;
rom[47042] = 12'h  0;
rom[47043] = 12'h  0;
rom[47044] = 12'h  0;
rom[47045] = 12'h  0;
rom[47046] = 12'h  0;
rom[47047] = 12'h  0;
rom[47048] = 12'h  0;
rom[47049] = 12'h  0;
rom[47050] = 12'h  0;
rom[47051] = 12'h  0;
rom[47052] = 12'h  0;
rom[47053] = 12'h  0;
rom[47054] = 12'h  0;
rom[47055] = 12'h  0;
rom[47056] = 12'h  0;
rom[47057] = 12'h  0;
rom[47058] = 12'h  0;
rom[47059] = 12'h  0;
rom[47060] = 12'h  0;
rom[47061] = 12'h  0;
rom[47062] = 12'h  0;
rom[47063] = 12'h  0;
rom[47064] = 12'h  0;
rom[47065] = 12'h  0;
rom[47066] = 12'h111;
rom[47067] = 12'h111;
rom[47068] = 12'h111;
rom[47069] = 12'h111;
rom[47070] = 12'h111;
rom[47071] = 12'h111;
rom[47072] = 12'h222;
rom[47073] = 12'h222;
rom[47074] = 12'h222;
rom[47075] = 12'h222;
rom[47076] = 12'h333;
rom[47077] = 12'h444;
rom[47078] = 12'h555;
rom[47079] = 12'h555;
rom[47080] = 12'h555;
rom[47081] = 12'h555;
rom[47082] = 12'h555;
rom[47083] = 12'h555;
rom[47084] = 12'h555;
rom[47085] = 12'h555;
rom[47086] = 12'h666;
rom[47087] = 12'h777;
rom[47088] = 12'h777;
rom[47089] = 12'h787;
rom[47090] = 12'h999;
rom[47091] = 12'haaa;
rom[47092] = 12'haaa;
rom[47093] = 12'haaa;
rom[47094] = 12'haaa;
rom[47095] = 12'haaa;
rom[47096] = 12'h888;
rom[47097] = 12'h655;
rom[47098] = 12'h433;
rom[47099] = 12'h222;
rom[47100] = 12'h211;
rom[47101] = 12'h100;
rom[47102] = 12'h100;
rom[47103] = 12'h100;
rom[47104] = 12'h  0;
rom[47105] = 12'h  0;
rom[47106] = 12'h  0;
rom[47107] = 12'h  0;
rom[47108] = 12'h  0;
rom[47109] = 12'h  0;
rom[47110] = 12'h  0;
rom[47111] = 12'h100;
rom[47112] = 12'h100;
rom[47113] = 12'h100;
rom[47114] = 12'h100;
rom[47115] = 12'h100;
rom[47116] = 12'h100;
rom[47117] = 12'h100;
rom[47118] = 12'h100;
rom[47119] = 12'h100;
rom[47120] = 12'h100;
rom[47121] = 12'h100;
rom[47122] = 12'h100;
rom[47123] = 12'h100;
rom[47124] = 12'h200;
rom[47125] = 12'h200;
rom[47126] = 12'h200;
rom[47127] = 12'h200;
rom[47128] = 12'h200;
rom[47129] = 12'h200;
rom[47130] = 12'h200;
rom[47131] = 12'h200;
rom[47132] = 12'h200;
rom[47133] = 12'h200;
rom[47134] = 12'h200;
rom[47135] = 12'h200;
rom[47136] = 12'h200;
rom[47137] = 12'h200;
rom[47138] = 12'h200;
rom[47139] = 12'h300;
rom[47140] = 12'h300;
rom[47141] = 12'h300;
rom[47142] = 12'h400;
rom[47143] = 12'h400;
rom[47144] = 12'h410;
rom[47145] = 12'h410;
rom[47146] = 12'h410;
rom[47147] = 12'h410;
rom[47148] = 12'h410;
rom[47149] = 12'h420;
rom[47150] = 12'h421;
rom[47151] = 12'h421;
rom[47152] = 12'h421;
rom[47153] = 12'h431;
rom[47154] = 12'h532;
rom[47155] = 12'h533;
rom[47156] = 12'h543;
rom[47157] = 12'h544;
rom[47158] = 12'h545;
rom[47159] = 12'h655;
rom[47160] = 12'h655;
rom[47161] = 12'h655;
rom[47162] = 12'h656;
rom[47163] = 12'h666;
rom[47164] = 12'h666;
rom[47165] = 12'h666;
rom[47166] = 12'h776;
rom[47167] = 12'h777;
rom[47168] = 12'h777;
rom[47169] = 12'h777;
rom[47170] = 12'h877;
rom[47171] = 12'h887;
rom[47172] = 12'h888;
rom[47173] = 12'h888;
rom[47174] = 12'h999;
rom[47175] = 12'h999;
rom[47176] = 12'haaa;
rom[47177] = 12'hbbb;
rom[47178] = 12'hcbb;
rom[47179] = 12'hccc;
rom[47180] = 12'hccc;
rom[47181] = 12'hccc;
rom[47182] = 12'hcbc;
rom[47183] = 12'hbbb;
rom[47184] = 12'hbbb;
rom[47185] = 12'hbbb;
rom[47186] = 12'hbbb;
rom[47187] = 12'hbbb;
rom[47188] = 12'haaa;
rom[47189] = 12'haaa;
rom[47190] = 12'haaa;
rom[47191] = 12'haaa;
rom[47192] = 12'haaa;
rom[47193] = 12'haaa;
rom[47194] = 12'haaa;
rom[47195] = 12'haaa;
rom[47196] = 12'haaa;
rom[47197] = 12'haaa;
rom[47198] = 12'haaa;
rom[47199] = 12'hbbb;
rom[47200] = 12'h999;
rom[47201] = 12'h999;
rom[47202] = 12'h999;
rom[47203] = 12'h888;
rom[47204] = 12'h888;
rom[47205] = 12'h888;
rom[47206] = 12'h777;
rom[47207] = 12'h777;
rom[47208] = 12'h777;
rom[47209] = 12'h777;
rom[47210] = 12'h666;
rom[47211] = 12'h666;
rom[47212] = 12'h666;
rom[47213] = 12'h666;
rom[47214] = 12'h666;
rom[47215] = 12'h666;
rom[47216] = 12'h666;
rom[47217] = 12'h666;
rom[47218] = 12'h666;
rom[47219] = 12'h666;
rom[47220] = 12'h666;
rom[47221] = 12'h666;
rom[47222] = 12'h777;
rom[47223] = 12'h777;
rom[47224] = 12'h777;
rom[47225] = 12'h777;
rom[47226] = 12'h777;
rom[47227] = 12'h777;
rom[47228] = 12'h777;
rom[47229] = 12'h777;
rom[47230] = 12'h777;
rom[47231] = 12'h777;
rom[47232] = 12'h777;
rom[47233] = 12'h777;
rom[47234] = 12'h777;
rom[47235] = 12'h777;
rom[47236] = 12'h777;
rom[47237] = 12'h777;
rom[47238] = 12'h777;
rom[47239] = 12'h777;
rom[47240] = 12'h777;
rom[47241] = 12'h777;
rom[47242] = 12'h777;
rom[47243] = 12'h777;
rom[47244] = 12'h777;
rom[47245] = 12'h777;
rom[47246] = 12'h777;
rom[47247] = 12'h777;
rom[47248] = 12'h777;
rom[47249] = 12'h888;
rom[47250] = 12'h888;
rom[47251] = 12'h888;
rom[47252] = 12'h888;
rom[47253] = 12'h888;
rom[47254] = 12'h888;
rom[47255] = 12'h888;
rom[47256] = 12'h999;
rom[47257] = 12'h999;
rom[47258] = 12'h999;
rom[47259] = 12'h999;
rom[47260] = 12'h999;
rom[47261] = 12'h999;
rom[47262] = 12'haaa;
rom[47263] = 12'haaa;
rom[47264] = 12'haaa;
rom[47265] = 12'haaa;
rom[47266] = 12'haaa;
rom[47267] = 12'haaa;
rom[47268] = 12'haaa;
rom[47269] = 12'h999;
rom[47270] = 12'h999;
rom[47271] = 12'h888;
rom[47272] = 12'h888;
rom[47273] = 12'h888;
rom[47274] = 12'h777;
rom[47275] = 12'h777;
rom[47276] = 12'h777;
rom[47277] = 12'h777;
rom[47278] = 12'h666;
rom[47279] = 12'h666;
rom[47280] = 12'h666;
rom[47281] = 12'h666;
rom[47282] = 12'h666;
rom[47283] = 12'h666;
rom[47284] = 12'h666;
rom[47285] = 12'h666;
rom[47286] = 12'h666;
rom[47287] = 12'h555;
rom[47288] = 12'h555;
rom[47289] = 12'h555;
rom[47290] = 12'h555;
rom[47291] = 12'h555;
rom[47292] = 12'h555;
rom[47293] = 12'h666;
rom[47294] = 12'h666;
rom[47295] = 12'h666;
rom[47296] = 12'h777;
rom[47297] = 12'h666;
rom[47298] = 12'h666;
rom[47299] = 12'h666;
rom[47300] = 12'h555;
rom[47301] = 12'h555;
rom[47302] = 12'h555;
rom[47303] = 12'h444;
rom[47304] = 12'h444;
rom[47305] = 12'h444;
rom[47306] = 12'h444;
rom[47307] = 12'h444;
rom[47308] = 12'h444;
rom[47309] = 12'h333;
rom[47310] = 12'h333;
rom[47311] = 12'h333;
rom[47312] = 12'h222;
rom[47313] = 12'h222;
rom[47314] = 12'h222;
rom[47315] = 12'h111;
rom[47316] = 12'h111;
rom[47317] = 12'h111;
rom[47318] = 12'h111;
rom[47319] = 12'h  0;
rom[47320] = 12'h  0;
rom[47321] = 12'h  0;
rom[47322] = 12'h  0;
rom[47323] = 12'h  0;
rom[47324] = 12'h  0;
rom[47325] = 12'h  0;
rom[47326] = 12'h  0;
rom[47327] = 12'h  0;
rom[47328] = 12'h  0;
rom[47329] = 12'h  0;
rom[47330] = 12'h  0;
rom[47331] = 12'h  0;
rom[47332] = 12'h  0;
rom[47333] = 12'h  0;
rom[47334] = 12'h  0;
rom[47335] = 12'h  0;
rom[47336] = 12'h  0;
rom[47337] = 12'h  0;
rom[47338] = 12'h  0;
rom[47339] = 12'h  0;
rom[47340] = 12'h  0;
rom[47341] = 12'h  0;
rom[47342] = 12'h  0;
rom[47343] = 12'h  0;
rom[47344] = 12'h  0;
rom[47345] = 12'h  0;
rom[47346] = 12'h  0;
rom[47347] = 12'h  0;
rom[47348] = 12'h  0;
rom[47349] = 12'h111;
rom[47350] = 12'h111;
rom[47351] = 12'h111;
rom[47352] = 12'h111;
rom[47353] = 12'h111;
rom[47354] = 12'h111;
rom[47355] = 12'h111;
rom[47356] = 12'h111;
rom[47357] = 12'h111;
rom[47358] = 12'h111;
rom[47359] = 12'h111;
rom[47360] = 12'h111;
rom[47361] = 12'h111;
rom[47362] = 12'h111;
rom[47363] = 12'h111;
rom[47364] = 12'h111;
rom[47365] = 12'h111;
rom[47366] = 12'h111;
rom[47367] = 12'h111;
rom[47368] = 12'h111;
rom[47369] = 12'h111;
rom[47370] = 12'h111;
rom[47371] = 12'h111;
rom[47372] = 12'h111;
rom[47373] = 12'h111;
rom[47374] = 12'h111;
rom[47375] = 12'h222;
rom[47376] = 12'h222;
rom[47377] = 12'h222;
rom[47378] = 12'h222;
rom[47379] = 12'h222;
rom[47380] = 12'h222;
rom[47381] = 12'h222;
rom[47382] = 12'h222;
rom[47383] = 12'h111;
rom[47384] = 12'h222;
rom[47385] = 12'h222;
rom[47386] = 12'h222;
rom[47387] = 12'h222;
rom[47388] = 12'h111;
rom[47389] = 12'h111;
rom[47390] = 12'h111;
rom[47391] = 12'h111;
rom[47392] = 12'h111;
rom[47393] = 12'h111;
rom[47394] = 12'h111;
rom[47395] = 12'h111;
rom[47396] = 12'h  0;
rom[47397] = 12'h  0;
rom[47398] = 12'h  0;
rom[47399] = 12'h  0;
rom[47400] = 12'h  0;
rom[47401] = 12'h  0;
rom[47402] = 12'h  0;
rom[47403] = 12'h  0;
rom[47404] = 12'h  0;
rom[47405] = 12'h  0;
rom[47406] = 12'h  0;
rom[47407] = 12'h  0;
rom[47408] = 12'h111;
rom[47409] = 12'h111;
rom[47410] = 12'h111;
rom[47411] = 12'h111;
rom[47412] = 12'h111;
rom[47413] = 12'h111;
rom[47414] = 12'h111;
rom[47415] = 12'h111;
rom[47416] = 12'h222;
rom[47417] = 12'h222;
rom[47418] = 12'h222;
rom[47419] = 12'h222;
rom[47420] = 12'h222;
rom[47421] = 12'h222;
rom[47422] = 12'h222;
rom[47423] = 12'h222;
rom[47424] = 12'h222;
rom[47425] = 12'h222;
rom[47426] = 12'h222;
rom[47427] = 12'h222;
rom[47428] = 12'h222;
rom[47429] = 12'h222;
rom[47430] = 12'h222;
rom[47431] = 12'h222;
rom[47432] = 12'h222;
rom[47433] = 12'h111;
rom[47434] = 12'h111;
rom[47435] = 12'h111;
rom[47436] = 12'h111;
rom[47437] = 12'h111;
rom[47438] = 12'h111;
rom[47439] = 12'h111;
rom[47440] = 12'h  0;
rom[47441] = 12'h  0;
rom[47442] = 12'h  0;
rom[47443] = 12'h  0;
rom[47444] = 12'h  0;
rom[47445] = 12'h  0;
rom[47446] = 12'h  0;
rom[47447] = 12'h  0;
rom[47448] = 12'h  0;
rom[47449] = 12'h  0;
rom[47450] = 12'h  0;
rom[47451] = 12'h  0;
rom[47452] = 12'h  0;
rom[47453] = 12'h  0;
rom[47454] = 12'h  0;
rom[47455] = 12'h  0;
rom[47456] = 12'h  0;
rom[47457] = 12'h  0;
rom[47458] = 12'h  0;
rom[47459] = 12'h  0;
rom[47460] = 12'h  0;
rom[47461] = 12'h  0;
rom[47462] = 12'h  0;
rom[47463] = 12'h  0;
rom[47464] = 12'h  0;
rom[47465] = 12'h  0;
rom[47466] = 12'h111;
rom[47467] = 12'h111;
rom[47468] = 12'h111;
rom[47469] = 12'h111;
rom[47470] = 12'h111;
rom[47471] = 12'h111;
rom[47472] = 12'h222;
rom[47473] = 12'h222;
rom[47474] = 12'h222;
rom[47475] = 12'h222;
rom[47476] = 12'h333;
rom[47477] = 12'h555;
rom[47478] = 12'h555;
rom[47479] = 12'h555;
rom[47480] = 12'h555;
rom[47481] = 12'h555;
rom[47482] = 12'h555;
rom[47483] = 12'h555;
rom[47484] = 12'h555;
rom[47485] = 12'h555;
rom[47486] = 12'h666;
rom[47487] = 12'h777;
rom[47488] = 12'h777;
rom[47489] = 12'h888;
rom[47490] = 12'h999;
rom[47491] = 12'h999;
rom[47492] = 12'h9aa;
rom[47493] = 12'h9aa;
rom[47494] = 12'h9aa;
rom[47495] = 12'haaa;
rom[47496] = 12'h888;
rom[47497] = 12'h666;
rom[47498] = 12'h433;
rom[47499] = 12'h322;
rom[47500] = 12'h211;
rom[47501] = 12'h100;
rom[47502] = 12'h100;
rom[47503] = 12'h100;
rom[47504] = 12'h  0;
rom[47505] = 12'h  0;
rom[47506] = 12'h  0;
rom[47507] = 12'h  0;
rom[47508] = 12'h  0;
rom[47509] = 12'h  0;
rom[47510] = 12'h100;
rom[47511] = 12'h100;
rom[47512] = 12'h100;
rom[47513] = 12'h100;
rom[47514] = 12'h100;
rom[47515] = 12'h100;
rom[47516] = 12'h100;
rom[47517] = 12'h100;
rom[47518] = 12'h100;
rom[47519] = 12'h100;
rom[47520] = 12'h100;
rom[47521] = 12'h200;
rom[47522] = 12'h200;
rom[47523] = 12'h200;
rom[47524] = 12'h200;
rom[47525] = 12'h200;
rom[47526] = 12'h200;
rom[47527] = 12'h200;
rom[47528] = 12'h200;
rom[47529] = 12'h200;
rom[47530] = 12'h200;
rom[47531] = 12'h200;
rom[47532] = 12'h200;
rom[47533] = 12'h200;
rom[47534] = 12'h200;
rom[47535] = 12'h200;
rom[47536] = 12'h200;
rom[47537] = 12'h200;
rom[47538] = 12'h200;
rom[47539] = 12'h200;
rom[47540] = 12'h300;
rom[47541] = 12'h300;
rom[47542] = 12'h300;
rom[47543] = 12'h410;
rom[47544] = 12'h410;
rom[47545] = 12'h410;
rom[47546] = 12'h410;
rom[47547] = 12'h410;
rom[47548] = 12'h421;
rom[47549] = 12'h421;
rom[47550] = 12'h421;
rom[47551] = 12'h421;
rom[47552] = 12'h532;
rom[47553] = 12'h532;
rom[47554] = 12'h543;
rom[47555] = 12'h543;
rom[47556] = 12'h544;
rom[47557] = 12'h544;
rom[47558] = 12'h655;
rom[47559] = 12'h655;
rom[47560] = 12'h655;
rom[47561] = 12'h656;
rom[47562] = 12'h656;
rom[47563] = 12'h666;
rom[47564] = 12'h666;
rom[47565] = 12'h666;
rom[47566] = 12'h777;
rom[47567] = 12'h777;
rom[47568] = 12'h777;
rom[47569] = 12'h777;
rom[47570] = 12'h877;
rom[47571] = 12'h888;
rom[47572] = 12'h888;
rom[47573] = 12'h989;
rom[47574] = 12'h999;
rom[47575] = 12'haaa;
rom[47576] = 12'hbbb;
rom[47577] = 12'hbbb;
rom[47578] = 12'hccc;
rom[47579] = 12'hccc;
rom[47580] = 12'hdcc;
rom[47581] = 12'hccc;
rom[47582] = 12'hccc;
rom[47583] = 12'hbbb;
rom[47584] = 12'hbbb;
rom[47585] = 12'hbbb;
rom[47586] = 12'hbbb;
rom[47587] = 12'hbbb;
rom[47588] = 12'haaa;
rom[47589] = 12'haaa;
rom[47590] = 12'haaa;
rom[47591] = 12'haaa;
rom[47592] = 12'haaa;
rom[47593] = 12'haaa;
rom[47594] = 12'haaa;
rom[47595] = 12'haaa;
rom[47596] = 12'haaa;
rom[47597] = 12'haaa;
rom[47598] = 12'haaa;
rom[47599] = 12'hbbb;
rom[47600] = 12'h999;
rom[47601] = 12'h999;
rom[47602] = 12'h999;
rom[47603] = 12'h999;
rom[47604] = 12'h888;
rom[47605] = 12'h888;
rom[47606] = 12'h888;
rom[47607] = 12'h777;
rom[47608] = 12'h777;
rom[47609] = 12'h777;
rom[47610] = 12'h666;
rom[47611] = 12'h666;
rom[47612] = 12'h666;
rom[47613] = 12'h666;
rom[47614] = 12'h666;
rom[47615] = 12'h666;
rom[47616] = 12'h777;
rom[47617] = 12'h666;
rom[47618] = 12'h666;
rom[47619] = 12'h666;
rom[47620] = 12'h666;
rom[47621] = 12'h666;
rom[47622] = 12'h777;
rom[47623] = 12'h777;
rom[47624] = 12'h777;
rom[47625] = 12'h777;
rom[47626] = 12'h777;
rom[47627] = 12'h777;
rom[47628] = 12'h777;
rom[47629] = 12'h777;
rom[47630] = 12'h777;
rom[47631] = 12'h777;
rom[47632] = 12'h777;
rom[47633] = 12'h777;
rom[47634] = 12'h777;
rom[47635] = 12'h777;
rom[47636] = 12'h777;
rom[47637] = 12'h777;
rom[47638] = 12'h777;
rom[47639] = 12'h888;
rom[47640] = 12'h777;
rom[47641] = 12'h777;
rom[47642] = 12'h777;
rom[47643] = 12'h777;
rom[47644] = 12'h777;
rom[47645] = 12'h777;
rom[47646] = 12'h777;
rom[47647] = 12'h777;
rom[47648] = 12'h777;
rom[47649] = 12'h888;
rom[47650] = 12'h888;
rom[47651] = 12'h888;
rom[47652] = 12'h888;
rom[47653] = 12'h888;
rom[47654] = 12'h888;
rom[47655] = 12'h888;
rom[47656] = 12'h999;
rom[47657] = 12'h999;
rom[47658] = 12'h999;
rom[47659] = 12'h999;
rom[47660] = 12'h999;
rom[47661] = 12'h999;
rom[47662] = 12'h999;
rom[47663] = 12'h999;
rom[47664] = 12'haaa;
rom[47665] = 12'haaa;
rom[47666] = 12'haaa;
rom[47667] = 12'haaa;
rom[47668] = 12'haaa;
rom[47669] = 12'h999;
rom[47670] = 12'h999;
rom[47671] = 12'h888;
rom[47672] = 12'h888;
rom[47673] = 12'h888;
rom[47674] = 12'h777;
rom[47675] = 12'h777;
rom[47676] = 12'h777;
rom[47677] = 12'h777;
rom[47678] = 12'h777;
rom[47679] = 12'h666;
rom[47680] = 12'h666;
rom[47681] = 12'h666;
rom[47682] = 12'h666;
rom[47683] = 12'h666;
rom[47684] = 12'h666;
rom[47685] = 12'h666;
rom[47686] = 12'h555;
rom[47687] = 12'h555;
rom[47688] = 12'h555;
rom[47689] = 12'h555;
rom[47690] = 12'h555;
rom[47691] = 12'h555;
rom[47692] = 12'h555;
rom[47693] = 12'h666;
rom[47694] = 12'h666;
rom[47695] = 12'h666;
rom[47696] = 12'h666;
rom[47697] = 12'h666;
rom[47698] = 12'h666;
rom[47699] = 12'h666;
rom[47700] = 12'h666;
rom[47701] = 12'h555;
rom[47702] = 12'h555;
rom[47703] = 12'h444;
rom[47704] = 12'h444;
rom[47705] = 12'h444;
rom[47706] = 12'h444;
rom[47707] = 12'h444;
rom[47708] = 12'h444;
rom[47709] = 12'h333;
rom[47710] = 12'h333;
rom[47711] = 12'h333;
rom[47712] = 12'h333;
rom[47713] = 12'h333;
rom[47714] = 12'h222;
rom[47715] = 12'h111;
rom[47716] = 12'h111;
rom[47717] = 12'h111;
rom[47718] = 12'h111;
rom[47719] = 12'h111;
rom[47720] = 12'h  0;
rom[47721] = 12'h  0;
rom[47722] = 12'h  0;
rom[47723] = 12'h  0;
rom[47724] = 12'h  0;
rom[47725] = 12'h  0;
rom[47726] = 12'h  0;
rom[47727] = 12'h  0;
rom[47728] = 12'h  0;
rom[47729] = 12'h  0;
rom[47730] = 12'h  0;
rom[47731] = 12'h  0;
rom[47732] = 12'h  0;
rom[47733] = 12'h  0;
rom[47734] = 12'h  0;
rom[47735] = 12'h  0;
rom[47736] = 12'h  0;
rom[47737] = 12'h  0;
rom[47738] = 12'h  0;
rom[47739] = 12'h  0;
rom[47740] = 12'h  0;
rom[47741] = 12'h  0;
rom[47742] = 12'h  0;
rom[47743] = 12'h  0;
rom[47744] = 12'h  0;
rom[47745] = 12'h  0;
rom[47746] = 12'h  0;
rom[47747] = 12'h  0;
rom[47748] = 12'h  0;
rom[47749] = 12'h  0;
rom[47750] = 12'h111;
rom[47751] = 12'h111;
rom[47752] = 12'h111;
rom[47753] = 12'h111;
rom[47754] = 12'h111;
rom[47755] = 12'h111;
rom[47756] = 12'h111;
rom[47757] = 12'h111;
rom[47758] = 12'h111;
rom[47759] = 12'h111;
rom[47760] = 12'h111;
rom[47761] = 12'h111;
rom[47762] = 12'h111;
rom[47763] = 12'h111;
rom[47764] = 12'h111;
rom[47765] = 12'h111;
rom[47766] = 12'h111;
rom[47767] = 12'h111;
rom[47768] = 12'h111;
rom[47769] = 12'h111;
rom[47770] = 12'h111;
rom[47771] = 12'h111;
rom[47772] = 12'h111;
rom[47773] = 12'h111;
rom[47774] = 12'h222;
rom[47775] = 12'h222;
rom[47776] = 12'h222;
rom[47777] = 12'h222;
rom[47778] = 12'h222;
rom[47779] = 12'h222;
rom[47780] = 12'h222;
rom[47781] = 12'h222;
rom[47782] = 12'h111;
rom[47783] = 12'h111;
rom[47784] = 12'h222;
rom[47785] = 12'h222;
rom[47786] = 12'h222;
rom[47787] = 12'h111;
rom[47788] = 12'h111;
rom[47789] = 12'h111;
rom[47790] = 12'h111;
rom[47791] = 12'h111;
rom[47792] = 12'h111;
rom[47793] = 12'h111;
rom[47794] = 12'h111;
rom[47795] = 12'h  0;
rom[47796] = 12'h  0;
rom[47797] = 12'h  0;
rom[47798] = 12'h  0;
rom[47799] = 12'h  0;
rom[47800] = 12'h111;
rom[47801] = 12'h  0;
rom[47802] = 12'h  0;
rom[47803] = 12'h  0;
rom[47804] = 12'h  0;
rom[47805] = 12'h  0;
rom[47806] = 12'h  0;
rom[47807] = 12'h111;
rom[47808] = 12'h111;
rom[47809] = 12'h111;
rom[47810] = 12'h111;
rom[47811] = 12'h111;
rom[47812] = 12'h111;
rom[47813] = 12'h111;
rom[47814] = 12'h111;
rom[47815] = 12'h111;
rom[47816] = 12'h111;
rom[47817] = 12'h222;
rom[47818] = 12'h222;
rom[47819] = 12'h222;
rom[47820] = 12'h222;
rom[47821] = 12'h222;
rom[47822] = 12'h222;
rom[47823] = 12'h222;
rom[47824] = 12'h222;
rom[47825] = 12'h222;
rom[47826] = 12'h222;
rom[47827] = 12'h222;
rom[47828] = 12'h222;
rom[47829] = 12'h222;
rom[47830] = 12'h222;
rom[47831] = 12'h111;
rom[47832] = 12'h222;
rom[47833] = 12'h111;
rom[47834] = 12'h111;
rom[47835] = 12'h111;
rom[47836] = 12'h111;
rom[47837] = 12'h111;
rom[47838] = 12'h111;
rom[47839] = 12'h  0;
rom[47840] = 12'h  0;
rom[47841] = 12'h  0;
rom[47842] = 12'h  0;
rom[47843] = 12'h  0;
rom[47844] = 12'h  0;
rom[47845] = 12'h  0;
rom[47846] = 12'h  0;
rom[47847] = 12'h  0;
rom[47848] = 12'h  0;
rom[47849] = 12'h  0;
rom[47850] = 12'h  0;
rom[47851] = 12'h  0;
rom[47852] = 12'h  0;
rom[47853] = 12'h  0;
rom[47854] = 12'h  0;
rom[47855] = 12'h  0;
rom[47856] = 12'h  0;
rom[47857] = 12'h  0;
rom[47858] = 12'h  0;
rom[47859] = 12'h  0;
rom[47860] = 12'h  0;
rom[47861] = 12'h  0;
rom[47862] = 12'h  0;
rom[47863] = 12'h  0;
rom[47864] = 12'h  0;
rom[47865] = 12'h  0;
rom[47866] = 12'h111;
rom[47867] = 12'h111;
rom[47868] = 12'h111;
rom[47869] = 12'h111;
rom[47870] = 12'h111;
rom[47871] = 12'h111;
rom[47872] = 12'h222;
rom[47873] = 12'h222;
rom[47874] = 12'h222;
rom[47875] = 12'h222;
rom[47876] = 12'h333;
rom[47877] = 12'h555;
rom[47878] = 12'h555;
rom[47879] = 12'h555;
rom[47880] = 12'h444;
rom[47881] = 12'h444;
rom[47882] = 12'h444;
rom[47883] = 12'h555;
rom[47884] = 12'h555;
rom[47885] = 12'h555;
rom[47886] = 12'h666;
rom[47887] = 12'h777;
rom[47888] = 12'h777;
rom[47889] = 12'h888;
rom[47890] = 12'h999;
rom[47891] = 12'h999;
rom[47892] = 12'h999;
rom[47893] = 12'h999;
rom[47894] = 12'h999;
rom[47895] = 12'h999;
rom[47896] = 12'h888;
rom[47897] = 12'h666;
rom[47898] = 12'h444;
rom[47899] = 12'h322;
rom[47900] = 12'h211;
rom[47901] = 12'h100;
rom[47902] = 12'h100;
rom[47903] = 12'h100;
rom[47904] = 12'h  0;
rom[47905] = 12'h  0;
rom[47906] = 12'h  0;
rom[47907] = 12'h  0;
rom[47908] = 12'h100;
rom[47909] = 12'h100;
rom[47910] = 12'h100;
rom[47911] = 12'h100;
rom[47912] = 12'h100;
rom[47913] = 12'h100;
rom[47914] = 12'h100;
rom[47915] = 12'h100;
rom[47916] = 12'h100;
rom[47917] = 12'h100;
rom[47918] = 12'h100;
rom[47919] = 12'h100;
rom[47920] = 12'h100;
rom[47921] = 12'h200;
rom[47922] = 12'h200;
rom[47923] = 12'h200;
rom[47924] = 12'h200;
rom[47925] = 12'h200;
rom[47926] = 12'h200;
rom[47927] = 12'h200;
rom[47928] = 12'h200;
rom[47929] = 12'h200;
rom[47930] = 12'h200;
rom[47931] = 12'h200;
rom[47932] = 12'h200;
rom[47933] = 12'h200;
rom[47934] = 12'h200;
rom[47935] = 12'h200;
rom[47936] = 12'h200;
rom[47937] = 12'h200;
rom[47938] = 12'h200;
rom[47939] = 12'h200;
rom[47940] = 12'h200;
rom[47941] = 12'h300;
rom[47942] = 12'h310;
rom[47943] = 12'h310;
rom[47944] = 12'h310;
rom[47945] = 12'h310;
rom[47946] = 12'h310;
rom[47947] = 12'h421;
rom[47948] = 12'h421;
rom[47949] = 12'h422;
rom[47950] = 12'h532;
rom[47951] = 12'h532;
rom[47952] = 12'h543;
rom[47953] = 12'h543;
rom[47954] = 12'h544;
rom[47955] = 12'h544;
rom[47956] = 12'h544;
rom[47957] = 12'h555;
rom[47958] = 12'h555;
rom[47959] = 12'h555;
rom[47960] = 12'h556;
rom[47961] = 12'h556;
rom[47962] = 12'h656;
rom[47963] = 12'h666;
rom[47964] = 12'h666;
rom[47965] = 12'h666;
rom[47966] = 12'h777;
rom[47967] = 12'h777;
rom[47968] = 12'h777;
rom[47969] = 12'h877;
rom[47970] = 12'h888;
rom[47971] = 12'h888;
rom[47972] = 12'h888;
rom[47973] = 12'h999;
rom[47974] = 12'haaa;
rom[47975] = 12'haaa;
rom[47976] = 12'hcbb;
rom[47977] = 12'hccc;
rom[47978] = 12'hccc;
rom[47979] = 12'hdcc;
rom[47980] = 12'hdcc;
rom[47981] = 12'hccc;
rom[47982] = 12'hccc;
rom[47983] = 12'hcbb;
rom[47984] = 12'hbbb;
rom[47985] = 12'hbbb;
rom[47986] = 12'hbbb;
rom[47987] = 12'hbbb;
rom[47988] = 12'haaa;
rom[47989] = 12'haaa;
rom[47990] = 12'haaa;
rom[47991] = 12'haaa;
rom[47992] = 12'haaa;
rom[47993] = 12'haaa;
rom[47994] = 12'haaa;
rom[47995] = 12'haaa;
rom[47996] = 12'haaa;
rom[47997] = 12'haaa;
rom[47998] = 12'hbbb;
rom[47999] = 12'hbbb;
rom[48000] = 12'h999;
rom[48001] = 12'h999;
rom[48002] = 12'h999;
rom[48003] = 12'h999;
rom[48004] = 12'h888;
rom[48005] = 12'h888;
rom[48006] = 12'h888;
rom[48007] = 12'h777;
rom[48008] = 12'h777;
rom[48009] = 12'h777;
rom[48010] = 12'h777;
rom[48011] = 12'h777;
rom[48012] = 12'h666;
rom[48013] = 12'h666;
rom[48014] = 12'h666;
rom[48015] = 12'h666;
rom[48016] = 12'h777;
rom[48017] = 12'h777;
rom[48018] = 12'h777;
rom[48019] = 12'h777;
rom[48020] = 12'h777;
rom[48021] = 12'h777;
rom[48022] = 12'h777;
rom[48023] = 12'h777;
rom[48024] = 12'h777;
rom[48025] = 12'h777;
rom[48026] = 12'h777;
rom[48027] = 12'h777;
rom[48028] = 12'h777;
rom[48029] = 12'h888;
rom[48030] = 12'h888;
rom[48031] = 12'h888;
rom[48032] = 12'h888;
rom[48033] = 12'h777;
rom[48034] = 12'h777;
rom[48035] = 12'h777;
rom[48036] = 12'h777;
rom[48037] = 12'h777;
rom[48038] = 12'h777;
rom[48039] = 12'h777;
rom[48040] = 12'h777;
rom[48041] = 12'h777;
rom[48042] = 12'h777;
rom[48043] = 12'h777;
rom[48044] = 12'h777;
rom[48045] = 12'h777;
rom[48046] = 12'h777;
rom[48047] = 12'h777;
rom[48048] = 12'h777;
rom[48049] = 12'h888;
rom[48050] = 12'h888;
rom[48051] = 12'h888;
rom[48052] = 12'h888;
rom[48053] = 12'h888;
rom[48054] = 12'h888;
rom[48055] = 12'h888;
rom[48056] = 12'h999;
rom[48057] = 12'h999;
rom[48058] = 12'h999;
rom[48059] = 12'h999;
rom[48060] = 12'h999;
rom[48061] = 12'h999;
rom[48062] = 12'h999;
rom[48063] = 12'haaa;
rom[48064] = 12'haaa;
rom[48065] = 12'haaa;
rom[48066] = 12'haaa;
rom[48067] = 12'haaa;
rom[48068] = 12'haaa;
rom[48069] = 12'haaa;
rom[48070] = 12'h999;
rom[48071] = 12'h999;
rom[48072] = 12'h999;
rom[48073] = 12'h888;
rom[48074] = 12'h888;
rom[48075] = 12'h777;
rom[48076] = 12'h777;
rom[48077] = 12'h777;
rom[48078] = 12'h777;
rom[48079] = 12'h777;
rom[48080] = 12'h777;
rom[48081] = 12'h666;
rom[48082] = 12'h666;
rom[48083] = 12'h666;
rom[48084] = 12'h666;
rom[48085] = 12'h666;
rom[48086] = 12'h666;
rom[48087] = 12'h666;
rom[48088] = 12'h555;
rom[48089] = 12'h555;
rom[48090] = 12'h555;
rom[48091] = 12'h555;
rom[48092] = 12'h666;
rom[48093] = 12'h666;
rom[48094] = 12'h666;
rom[48095] = 12'h666;
rom[48096] = 12'h666;
rom[48097] = 12'h666;
rom[48098] = 12'h666;
rom[48099] = 12'h666;
rom[48100] = 12'h666;
rom[48101] = 12'h666;
rom[48102] = 12'h555;
rom[48103] = 12'h444;
rom[48104] = 12'h444;
rom[48105] = 12'h444;
rom[48106] = 12'h444;
rom[48107] = 12'h444;
rom[48108] = 12'h444;
rom[48109] = 12'h444;
rom[48110] = 12'h333;
rom[48111] = 12'h333;
rom[48112] = 12'h333;
rom[48113] = 12'h333;
rom[48114] = 12'h333;
rom[48115] = 12'h222;
rom[48116] = 12'h111;
rom[48117] = 12'h111;
rom[48118] = 12'h111;
rom[48119] = 12'h111;
rom[48120] = 12'h111;
rom[48121] = 12'h  0;
rom[48122] = 12'h  0;
rom[48123] = 12'h  0;
rom[48124] = 12'h  0;
rom[48125] = 12'h  0;
rom[48126] = 12'h  0;
rom[48127] = 12'h  0;
rom[48128] = 12'h  0;
rom[48129] = 12'h  0;
rom[48130] = 12'h  0;
rom[48131] = 12'h  0;
rom[48132] = 12'h  0;
rom[48133] = 12'h  0;
rom[48134] = 12'h  0;
rom[48135] = 12'h  0;
rom[48136] = 12'h  0;
rom[48137] = 12'h  0;
rom[48138] = 12'h  0;
rom[48139] = 12'h  0;
rom[48140] = 12'h  0;
rom[48141] = 12'h  0;
rom[48142] = 12'h  0;
rom[48143] = 12'h  0;
rom[48144] = 12'h  0;
rom[48145] = 12'h  0;
rom[48146] = 12'h  0;
rom[48147] = 12'h  0;
rom[48148] = 12'h  0;
rom[48149] = 12'h  0;
rom[48150] = 12'h  0;
rom[48151] = 12'h111;
rom[48152] = 12'h111;
rom[48153] = 12'h111;
rom[48154] = 12'h111;
rom[48155] = 12'h111;
rom[48156] = 12'h111;
rom[48157] = 12'h111;
rom[48158] = 12'h111;
rom[48159] = 12'h111;
rom[48160] = 12'h111;
rom[48161] = 12'h111;
rom[48162] = 12'h111;
rom[48163] = 12'h111;
rom[48164] = 12'h111;
rom[48165] = 12'h111;
rom[48166] = 12'h111;
rom[48167] = 12'h111;
rom[48168] = 12'h111;
rom[48169] = 12'h111;
rom[48170] = 12'h111;
rom[48171] = 12'h222;
rom[48172] = 12'h222;
rom[48173] = 12'h222;
rom[48174] = 12'h222;
rom[48175] = 12'h222;
rom[48176] = 12'h111;
rom[48177] = 12'h111;
rom[48178] = 12'h111;
rom[48179] = 12'h111;
rom[48180] = 12'h111;
rom[48181] = 12'h111;
rom[48182] = 12'h111;
rom[48183] = 12'h111;
rom[48184] = 12'h111;
rom[48185] = 12'h111;
rom[48186] = 12'h111;
rom[48187] = 12'h111;
rom[48188] = 12'h111;
rom[48189] = 12'h111;
rom[48190] = 12'h111;
rom[48191] = 12'h111;
rom[48192] = 12'h111;
rom[48193] = 12'h  0;
rom[48194] = 12'h  0;
rom[48195] = 12'h  0;
rom[48196] = 12'h  0;
rom[48197] = 12'h  0;
rom[48198] = 12'h  0;
rom[48199] = 12'h  0;
rom[48200] = 12'h  0;
rom[48201] = 12'h  0;
rom[48202] = 12'h  0;
rom[48203] = 12'h  0;
rom[48204] = 12'h  0;
rom[48205] = 12'h  0;
rom[48206] = 12'h  0;
rom[48207] = 12'h  0;
rom[48208] = 12'h111;
rom[48209] = 12'h111;
rom[48210] = 12'h111;
rom[48211] = 12'h111;
rom[48212] = 12'h111;
rom[48213] = 12'h111;
rom[48214] = 12'h111;
rom[48215] = 12'h111;
rom[48216] = 12'h222;
rom[48217] = 12'h222;
rom[48218] = 12'h222;
rom[48219] = 12'h222;
rom[48220] = 12'h222;
rom[48221] = 12'h222;
rom[48222] = 12'h222;
rom[48223] = 12'h222;
rom[48224] = 12'h222;
rom[48225] = 12'h222;
rom[48226] = 12'h222;
rom[48227] = 12'h222;
rom[48228] = 12'h222;
rom[48229] = 12'h222;
rom[48230] = 12'h222;
rom[48231] = 12'h111;
rom[48232] = 12'h111;
rom[48233] = 12'h111;
rom[48234] = 12'h111;
rom[48235] = 12'h111;
rom[48236] = 12'h111;
rom[48237] = 12'h  0;
rom[48238] = 12'h  0;
rom[48239] = 12'h  0;
rom[48240] = 12'h  0;
rom[48241] = 12'h  0;
rom[48242] = 12'h  0;
rom[48243] = 12'h  0;
rom[48244] = 12'h  0;
rom[48245] = 12'h  0;
rom[48246] = 12'h  0;
rom[48247] = 12'h  0;
rom[48248] = 12'h  0;
rom[48249] = 12'h  0;
rom[48250] = 12'h  0;
rom[48251] = 12'h  0;
rom[48252] = 12'h  0;
rom[48253] = 12'h  0;
rom[48254] = 12'h  0;
rom[48255] = 12'h  0;
rom[48256] = 12'h  0;
rom[48257] = 12'h  0;
rom[48258] = 12'h  0;
rom[48259] = 12'h  0;
rom[48260] = 12'h  0;
rom[48261] = 12'h  0;
rom[48262] = 12'h  0;
rom[48263] = 12'h  0;
rom[48264] = 12'h  0;
rom[48265] = 12'h  0;
rom[48266] = 12'h  0;
rom[48267] = 12'h  0;
rom[48268] = 12'h111;
rom[48269] = 12'h111;
rom[48270] = 12'h111;
rom[48271] = 12'h111;
rom[48272] = 12'h222;
rom[48273] = 12'h222;
rom[48274] = 12'h222;
rom[48275] = 12'h222;
rom[48276] = 12'h333;
rom[48277] = 12'h555;
rom[48278] = 12'h555;
rom[48279] = 12'h444;
rom[48280] = 12'h444;
rom[48281] = 12'h444;
rom[48282] = 12'h444;
rom[48283] = 12'h555;
rom[48284] = 12'h555;
rom[48285] = 12'h555;
rom[48286] = 12'h666;
rom[48287] = 12'h666;
rom[48288] = 12'h777;
rom[48289] = 12'h888;
rom[48290] = 12'h999;
rom[48291] = 12'h999;
rom[48292] = 12'h888;
rom[48293] = 12'h888;
rom[48294] = 12'h999;
rom[48295] = 12'h9a9;
rom[48296] = 12'h888;
rom[48297] = 12'h666;
rom[48298] = 12'h444;
rom[48299] = 12'h333;
rom[48300] = 12'h322;
rom[48301] = 12'h111;
rom[48302] = 12'h100;
rom[48303] = 12'h100;
rom[48304] = 12'h100;
rom[48305] = 12'h100;
rom[48306] = 12'h100;
rom[48307] = 12'h100;
rom[48308] = 12'h100;
rom[48309] = 12'h100;
rom[48310] = 12'h100;
rom[48311] = 12'h100;
rom[48312] = 12'h100;
rom[48313] = 12'h100;
rom[48314] = 12'h100;
rom[48315] = 12'h100;
rom[48316] = 12'h100;
rom[48317] = 12'h100;
rom[48318] = 12'h100;
rom[48319] = 12'h100;
rom[48320] = 12'h200;
rom[48321] = 12'h200;
rom[48322] = 12'h200;
rom[48323] = 12'h200;
rom[48324] = 12'h200;
rom[48325] = 12'h200;
rom[48326] = 12'h200;
rom[48327] = 12'h200;
rom[48328] = 12'h200;
rom[48329] = 12'h200;
rom[48330] = 12'h200;
rom[48331] = 12'h200;
rom[48332] = 12'h200;
rom[48333] = 12'h200;
rom[48334] = 12'h200;
rom[48335] = 12'h200;
rom[48336] = 12'h100;
rom[48337] = 12'h200;
rom[48338] = 12'h200;
rom[48339] = 12'h200;
rom[48340] = 12'h200;
rom[48341] = 12'h200;
rom[48342] = 12'h310;
rom[48343] = 12'h310;
rom[48344] = 12'h310;
rom[48345] = 12'h310;
rom[48346] = 12'h321;
rom[48347] = 12'h421;
rom[48348] = 12'h422;
rom[48349] = 12'h532;
rom[48350] = 12'h643;
rom[48351] = 12'h644;
rom[48352] = 12'h544;
rom[48353] = 12'h544;
rom[48354] = 12'h554;
rom[48355] = 12'h554;
rom[48356] = 12'h554;
rom[48357] = 12'h555;
rom[48358] = 12'h555;
rom[48359] = 12'h555;
rom[48360] = 12'h555;
rom[48361] = 12'h556;
rom[48362] = 12'h666;
rom[48363] = 12'h666;
rom[48364] = 12'h667;
rom[48365] = 12'h777;
rom[48366] = 12'h777;
rom[48367] = 12'h777;
rom[48368] = 12'h878;
rom[48369] = 12'h888;
rom[48370] = 12'h888;
rom[48371] = 12'h999;
rom[48372] = 12'h999;
rom[48373] = 12'h999;
rom[48374] = 12'haaa;
rom[48375] = 12'hbbb;
rom[48376] = 12'hccc;
rom[48377] = 12'hccc;
rom[48378] = 12'hddd;
rom[48379] = 12'hddd;
rom[48380] = 12'hccc;
rom[48381] = 12'hccc;
rom[48382] = 12'hcbb;
rom[48383] = 12'hbbb;
rom[48384] = 12'hbbb;
rom[48385] = 12'hbbb;
rom[48386] = 12'hbbb;
rom[48387] = 12'hbbb;
rom[48388] = 12'haaa;
rom[48389] = 12'haaa;
rom[48390] = 12'haaa;
rom[48391] = 12'haaa;
rom[48392] = 12'haaa;
rom[48393] = 12'haaa;
rom[48394] = 12'haaa;
rom[48395] = 12'haaa;
rom[48396] = 12'haaa;
rom[48397] = 12'haaa;
rom[48398] = 12'hbbb;
rom[48399] = 12'hbbb;
rom[48400] = 12'haaa;
rom[48401] = 12'h999;
rom[48402] = 12'h999;
rom[48403] = 12'h999;
rom[48404] = 12'h888;
rom[48405] = 12'h888;
rom[48406] = 12'h888;
rom[48407] = 12'h888;
rom[48408] = 12'h777;
rom[48409] = 12'h777;
rom[48410] = 12'h777;
rom[48411] = 12'h777;
rom[48412] = 12'h777;
rom[48413] = 12'h777;
rom[48414] = 12'h777;
rom[48415] = 12'h777;
rom[48416] = 12'h777;
rom[48417] = 12'h777;
rom[48418] = 12'h777;
rom[48419] = 12'h777;
rom[48420] = 12'h777;
rom[48421] = 12'h777;
rom[48422] = 12'h777;
rom[48423] = 12'h777;
rom[48424] = 12'h777;
rom[48425] = 12'h777;
rom[48426] = 12'h777;
rom[48427] = 12'h777;
rom[48428] = 12'h777;
rom[48429] = 12'h888;
rom[48430] = 12'h888;
rom[48431] = 12'h888;
rom[48432] = 12'h888;
rom[48433] = 12'h777;
rom[48434] = 12'h777;
rom[48435] = 12'h777;
rom[48436] = 12'h777;
rom[48437] = 12'h777;
rom[48438] = 12'h777;
rom[48439] = 12'h777;
rom[48440] = 12'h777;
rom[48441] = 12'h777;
rom[48442] = 12'h777;
rom[48443] = 12'h777;
rom[48444] = 12'h777;
rom[48445] = 12'h777;
rom[48446] = 12'h777;
rom[48447] = 12'h777;
rom[48448] = 12'h777;
rom[48449] = 12'h888;
rom[48450] = 12'h888;
rom[48451] = 12'h888;
rom[48452] = 12'h888;
rom[48453] = 12'h888;
rom[48454] = 12'h888;
rom[48455] = 12'h888;
rom[48456] = 12'h999;
rom[48457] = 12'h999;
rom[48458] = 12'h999;
rom[48459] = 12'h999;
rom[48460] = 12'h999;
rom[48461] = 12'h999;
rom[48462] = 12'h999;
rom[48463] = 12'haaa;
rom[48464] = 12'haaa;
rom[48465] = 12'haaa;
rom[48466] = 12'haaa;
rom[48467] = 12'haaa;
rom[48468] = 12'haaa;
rom[48469] = 12'haaa;
rom[48470] = 12'h999;
rom[48471] = 12'h999;
rom[48472] = 12'h999;
rom[48473] = 12'h999;
rom[48474] = 12'h888;
rom[48475] = 12'h888;
rom[48476] = 12'h888;
rom[48477] = 12'h888;
rom[48478] = 12'h777;
rom[48479] = 12'h777;
rom[48480] = 12'h777;
rom[48481] = 12'h666;
rom[48482] = 12'h666;
rom[48483] = 12'h666;
rom[48484] = 12'h666;
rom[48485] = 12'h666;
rom[48486] = 12'h666;
rom[48487] = 12'h666;
rom[48488] = 12'h666;
rom[48489] = 12'h666;
rom[48490] = 12'h666;
rom[48491] = 12'h666;
rom[48492] = 12'h666;
rom[48493] = 12'h666;
rom[48494] = 12'h666;
rom[48495] = 12'h666;
rom[48496] = 12'h666;
rom[48497] = 12'h666;
rom[48498] = 12'h666;
rom[48499] = 12'h666;
rom[48500] = 12'h666;
rom[48501] = 12'h666;
rom[48502] = 12'h555;
rom[48503] = 12'h444;
rom[48504] = 12'h444;
rom[48505] = 12'h444;
rom[48506] = 12'h444;
rom[48507] = 12'h444;
rom[48508] = 12'h444;
rom[48509] = 12'h444;
rom[48510] = 12'h444;
rom[48511] = 12'h444;
rom[48512] = 12'h444;
rom[48513] = 12'h333;
rom[48514] = 12'h333;
rom[48515] = 12'h222;
rom[48516] = 12'h222;
rom[48517] = 12'h222;
rom[48518] = 12'h111;
rom[48519] = 12'h111;
rom[48520] = 12'h111;
rom[48521] = 12'h  0;
rom[48522] = 12'h  0;
rom[48523] = 12'h  0;
rom[48524] = 12'h  0;
rom[48525] = 12'h  0;
rom[48526] = 12'h  0;
rom[48527] = 12'h  0;
rom[48528] = 12'h  0;
rom[48529] = 12'h  0;
rom[48530] = 12'h  0;
rom[48531] = 12'h  0;
rom[48532] = 12'h  0;
rom[48533] = 12'h  0;
rom[48534] = 12'h  0;
rom[48535] = 12'h  0;
rom[48536] = 12'h  0;
rom[48537] = 12'h  0;
rom[48538] = 12'h  0;
rom[48539] = 12'h  0;
rom[48540] = 12'h  0;
rom[48541] = 12'h  0;
rom[48542] = 12'h  0;
rom[48543] = 12'h  0;
rom[48544] = 12'h  0;
rom[48545] = 12'h  0;
rom[48546] = 12'h  0;
rom[48547] = 12'h  0;
rom[48548] = 12'h  0;
rom[48549] = 12'h  0;
rom[48550] = 12'h  0;
rom[48551] = 12'h111;
rom[48552] = 12'h111;
rom[48553] = 12'h111;
rom[48554] = 12'h111;
rom[48555] = 12'h111;
rom[48556] = 12'h111;
rom[48557] = 12'h111;
rom[48558] = 12'h111;
rom[48559] = 12'h111;
rom[48560] = 12'h111;
rom[48561] = 12'h111;
rom[48562] = 12'h111;
rom[48563] = 12'h111;
rom[48564] = 12'h111;
rom[48565] = 12'h111;
rom[48566] = 12'h111;
rom[48567] = 12'h111;
rom[48568] = 12'h111;
rom[48569] = 12'h111;
rom[48570] = 12'h111;
rom[48571] = 12'h111;
rom[48572] = 12'h222;
rom[48573] = 12'h222;
rom[48574] = 12'h111;
rom[48575] = 12'h111;
rom[48576] = 12'h111;
rom[48577] = 12'h111;
rom[48578] = 12'h111;
rom[48579] = 12'h111;
rom[48580] = 12'h111;
rom[48581] = 12'h111;
rom[48582] = 12'h111;
rom[48583] = 12'h111;
rom[48584] = 12'h111;
rom[48585] = 12'h111;
rom[48586] = 12'h111;
rom[48587] = 12'h111;
rom[48588] = 12'h111;
rom[48589] = 12'h111;
rom[48590] = 12'h111;
rom[48591] = 12'h111;
rom[48592] = 12'h  0;
rom[48593] = 12'h  0;
rom[48594] = 12'h  0;
rom[48595] = 12'h  0;
rom[48596] = 12'h  0;
rom[48597] = 12'h  0;
rom[48598] = 12'h  0;
rom[48599] = 12'h  0;
rom[48600] = 12'h  0;
rom[48601] = 12'h  0;
rom[48602] = 12'h  0;
rom[48603] = 12'h  0;
rom[48604] = 12'h  0;
rom[48605] = 12'h  0;
rom[48606] = 12'h  0;
rom[48607] = 12'h  0;
rom[48608] = 12'h111;
rom[48609] = 12'h111;
rom[48610] = 12'h111;
rom[48611] = 12'h111;
rom[48612] = 12'h111;
rom[48613] = 12'h111;
rom[48614] = 12'h111;
rom[48615] = 12'h111;
rom[48616] = 12'h222;
rom[48617] = 12'h222;
rom[48618] = 12'h222;
rom[48619] = 12'h222;
rom[48620] = 12'h222;
rom[48621] = 12'h222;
rom[48622] = 12'h222;
rom[48623] = 12'h222;
rom[48624] = 12'h222;
rom[48625] = 12'h222;
rom[48626] = 12'h222;
rom[48627] = 12'h222;
rom[48628] = 12'h222;
rom[48629] = 12'h222;
rom[48630] = 12'h111;
rom[48631] = 12'h111;
rom[48632] = 12'h111;
rom[48633] = 12'h111;
rom[48634] = 12'h111;
rom[48635] = 12'h111;
rom[48636] = 12'h111;
rom[48637] = 12'h  0;
rom[48638] = 12'h  0;
rom[48639] = 12'h  0;
rom[48640] = 12'h  0;
rom[48641] = 12'h  0;
rom[48642] = 12'h  0;
rom[48643] = 12'h  0;
rom[48644] = 12'h  0;
rom[48645] = 12'h  0;
rom[48646] = 12'h  0;
rom[48647] = 12'h  0;
rom[48648] = 12'h  0;
rom[48649] = 12'h  0;
rom[48650] = 12'h  0;
rom[48651] = 12'h  0;
rom[48652] = 12'h  0;
rom[48653] = 12'h  0;
rom[48654] = 12'h  0;
rom[48655] = 12'h  0;
rom[48656] = 12'h  0;
rom[48657] = 12'h  0;
rom[48658] = 12'h  0;
rom[48659] = 12'h  0;
rom[48660] = 12'h  0;
rom[48661] = 12'h  0;
rom[48662] = 12'h  0;
rom[48663] = 12'h  0;
rom[48664] = 12'h  0;
rom[48665] = 12'h  0;
rom[48666] = 12'h  0;
rom[48667] = 12'h  0;
rom[48668] = 12'h111;
rom[48669] = 12'h111;
rom[48670] = 12'h111;
rom[48671] = 12'h111;
rom[48672] = 12'h222;
rom[48673] = 12'h222;
rom[48674] = 12'h222;
rom[48675] = 12'h222;
rom[48676] = 12'h333;
rom[48677] = 12'h555;
rom[48678] = 12'h555;
rom[48679] = 12'h444;
rom[48680] = 12'h444;
rom[48681] = 12'h444;
rom[48682] = 12'h444;
rom[48683] = 12'h555;
rom[48684] = 12'h555;
rom[48685] = 12'h555;
rom[48686] = 12'h666;
rom[48687] = 12'h666;
rom[48688] = 12'h777;
rom[48689] = 12'h888;
rom[48690] = 12'h999;
rom[48691] = 12'h888;
rom[48692] = 12'h888;
rom[48693] = 12'h888;
rom[48694] = 12'h899;
rom[48695] = 12'h999;
rom[48696] = 12'h888;
rom[48697] = 12'h666;
rom[48698] = 12'h444;
rom[48699] = 12'h433;
rom[48700] = 12'h322;
rom[48701] = 12'h211;
rom[48702] = 12'h100;
rom[48703] = 12'h100;
rom[48704] = 12'h100;
rom[48705] = 12'h100;
rom[48706] = 12'h100;
rom[48707] = 12'h100;
rom[48708] = 12'h100;
rom[48709] = 12'h100;
rom[48710] = 12'h100;
rom[48711] = 12'h100;
rom[48712] = 12'h100;
rom[48713] = 12'h100;
rom[48714] = 12'h100;
rom[48715] = 12'h100;
rom[48716] = 12'h100;
rom[48717] = 12'h100;
rom[48718] = 12'h200;
rom[48719] = 12'h200;
rom[48720] = 12'h200;
rom[48721] = 12'h200;
rom[48722] = 12'h200;
rom[48723] = 12'h200;
rom[48724] = 12'h200;
rom[48725] = 12'h200;
rom[48726] = 12'h200;
rom[48727] = 12'h200;
rom[48728] = 12'h200;
rom[48729] = 12'h200;
rom[48730] = 12'h200;
rom[48731] = 12'h200;
rom[48732] = 12'h200;
rom[48733] = 12'h200;
rom[48734] = 12'h200;
rom[48735] = 12'h200;
rom[48736] = 12'h200;
rom[48737] = 12'h200;
rom[48738] = 12'h200;
rom[48739] = 12'h200;
rom[48740] = 12'h200;
rom[48741] = 12'h200;
rom[48742] = 12'h210;
rom[48743] = 12'h310;
rom[48744] = 12'h321;
rom[48745] = 12'h321;
rom[48746] = 12'h422;
rom[48747] = 12'h432;
rom[48748] = 12'h532;
rom[48749] = 12'h533;
rom[48750] = 12'h543;
rom[48751] = 12'h544;
rom[48752] = 12'h544;
rom[48753] = 12'h544;
rom[48754] = 12'h554;
rom[48755] = 12'h554;
rom[48756] = 12'h555;
rom[48757] = 12'h555;
rom[48758] = 12'h555;
rom[48759] = 12'h555;
rom[48760] = 12'h556;
rom[48761] = 12'h666;
rom[48762] = 12'h666;
rom[48763] = 12'h667;
rom[48764] = 12'h777;
rom[48765] = 12'h777;
rom[48766] = 12'h777;
rom[48767] = 12'h778;
rom[48768] = 12'h888;
rom[48769] = 12'h888;
rom[48770] = 12'h989;
rom[48771] = 12'h999;
rom[48772] = 12'ha9a;
rom[48773] = 12'haaa;
rom[48774] = 12'hbbb;
rom[48775] = 12'hcbb;
rom[48776] = 12'hccc;
rom[48777] = 12'hddd;
rom[48778] = 12'hddd;
rom[48779] = 12'hddd;
rom[48780] = 12'hccc;
rom[48781] = 12'hccc;
rom[48782] = 12'hcbb;
rom[48783] = 12'hcbb;
rom[48784] = 12'hbbb;
rom[48785] = 12'hbbb;
rom[48786] = 12'hbbb;
rom[48787] = 12'hbbb;
rom[48788] = 12'haaa;
rom[48789] = 12'haaa;
rom[48790] = 12'haaa;
rom[48791] = 12'haaa;
rom[48792] = 12'haaa;
rom[48793] = 12'haaa;
rom[48794] = 12'haaa;
rom[48795] = 12'haaa;
rom[48796] = 12'haaa;
rom[48797] = 12'haaa;
rom[48798] = 12'hbbb;
rom[48799] = 12'hbbb;
rom[48800] = 12'haaa;
rom[48801] = 12'haaa;
rom[48802] = 12'h999;
rom[48803] = 12'h999;
rom[48804] = 12'h999;
rom[48805] = 12'h888;
rom[48806] = 12'h888;
rom[48807] = 12'h888;
rom[48808] = 12'h777;
rom[48809] = 12'h777;
rom[48810] = 12'h777;
rom[48811] = 12'h777;
rom[48812] = 12'h777;
rom[48813] = 12'h777;
rom[48814] = 12'h777;
rom[48815] = 12'h777;
rom[48816] = 12'h777;
rom[48817] = 12'h777;
rom[48818] = 12'h777;
rom[48819] = 12'h777;
rom[48820] = 12'h777;
rom[48821] = 12'h777;
rom[48822] = 12'h777;
rom[48823] = 12'h777;
rom[48824] = 12'h777;
rom[48825] = 12'h777;
rom[48826] = 12'h777;
rom[48827] = 12'h777;
rom[48828] = 12'h888;
rom[48829] = 12'h888;
rom[48830] = 12'h888;
rom[48831] = 12'h888;
rom[48832] = 12'h888;
rom[48833] = 12'h777;
rom[48834] = 12'h777;
rom[48835] = 12'h777;
rom[48836] = 12'h777;
rom[48837] = 12'h777;
rom[48838] = 12'h888;
rom[48839] = 12'h888;
rom[48840] = 12'h777;
rom[48841] = 12'h777;
rom[48842] = 12'h777;
rom[48843] = 12'h777;
rom[48844] = 12'h777;
rom[48845] = 12'h777;
rom[48846] = 12'h777;
rom[48847] = 12'h888;
rom[48848] = 12'h888;
rom[48849] = 12'h888;
rom[48850] = 12'h888;
rom[48851] = 12'h888;
rom[48852] = 12'h888;
rom[48853] = 12'h888;
rom[48854] = 12'h888;
rom[48855] = 12'h888;
rom[48856] = 12'h999;
rom[48857] = 12'h999;
rom[48858] = 12'h999;
rom[48859] = 12'h999;
rom[48860] = 12'h999;
rom[48861] = 12'h999;
rom[48862] = 12'h999;
rom[48863] = 12'h999;
rom[48864] = 12'haaa;
rom[48865] = 12'haaa;
rom[48866] = 12'haaa;
rom[48867] = 12'haaa;
rom[48868] = 12'haaa;
rom[48869] = 12'haaa;
rom[48870] = 12'haaa;
rom[48871] = 12'haaa;
rom[48872] = 12'h999;
rom[48873] = 12'h999;
rom[48874] = 12'h999;
rom[48875] = 12'h999;
rom[48876] = 12'h999;
rom[48877] = 12'h999;
rom[48878] = 12'h888;
rom[48879] = 12'h888;
rom[48880] = 12'h777;
rom[48881] = 12'h777;
rom[48882] = 12'h777;
rom[48883] = 12'h777;
rom[48884] = 12'h777;
rom[48885] = 12'h666;
rom[48886] = 12'h666;
rom[48887] = 12'h666;
rom[48888] = 12'h666;
rom[48889] = 12'h666;
rom[48890] = 12'h666;
rom[48891] = 12'h666;
rom[48892] = 12'h666;
rom[48893] = 12'h666;
rom[48894] = 12'h666;
rom[48895] = 12'h666;
rom[48896] = 12'h666;
rom[48897] = 12'h666;
rom[48898] = 12'h666;
rom[48899] = 12'h666;
rom[48900] = 12'h666;
rom[48901] = 12'h666;
rom[48902] = 12'h555;
rom[48903] = 12'h555;
rom[48904] = 12'h444;
rom[48905] = 12'h444;
rom[48906] = 12'h444;
rom[48907] = 12'h444;
rom[48908] = 12'h444;
rom[48909] = 12'h555;
rom[48910] = 12'h444;
rom[48911] = 12'h444;
rom[48912] = 12'h444;
rom[48913] = 12'h333;
rom[48914] = 12'h333;
rom[48915] = 12'h222;
rom[48916] = 12'h222;
rom[48917] = 12'h222;
rom[48918] = 12'h222;
rom[48919] = 12'h111;
rom[48920] = 12'h111;
rom[48921] = 12'h111;
rom[48922] = 12'h  0;
rom[48923] = 12'h  0;
rom[48924] = 12'h  0;
rom[48925] = 12'h  0;
rom[48926] = 12'h  0;
rom[48927] = 12'h  0;
rom[48928] = 12'h  0;
rom[48929] = 12'h  0;
rom[48930] = 12'h  0;
rom[48931] = 12'h  0;
rom[48932] = 12'h  0;
rom[48933] = 12'h  0;
rom[48934] = 12'h  0;
rom[48935] = 12'h  0;
rom[48936] = 12'h  0;
rom[48937] = 12'h  0;
rom[48938] = 12'h  0;
rom[48939] = 12'h  0;
rom[48940] = 12'h  0;
rom[48941] = 12'h  0;
rom[48942] = 12'h  0;
rom[48943] = 12'h  0;
rom[48944] = 12'h  0;
rom[48945] = 12'h  0;
rom[48946] = 12'h  0;
rom[48947] = 12'h  0;
rom[48948] = 12'h  0;
rom[48949] = 12'h  0;
rom[48950] = 12'h  0;
rom[48951] = 12'h111;
rom[48952] = 12'h111;
rom[48953] = 12'h111;
rom[48954] = 12'h111;
rom[48955] = 12'h111;
rom[48956] = 12'h111;
rom[48957] = 12'h111;
rom[48958] = 12'h111;
rom[48959] = 12'h111;
rom[48960] = 12'h111;
rom[48961] = 12'h111;
rom[48962] = 12'h111;
rom[48963] = 12'h111;
rom[48964] = 12'h111;
rom[48965] = 12'h111;
rom[48966] = 12'h111;
rom[48967] = 12'h111;
rom[48968] = 12'h111;
rom[48969] = 12'h111;
rom[48970] = 12'h111;
rom[48971] = 12'h111;
rom[48972] = 12'h111;
rom[48973] = 12'h111;
rom[48974] = 12'h111;
rom[48975] = 12'h111;
rom[48976] = 12'h111;
rom[48977] = 12'h111;
rom[48978] = 12'h111;
rom[48979] = 12'h111;
rom[48980] = 12'h111;
rom[48981] = 12'h111;
rom[48982] = 12'h111;
rom[48983] = 12'h111;
rom[48984] = 12'h111;
rom[48985] = 12'h111;
rom[48986] = 12'h111;
rom[48987] = 12'h111;
rom[48988] = 12'h111;
rom[48989] = 12'h111;
rom[48990] = 12'h111;
rom[48991] = 12'h  0;
rom[48992] = 12'h  0;
rom[48993] = 12'h  0;
rom[48994] = 12'h  0;
rom[48995] = 12'h  0;
rom[48996] = 12'h  0;
rom[48997] = 12'h  0;
rom[48998] = 12'h  0;
rom[48999] = 12'h  0;
rom[49000] = 12'h  0;
rom[49001] = 12'h  0;
rom[49002] = 12'h  0;
rom[49003] = 12'h  0;
rom[49004] = 12'h  0;
rom[49005] = 12'h  0;
rom[49006] = 12'h  0;
rom[49007] = 12'h  0;
rom[49008] = 12'h111;
rom[49009] = 12'h111;
rom[49010] = 12'h111;
rom[49011] = 12'h111;
rom[49012] = 12'h111;
rom[49013] = 12'h111;
rom[49014] = 12'h111;
rom[49015] = 12'h111;
rom[49016] = 12'h111;
rom[49017] = 12'h111;
rom[49018] = 12'h111;
rom[49019] = 12'h222;
rom[49020] = 12'h222;
rom[49021] = 12'h222;
rom[49022] = 12'h222;
rom[49023] = 12'h222;
rom[49024] = 12'h222;
rom[49025] = 12'h222;
rom[49026] = 12'h222;
rom[49027] = 12'h222;
rom[49028] = 12'h222;
rom[49029] = 12'h222;
rom[49030] = 12'h111;
rom[49031] = 12'h111;
rom[49032] = 12'h111;
rom[49033] = 12'h111;
rom[49034] = 12'h111;
rom[49035] = 12'h111;
rom[49036] = 12'h  0;
rom[49037] = 12'h  0;
rom[49038] = 12'h  0;
rom[49039] = 12'h  0;
rom[49040] = 12'h  0;
rom[49041] = 12'h  0;
rom[49042] = 12'h  0;
rom[49043] = 12'h  0;
rom[49044] = 12'h  0;
rom[49045] = 12'h  0;
rom[49046] = 12'h  0;
rom[49047] = 12'h  0;
rom[49048] = 12'h  0;
rom[49049] = 12'h  0;
rom[49050] = 12'h  0;
rom[49051] = 12'h  0;
rom[49052] = 12'h  0;
rom[49053] = 12'h  0;
rom[49054] = 12'h  0;
rom[49055] = 12'h  0;
rom[49056] = 12'h  0;
rom[49057] = 12'h  0;
rom[49058] = 12'h  0;
rom[49059] = 12'h  0;
rom[49060] = 12'h  0;
rom[49061] = 12'h  0;
rom[49062] = 12'h  0;
rom[49063] = 12'h  0;
rom[49064] = 12'h  0;
rom[49065] = 12'h  0;
rom[49066] = 12'h  0;
rom[49067] = 12'h  0;
rom[49068] = 12'h111;
rom[49069] = 12'h111;
rom[49070] = 12'h111;
rom[49071] = 12'h111;
rom[49072] = 12'h222;
rom[49073] = 12'h222;
rom[49074] = 12'h222;
rom[49075] = 12'h222;
rom[49076] = 12'h444;
rom[49077] = 12'h555;
rom[49078] = 12'h555;
rom[49079] = 12'h444;
rom[49080] = 12'h444;
rom[49081] = 12'h444;
rom[49082] = 12'h444;
rom[49083] = 12'h555;
rom[49084] = 12'h555;
rom[49085] = 12'h555;
rom[49086] = 12'h666;
rom[49087] = 12'h666;
rom[49088] = 12'h777;
rom[49089] = 12'h888;
rom[49090] = 12'h888;
rom[49091] = 12'h888;
rom[49092] = 12'h777;
rom[49093] = 12'h777;
rom[49094] = 12'h888;
rom[49095] = 12'h999;
rom[49096] = 12'h888;
rom[49097] = 12'h777;
rom[49098] = 12'h555;
rom[49099] = 12'h444;
rom[49100] = 12'h333;
rom[49101] = 12'h222;
rom[49102] = 12'h111;
rom[49103] = 12'h100;
rom[49104] = 12'h100;
rom[49105] = 12'h100;
rom[49106] = 12'h100;
rom[49107] = 12'h100;
rom[49108] = 12'h100;
rom[49109] = 12'h100;
rom[49110] = 12'h100;
rom[49111] = 12'h100;
rom[49112] = 12'h100;
rom[49113] = 12'h100;
rom[49114] = 12'h100;
rom[49115] = 12'h100;
rom[49116] = 12'h200;
rom[49117] = 12'h200;
rom[49118] = 12'h200;
rom[49119] = 12'h200;
rom[49120] = 12'h200;
rom[49121] = 12'h200;
rom[49122] = 12'h200;
rom[49123] = 12'h200;
rom[49124] = 12'h200;
rom[49125] = 12'h200;
rom[49126] = 12'h200;
rom[49127] = 12'h200;
rom[49128] = 12'h200;
rom[49129] = 12'h200;
rom[49130] = 12'h200;
rom[49131] = 12'h200;
rom[49132] = 12'h200;
rom[49133] = 12'h200;
rom[49134] = 12'h200;
rom[49135] = 12'h200;
rom[49136] = 12'h200;
rom[49137] = 12'h200;
rom[49138] = 12'h100;
rom[49139] = 12'h100;
rom[49140] = 12'h100;
rom[49141] = 12'h200;
rom[49142] = 12'h211;
rom[49143] = 12'h321;
rom[49144] = 12'h422;
rom[49145] = 12'h432;
rom[49146] = 12'h433;
rom[49147] = 12'h543;
rom[49148] = 12'h543;
rom[49149] = 12'h543;
rom[49150] = 12'h544;
rom[49151] = 12'h544;
rom[49152] = 12'h544;
rom[49153] = 12'h554;
rom[49154] = 12'h555;
rom[49155] = 12'h555;
rom[49156] = 12'h555;
rom[49157] = 12'h555;
rom[49158] = 12'h555;
rom[49159] = 12'h566;
rom[49160] = 12'h666;
rom[49161] = 12'h666;
rom[49162] = 12'h677;
rom[49163] = 12'h777;
rom[49164] = 12'h777;
rom[49165] = 12'h777;
rom[49166] = 12'h888;
rom[49167] = 12'h888;
rom[49168] = 12'h888;
rom[49169] = 12'h889;
rom[49170] = 12'h999;
rom[49171] = 12'haaa;
rom[49172] = 12'haaa;
rom[49173] = 12'hbab;
rom[49174] = 12'hbbb;
rom[49175] = 12'hccc;
rom[49176] = 12'hddd;
rom[49177] = 12'hddd;
rom[49178] = 12'hddd;
rom[49179] = 12'hcdc;
rom[49180] = 12'hccc;
rom[49181] = 12'hccb;
rom[49182] = 12'hbcb;
rom[49183] = 12'hbbb;
rom[49184] = 12'hbbb;
rom[49185] = 12'hbbb;
rom[49186] = 12'hbbb;
rom[49187] = 12'hbbb;
rom[49188] = 12'hbbb;
rom[49189] = 12'hbbb;
rom[49190] = 12'hbbb;
rom[49191] = 12'hbbb;
rom[49192] = 12'hbbb;
rom[49193] = 12'haaa;
rom[49194] = 12'haaa;
rom[49195] = 12'haaa;
rom[49196] = 12'haaa;
rom[49197] = 12'haaa;
rom[49198] = 12'haaa;
rom[49199] = 12'hbbb;
rom[49200] = 12'haaa;
rom[49201] = 12'haaa;
rom[49202] = 12'h999;
rom[49203] = 12'h999;
rom[49204] = 12'h999;
rom[49205] = 12'h999;
rom[49206] = 12'h888;
rom[49207] = 12'h888;
rom[49208] = 12'h777;
rom[49209] = 12'h777;
rom[49210] = 12'h777;
rom[49211] = 12'h777;
rom[49212] = 12'h777;
rom[49213] = 12'h777;
rom[49214] = 12'h777;
rom[49215] = 12'h777;
rom[49216] = 12'h777;
rom[49217] = 12'h777;
rom[49218] = 12'h777;
rom[49219] = 12'h777;
rom[49220] = 12'h777;
rom[49221] = 12'h777;
rom[49222] = 12'h777;
rom[49223] = 12'h777;
rom[49224] = 12'h777;
rom[49225] = 12'h777;
rom[49226] = 12'h888;
rom[49227] = 12'h888;
rom[49228] = 12'h888;
rom[49229] = 12'h888;
rom[49230] = 12'h888;
rom[49231] = 12'h888;
rom[49232] = 12'h888;
rom[49233] = 12'h777;
rom[49234] = 12'h777;
rom[49235] = 12'h777;
rom[49236] = 12'h777;
rom[49237] = 12'h888;
rom[49238] = 12'h888;
rom[49239] = 12'h888;
rom[49240] = 12'h888;
rom[49241] = 12'h888;
rom[49242] = 12'h777;
rom[49243] = 12'h777;
rom[49244] = 12'h777;
rom[49245] = 12'h777;
rom[49246] = 12'h888;
rom[49247] = 12'h888;
rom[49248] = 12'h888;
rom[49249] = 12'h888;
rom[49250] = 12'h888;
rom[49251] = 12'h888;
rom[49252] = 12'h888;
rom[49253] = 12'h888;
rom[49254] = 12'h888;
rom[49255] = 12'h888;
rom[49256] = 12'h999;
rom[49257] = 12'h999;
rom[49258] = 12'h999;
rom[49259] = 12'h999;
rom[49260] = 12'h999;
rom[49261] = 12'h999;
rom[49262] = 12'h999;
rom[49263] = 12'h999;
rom[49264] = 12'haaa;
rom[49265] = 12'haaa;
rom[49266] = 12'haaa;
rom[49267] = 12'haaa;
rom[49268] = 12'hbbb;
rom[49269] = 12'hbbb;
rom[49270] = 12'haaa;
rom[49271] = 12'haaa;
rom[49272] = 12'h999;
rom[49273] = 12'h999;
rom[49274] = 12'h999;
rom[49275] = 12'h999;
rom[49276] = 12'h999;
rom[49277] = 12'h999;
rom[49278] = 12'h888;
rom[49279] = 12'h888;
rom[49280] = 12'h888;
rom[49281] = 12'h888;
rom[49282] = 12'h888;
rom[49283] = 12'h888;
rom[49284] = 12'h777;
rom[49285] = 12'h777;
rom[49286] = 12'h777;
rom[49287] = 12'h666;
rom[49288] = 12'h666;
rom[49289] = 12'h666;
rom[49290] = 12'h666;
rom[49291] = 12'h666;
rom[49292] = 12'h666;
rom[49293] = 12'h666;
rom[49294] = 12'h666;
rom[49295] = 12'h666;
rom[49296] = 12'h666;
rom[49297] = 12'h666;
rom[49298] = 12'h666;
rom[49299] = 12'h666;
rom[49300] = 12'h666;
rom[49301] = 12'h666;
rom[49302] = 12'h666;
rom[49303] = 12'h666;
rom[49304] = 12'h555;
rom[49305] = 12'h444;
rom[49306] = 12'h444;
rom[49307] = 12'h444;
rom[49308] = 12'h444;
rom[49309] = 12'h444;
rom[49310] = 12'h444;
rom[49311] = 12'h444;
rom[49312] = 12'h444;
rom[49313] = 12'h444;
rom[49314] = 12'h333;
rom[49315] = 12'h333;
rom[49316] = 12'h333;
rom[49317] = 12'h222;
rom[49318] = 12'h222;
rom[49319] = 12'h111;
rom[49320] = 12'h111;
rom[49321] = 12'h111;
rom[49322] = 12'h  0;
rom[49323] = 12'h  0;
rom[49324] = 12'h  0;
rom[49325] = 12'h  0;
rom[49326] = 12'h  0;
rom[49327] = 12'h  0;
rom[49328] = 12'h  0;
rom[49329] = 12'h  0;
rom[49330] = 12'h  0;
rom[49331] = 12'h  0;
rom[49332] = 12'h  0;
rom[49333] = 12'h  0;
rom[49334] = 12'h  0;
rom[49335] = 12'h  0;
rom[49336] = 12'h  0;
rom[49337] = 12'h  0;
rom[49338] = 12'h  0;
rom[49339] = 12'h  0;
rom[49340] = 12'h  0;
rom[49341] = 12'h  0;
rom[49342] = 12'h  0;
rom[49343] = 12'h  0;
rom[49344] = 12'h  0;
rom[49345] = 12'h  0;
rom[49346] = 12'h  0;
rom[49347] = 12'h  0;
rom[49348] = 12'h  0;
rom[49349] = 12'h  0;
rom[49350] = 12'h  0;
rom[49351] = 12'h111;
rom[49352] = 12'h111;
rom[49353] = 12'h111;
rom[49354] = 12'h111;
rom[49355] = 12'h111;
rom[49356] = 12'h111;
rom[49357] = 12'h111;
rom[49358] = 12'h111;
rom[49359] = 12'h111;
rom[49360] = 12'h111;
rom[49361] = 12'h111;
rom[49362] = 12'h111;
rom[49363] = 12'h111;
rom[49364] = 12'h111;
rom[49365] = 12'h111;
rom[49366] = 12'h111;
rom[49367] = 12'h111;
rom[49368] = 12'h111;
rom[49369] = 12'h111;
rom[49370] = 12'h111;
rom[49371] = 12'h111;
rom[49372] = 12'h111;
rom[49373] = 12'h111;
rom[49374] = 12'h111;
rom[49375] = 12'h111;
rom[49376] = 12'h111;
rom[49377] = 12'h111;
rom[49378] = 12'h111;
rom[49379] = 12'h111;
rom[49380] = 12'h111;
rom[49381] = 12'h111;
rom[49382] = 12'h111;
rom[49383] = 12'h111;
rom[49384] = 12'h111;
rom[49385] = 12'h111;
rom[49386] = 12'h111;
rom[49387] = 12'h111;
rom[49388] = 12'h111;
rom[49389] = 12'h  0;
rom[49390] = 12'h  0;
rom[49391] = 12'h  0;
rom[49392] = 12'h  0;
rom[49393] = 12'h  0;
rom[49394] = 12'h  0;
rom[49395] = 12'h  0;
rom[49396] = 12'h  0;
rom[49397] = 12'h  0;
rom[49398] = 12'h  0;
rom[49399] = 12'h  0;
rom[49400] = 12'h  0;
rom[49401] = 12'h  0;
rom[49402] = 12'h  0;
rom[49403] = 12'h  0;
rom[49404] = 12'h  0;
rom[49405] = 12'h  0;
rom[49406] = 12'h  0;
rom[49407] = 12'h  0;
rom[49408] = 12'h111;
rom[49409] = 12'h111;
rom[49410] = 12'h111;
rom[49411] = 12'h111;
rom[49412] = 12'h111;
rom[49413] = 12'h111;
rom[49414] = 12'h111;
rom[49415] = 12'h111;
rom[49416] = 12'h111;
rom[49417] = 12'h111;
rom[49418] = 12'h111;
rom[49419] = 12'h111;
rom[49420] = 12'h111;
rom[49421] = 12'h222;
rom[49422] = 12'h222;
rom[49423] = 12'h222;
rom[49424] = 12'h222;
rom[49425] = 12'h222;
rom[49426] = 12'h222;
rom[49427] = 12'h222;
rom[49428] = 12'h222;
rom[49429] = 12'h222;
rom[49430] = 12'h111;
rom[49431] = 12'h111;
rom[49432] = 12'h111;
rom[49433] = 12'h111;
rom[49434] = 12'h111;
rom[49435] = 12'h111;
rom[49436] = 12'h  0;
rom[49437] = 12'h  0;
rom[49438] = 12'h  0;
rom[49439] = 12'h  0;
rom[49440] = 12'h  0;
rom[49441] = 12'h  0;
rom[49442] = 12'h  0;
rom[49443] = 12'h  0;
rom[49444] = 12'h  0;
rom[49445] = 12'h  0;
rom[49446] = 12'h  0;
rom[49447] = 12'h  0;
rom[49448] = 12'h  0;
rom[49449] = 12'h  0;
rom[49450] = 12'h  0;
rom[49451] = 12'h  0;
rom[49452] = 12'h  0;
rom[49453] = 12'h  0;
rom[49454] = 12'h  0;
rom[49455] = 12'h  0;
rom[49456] = 12'h  0;
rom[49457] = 12'h  0;
rom[49458] = 12'h  0;
rom[49459] = 12'h  0;
rom[49460] = 12'h  0;
rom[49461] = 12'h  0;
rom[49462] = 12'h  0;
rom[49463] = 12'h  0;
rom[49464] = 12'h  0;
rom[49465] = 12'h  0;
rom[49466] = 12'h  0;
rom[49467] = 12'h  0;
rom[49468] = 12'h  0;
rom[49469] = 12'h111;
rom[49470] = 12'h111;
rom[49471] = 12'h111;
rom[49472] = 12'h111;
rom[49473] = 12'h222;
rom[49474] = 12'h222;
rom[49475] = 12'h333;
rom[49476] = 12'h444;
rom[49477] = 12'h555;
rom[49478] = 12'h444;
rom[49479] = 12'h444;
rom[49480] = 12'h333;
rom[49481] = 12'h444;
rom[49482] = 12'h444;
rom[49483] = 12'h555;
rom[49484] = 12'h555;
rom[49485] = 12'h555;
rom[49486] = 12'h666;
rom[49487] = 12'h666;
rom[49488] = 12'h777;
rom[49489] = 12'h888;
rom[49490] = 12'h888;
rom[49491] = 12'h777;
rom[49492] = 12'h777;
rom[49493] = 12'h777;
rom[49494] = 12'h888;
rom[49495] = 12'h899;
rom[49496] = 12'h888;
rom[49497] = 12'h777;
rom[49498] = 12'h565;
rom[49499] = 12'h454;
rom[49500] = 12'h433;
rom[49501] = 12'h322;
rom[49502] = 12'h211;
rom[49503] = 12'h111;
rom[49504] = 12'h100;
rom[49505] = 12'h100;
rom[49506] = 12'h100;
rom[49507] = 12'h100;
rom[49508] = 12'h100;
rom[49509] = 12'h100;
rom[49510] = 12'h100;
rom[49511] = 12'h100;
rom[49512] = 12'h100;
rom[49513] = 12'h100;
rom[49514] = 12'h100;
rom[49515] = 12'h100;
rom[49516] = 12'h100;
rom[49517] = 12'h100;
rom[49518] = 12'h200;
rom[49519] = 12'h200;
rom[49520] = 12'h200;
rom[49521] = 12'h200;
rom[49522] = 12'h200;
rom[49523] = 12'h200;
rom[49524] = 12'h200;
rom[49525] = 12'h200;
rom[49526] = 12'h200;
rom[49527] = 12'h100;
rom[49528] = 12'h200;
rom[49529] = 12'h100;
rom[49530] = 12'h200;
rom[49531] = 12'h100;
rom[49532] = 12'h100;
rom[49533] = 12'h200;
rom[49534] = 12'h200;
rom[49535] = 12'h100;
rom[49536] = 12'h100;
rom[49537] = 12'h100;
rom[49538] = 12'h200;
rom[49539] = 12'h200;
rom[49540] = 12'h211;
rom[49541] = 12'h211;
rom[49542] = 12'h322;
rom[49543] = 12'h332;
rom[49544] = 12'h433;
rom[49545] = 12'h443;
rom[49546] = 12'h543;
rom[49547] = 12'h544;
rom[49548] = 12'h544;
rom[49549] = 12'h544;
rom[49550] = 12'h544;
rom[49551] = 12'h544;
rom[49552] = 12'h554;
rom[49553] = 12'h555;
rom[49554] = 12'h555;
rom[49555] = 12'h555;
rom[49556] = 12'h555;
rom[49557] = 12'h555;
rom[49558] = 12'h566;
rom[49559] = 12'h666;
rom[49560] = 12'h666;
rom[49561] = 12'h677;
rom[49562] = 12'h777;
rom[49563] = 12'h777;
rom[49564] = 12'h777;
rom[49565] = 12'h778;
rom[49566] = 12'h888;
rom[49567] = 12'h888;
rom[49568] = 12'h889;
rom[49569] = 12'h999;
rom[49570] = 12'h99a;
rom[49571] = 12'haaa;
rom[49572] = 12'hbbb;
rom[49573] = 12'hbbb;
rom[49574] = 12'hccc;
rom[49575] = 12'hccc;
rom[49576] = 12'hddd;
rom[49577] = 12'hddd;
rom[49578] = 12'hddc;
rom[49579] = 12'hccc;
rom[49580] = 12'hccc;
rom[49581] = 12'hccb;
rom[49582] = 12'hbbb;
rom[49583] = 12'hbbb;
rom[49584] = 12'hbbb;
rom[49585] = 12'hbbb;
rom[49586] = 12'hbbb;
rom[49587] = 12'hbbb;
rom[49588] = 12'hbbb;
rom[49589] = 12'hbbb;
rom[49590] = 12'hbbb;
rom[49591] = 12'hbbb;
rom[49592] = 12'hbbb;
rom[49593] = 12'hbbb;
rom[49594] = 12'hbbb;
rom[49595] = 12'haaa;
rom[49596] = 12'haaa;
rom[49597] = 12'haaa;
rom[49598] = 12'haaa;
rom[49599] = 12'hbbb;
rom[49600] = 12'haaa;
rom[49601] = 12'haaa;
rom[49602] = 12'haaa;
rom[49603] = 12'h999;
rom[49604] = 12'h999;
rom[49605] = 12'h999;
rom[49606] = 12'h888;
rom[49607] = 12'h888;
rom[49608] = 12'h888;
rom[49609] = 12'h888;
rom[49610] = 12'h777;
rom[49611] = 12'h777;
rom[49612] = 12'h777;
rom[49613] = 12'h777;
rom[49614] = 12'h777;
rom[49615] = 12'h777;
rom[49616] = 12'h777;
rom[49617] = 12'h777;
rom[49618] = 12'h777;
rom[49619] = 12'h777;
rom[49620] = 12'h777;
rom[49621] = 12'h777;
rom[49622] = 12'h777;
rom[49623] = 12'h777;
rom[49624] = 12'h888;
rom[49625] = 12'h888;
rom[49626] = 12'h888;
rom[49627] = 12'h888;
rom[49628] = 12'h888;
rom[49629] = 12'h888;
rom[49630] = 12'h888;
rom[49631] = 12'h888;
rom[49632] = 12'h888;
rom[49633] = 12'h888;
rom[49634] = 12'h777;
rom[49635] = 12'h777;
rom[49636] = 12'h888;
rom[49637] = 12'h888;
rom[49638] = 12'h888;
rom[49639] = 12'h888;
rom[49640] = 12'h888;
rom[49641] = 12'h888;
rom[49642] = 12'h888;
rom[49643] = 12'h888;
rom[49644] = 12'h888;
rom[49645] = 12'h888;
rom[49646] = 12'h888;
rom[49647] = 12'h888;
rom[49648] = 12'h888;
rom[49649] = 12'h888;
rom[49650] = 12'h888;
rom[49651] = 12'h888;
rom[49652] = 12'h888;
rom[49653] = 12'h888;
rom[49654] = 12'h999;
rom[49655] = 12'h999;
rom[49656] = 12'h999;
rom[49657] = 12'h999;
rom[49658] = 12'h999;
rom[49659] = 12'h999;
rom[49660] = 12'h999;
rom[49661] = 12'h999;
rom[49662] = 12'h999;
rom[49663] = 12'haaa;
rom[49664] = 12'haaa;
rom[49665] = 12'haaa;
rom[49666] = 12'haaa;
rom[49667] = 12'haaa;
rom[49668] = 12'hbbb;
rom[49669] = 12'hbbb;
rom[49670] = 12'hbbb;
rom[49671] = 12'haaa;
rom[49672] = 12'haaa;
rom[49673] = 12'h999;
rom[49674] = 12'h999;
rom[49675] = 12'h888;
rom[49676] = 12'h888;
rom[49677] = 12'h888;
rom[49678] = 12'h888;
rom[49679] = 12'h888;
rom[49680] = 12'h888;
rom[49681] = 12'h888;
rom[49682] = 12'h888;
rom[49683] = 12'h888;
rom[49684] = 12'h888;
rom[49685] = 12'h888;
rom[49686] = 12'h888;
rom[49687] = 12'h777;
rom[49688] = 12'h777;
rom[49689] = 12'h777;
rom[49690] = 12'h666;
rom[49691] = 12'h666;
rom[49692] = 12'h666;
rom[49693] = 12'h666;
rom[49694] = 12'h666;
rom[49695] = 12'h666;
rom[49696] = 12'h666;
rom[49697] = 12'h666;
rom[49698] = 12'h666;
rom[49699] = 12'h666;
rom[49700] = 12'h666;
rom[49701] = 12'h666;
rom[49702] = 12'h666;
rom[49703] = 12'h666;
rom[49704] = 12'h555;
rom[49705] = 12'h555;
rom[49706] = 12'h555;
rom[49707] = 12'h444;
rom[49708] = 12'h444;
rom[49709] = 12'h444;
rom[49710] = 12'h444;
rom[49711] = 12'h444;
rom[49712] = 12'h444;
rom[49713] = 12'h444;
rom[49714] = 12'h444;
rom[49715] = 12'h333;
rom[49716] = 12'h333;
rom[49717] = 12'h222;
rom[49718] = 12'h222;
rom[49719] = 12'h111;
rom[49720] = 12'h111;
rom[49721] = 12'h111;
rom[49722] = 12'h111;
rom[49723] = 12'h111;
rom[49724] = 12'h  0;
rom[49725] = 12'h  0;
rom[49726] = 12'h  0;
rom[49727] = 12'h  0;
rom[49728] = 12'h  0;
rom[49729] = 12'h  0;
rom[49730] = 12'h  0;
rom[49731] = 12'h  0;
rom[49732] = 12'h  0;
rom[49733] = 12'h  0;
rom[49734] = 12'h  0;
rom[49735] = 12'h  0;
rom[49736] = 12'h  0;
rom[49737] = 12'h  0;
rom[49738] = 12'h  0;
rom[49739] = 12'h  0;
rom[49740] = 12'h  0;
rom[49741] = 12'h  0;
rom[49742] = 12'h  0;
rom[49743] = 12'h  0;
rom[49744] = 12'h  0;
rom[49745] = 12'h  0;
rom[49746] = 12'h  0;
rom[49747] = 12'h  0;
rom[49748] = 12'h  0;
rom[49749] = 12'h111;
rom[49750] = 12'h111;
rom[49751] = 12'h111;
rom[49752] = 12'h111;
rom[49753] = 12'h111;
rom[49754] = 12'h111;
rom[49755] = 12'h111;
rom[49756] = 12'h111;
rom[49757] = 12'h111;
rom[49758] = 12'h111;
rom[49759] = 12'h111;
rom[49760] = 12'h111;
rom[49761] = 12'h111;
rom[49762] = 12'h111;
rom[49763] = 12'h111;
rom[49764] = 12'h111;
rom[49765] = 12'h111;
rom[49766] = 12'h111;
rom[49767] = 12'h111;
rom[49768] = 12'h111;
rom[49769] = 12'h111;
rom[49770] = 12'h111;
rom[49771] = 12'h111;
rom[49772] = 12'h111;
rom[49773] = 12'h111;
rom[49774] = 12'h111;
rom[49775] = 12'h111;
rom[49776] = 12'h111;
rom[49777] = 12'h111;
rom[49778] = 12'h111;
rom[49779] = 12'h111;
rom[49780] = 12'h111;
rom[49781] = 12'h111;
rom[49782] = 12'h111;
rom[49783] = 12'h111;
rom[49784] = 12'h111;
rom[49785] = 12'h111;
rom[49786] = 12'h111;
rom[49787] = 12'h  0;
rom[49788] = 12'h  0;
rom[49789] = 12'h  0;
rom[49790] = 12'h  0;
rom[49791] = 12'h  0;
rom[49792] = 12'h  0;
rom[49793] = 12'h  0;
rom[49794] = 12'h  0;
rom[49795] = 12'h  0;
rom[49796] = 12'h  0;
rom[49797] = 12'h  0;
rom[49798] = 12'h  0;
rom[49799] = 12'h  0;
rom[49800] = 12'h  0;
rom[49801] = 12'h  0;
rom[49802] = 12'h  0;
rom[49803] = 12'h  0;
rom[49804] = 12'h  0;
rom[49805] = 12'h  0;
rom[49806] = 12'h  0;
rom[49807] = 12'h  0;
rom[49808] = 12'h111;
rom[49809] = 12'h111;
rom[49810] = 12'h111;
rom[49811] = 12'h111;
rom[49812] = 12'h111;
rom[49813] = 12'h111;
rom[49814] = 12'h111;
rom[49815] = 12'h111;
rom[49816] = 12'h111;
rom[49817] = 12'h111;
rom[49818] = 12'h111;
rom[49819] = 12'h111;
rom[49820] = 12'h111;
rom[49821] = 12'h222;
rom[49822] = 12'h222;
rom[49823] = 12'h222;
rom[49824] = 12'h222;
rom[49825] = 12'h222;
rom[49826] = 12'h222;
rom[49827] = 12'h222;
rom[49828] = 12'h222;
rom[49829] = 12'h111;
rom[49830] = 12'h111;
rom[49831] = 12'h111;
rom[49832] = 12'h111;
rom[49833] = 12'h111;
rom[49834] = 12'h111;
rom[49835] = 12'h  0;
rom[49836] = 12'h  0;
rom[49837] = 12'h  0;
rom[49838] = 12'h  0;
rom[49839] = 12'h  0;
rom[49840] = 12'h  0;
rom[49841] = 12'h  0;
rom[49842] = 12'h  0;
rom[49843] = 12'h  0;
rom[49844] = 12'h  0;
rom[49845] = 12'h  0;
rom[49846] = 12'h  0;
rom[49847] = 12'h  0;
rom[49848] = 12'h  0;
rom[49849] = 12'h  0;
rom[49850] = 12'h  0;
rom[49851] = 12'h  0;
rom[49852] = 12'h  0;
rom[49853] = 12'h  0;
rom[49854] = 12'h  0;
rom[49855] = 12'h  0;
rom[49856] = 12'h  0;
rom[49857] = 12'h  0;
rom[49858] = 12'h  0;
rom[49859] = 12'h  0;
rom[49860] = 12'h  0;
rom[49861] = 12'h  0;
rom[49862] = 12'h  0;
rom[49863] = 12'h  0;
rom[49864] = 12'h  0;
rom[49865] = 12'h  0;
rom[49866] = 12'h  0;
rom[49867] = 12'h  0;
rom[49868] = 12'h  0;
rom[49869] = 12'h111;
rom[49870] = 12'h111;
rom[49871] = 12'h111;
rom[49872] = 12'h111;
rom[49873] = 12'h222;
rom[49874] = 12'h222;
rom[49875] = 12'h333;
rom[49876] = 12'h444;
rom[49877] = 12'h555;
rom[49878] = 12'h444;
rom[49879] = 12'h444;
rom[49880] = 12'h333;
rom[49881] = 12'h444;
rom[49882] = 12'h444;
rom[49883] = 12'h555;
rom[49884] = 12'h555;
rom[49885] = 12'h555;
rom[49886] = 12'h666;
rom[49887] = 12'h666;
rom[49888] = 12'h777;
rom[49889] = 12'h888;
rom[49890] = 12'h887;
rom[49891] = 12'h777;
rom[49892] = 12'h666;
rom[49893] = 12'h777;
rom[49894] = 12'h788;
rom[49895] = 12'h888;
rom[49896] = 12'h888;
rom[49897] = 12'h777;
rom[49898] = 12'h666;
rom[49899] = 12'h555;
rom[49900] = 12'h444;
rom[49901] = 12'h333;
rom[49902] = 12'h222;
rom[49903] = 12'h211;
rom[49904] = 12'h110;
rom[49905] = 12'h100;
rom[49906] = 12'h100;
rom[49907] = 12'h  0;
rom[49908] = 12'h100;
rom[49909] = 12'h100;
rom[49910] = 12'h100;
rom[49911] = 12'h100;
rom[49912] = 12'h100;
rom[49913] = 12'h100;
rom[49914] = 12'h100;
rom[49915] = 12'h100;
rom[49916] = 12'h100;
rom[49917] = 12'h100;
rom[49918] = 12'h100;
rom[49919] = 12'h100;
rom[49920] = 12'h100;
rom[49921] = 12'h100;
rom[49922] = 12'h100;
rom[49923] = 12'h100;
rom[49924] = 12'h100;
rom[49925] = 12'h100;
rom[49926] = 12'h100;
rom[49927] = 12'h100;
rom[49928] = 12'h100;
rom[49929] = 12'h100;
rom[49930] = 12'h100;
rom[49931] = 12'h100;
rom[49932] = 12'h100;
rom[49933] = 12'h100;
rom[49934] = 12'h100;
rom[49935] = 12'h100;
rom[49936] = 12'h100;
rom[49937] = 12'h201;
rom[49938] = 12'h211;
rom[49939] = 12'h212;
rom[49940] = 12'h322;
rom[49941] = 12'h332;
rom[49942] = 12'h433;
rom[49943] = 12'h443;
rom[49944] = 12'h443;
rom[49945] = 12'h544;
rom[49946] = 12'h544;
rom[49947] = 12'h544;
rom[49948] = 12'h544;
rom[49949] = 12'h544;
rom[49950] = 12'h554;
rom[49951] = 12'h555;
rom[49952] = 12'h555;
rom[49953] = 12'h555;
rom[49954] = 12'h555;
rom[49955] = 12'h555;
rom[49956] = 12'h565;
rom[49957] = 12'h666;
rom[49958] = 12'h666;
rom[49959] = 12'h666;
rom[49960] = 12'h676;
rom[49961] = 12'h677;
rom[49962] = 12'h777;
rom[49963] = 12'h777;
rom[49964] = 12'h777;
rom[49965] = 12'h888;
rom[49966] = 12'h888;
rom[49967] = 12'h989;
rom[49968] = 12'h999;
rom[49969] = 12'h999;
rom[49970] = 12'haaa;
rom[49971] = 12'haab;
rom[49972] = 12'hbbb;
rom[49973] = 12'hccc;
rom[49974] = 12'hccc;
rom[49975] = 12'hccc;
rom[49976] = 12'hddd;
rom[49977] = 12'hddd;
rom[49978] = 12'hccc;
rom[49979] = 12'hccc;
rom[49980] = 12'hccb;
rom[49981] = 12'hbbb;
rom[49982] = 12'hbbb;
rom[49983] = 12'hbbb;
rom[49984] = 12'hbbb;
rom[49985] = 12'hbbb;
rom[49986] = 12'hbbb;
rom[49987] = 12'hbbb;
rom[49988] = 12'hbbb;
rom[49989] = 12'hbbb;
rom[49990] = 12'hbbb;
rom[49991] = 12'hbbb;
rom[49992] = 12'hbbb;
rom[49993] = 12'hbbb;
rom[49994] = 12'hbbb;
rom[49995] = 12'hbbb;
rom[49996] = 12'hbbb;
rom[49997] = 12'hbbb;
rom[49998] = 12'hbbb;
rom[49999] = 12'hbbb;
rom[50000] = 12'hbbb;
rom[50001] = 12'haaa;
rom[50002] = 12'haaa;
rom[50003] = 12'haaa;
rom[50004] = 12'h999;
rom[50005] = 12'h999;
rom[50006] = 12'h999;
rom[50007] = 12'h888;
rom[50008] = 12'h888;
rom[50009] = 12'h888;
rom[50010] = 12'h888;
rom[50011] = 12'h888;
rom[50012] = 12'h777;
rom[50013] = 12'h777;
rom[50014] = 12'h777;
rom[50015] = 12'h777;
rom[50016] = 12'h888;
rom[50017] = 12'h888;
rom[50018] = 12'h888;
rom[50019] = 12'h888;
rom[50020] = 12'h888;
rom[50021] = 12'h888;
rom[50022] = 12'h888;
rom[50023] = 12'h888;
rom[50024] = 12'h888;
rom[50025] = 12'h888;
rom[50026] = 12'h888;
rom[50027] = 12'h888;
rom[50028] = 12'h888;
rom[50029] = 12'h888;
rom[50030] = 12'h888;
rom[50031] = 12'h888;
rom[50032] = 12'h888;
rom[50033] = 12'h888;
rom[50034] = 12'h888;
rom[50035] = 12'h888;
rom[50036] = 12'h888;
rom[50037] = 12'h888;
rom[50038] = 12'h888;
rom[50039] = 12'h888;
rom[50040] = 12'h888;
rom[50041] = 12'h888;
rom[50042] = 12'h888;
rom[50043] = 12'h888;
rom[50044] = 12'h888;
rom[50045] = 12'h888;
rom[50046] = 12'h888;
rom[50047] = 12'h888;
rom[50048] = 12'h888;
rom[50049] = 12'h888;
rom[50050] = 12'h888;
rom[50051] = 12'h888;
rom[50052] = 12'h888;
rom[50053] = 12'h999;
rom[50054] = 12'h999;
rom[50055] = 12'h999;
rom[50056] = 12'h999;
rom[50057] = 12'h999;
rom[50058] = 12'h999;
rom[50059] = 12'h999;
rom[50060] = 12'h999;
rom[50061] = 12'haaa;
rom[50062] = 12'haaa;
rom[50063] = 12'haaa;
rom[50064] = 12'haaa;
rom[50065] = 12'haaa;
rom[50066] = 12'haaa;
rom[50067] = 12'hbbb;
rom[50068] = 12'hbbb;
rom[50069] = 12'hbbb;
rom[50070] = 12'hbbb;
rom[50071] = 12'hbbb;
rom[50072] = 12'haaa;
rom[50073] = 12'h999;
rom[50074] = 12'h999;
rom[50075] = 12'h888;
rom[50076] = 12'h888;
rom[50077] = 12'h888;
rom[50078] = 12'h888;
rom[50079] = 12'h888;
rom[50080] = 12'h888;
rom[50081] = 12'h888;
rom[50082] = 12'h888;
rom[50083] = 12'h888;
rom[50084] = 12'h888;
rom[50085] = 12'h888;
rom[50086] = 12'h888;
rom[50087] = 12'h888;
rom[50088] = 12'h888;
rom[50089] = 12'h888;
rom[50090] = 12'h777;
rom[50091] = 12'h777;
rom[50092] = 12'h777;
rom[50093] = 12'h777;
rom[50094] = 12'h666;
rom[50095] = 12'h666;
rom[50096] = 12'h777;
rom[50097] = 12'h666;
rom[50098] = 12'h666;
rom[50099] = 12'h666;
rom[50100] = 12'h666;
rom[50101] = 12'h666;
rom[50102] = 12'h666;
rom[50103] = 12'h666;
rom[50104] = 12'h666;
rom[50105] = 12'h666;
rom[50106] = 12'h555;
rom[50107] = 12'h555;
rom[50108] = 12'h444;
rom[50109] = 12'h444;
rom[50110] = 12'h444;
rom[50111] = 12'h444;
rom[50112] = 12'h444;
rom[50113] = 12'h444;
rom[50114] = 12'h444;
rom[50115] = 12'h444;
rom[50116] = 12'h333;
rom[50117] = 12'h333;
rom[50118] = 12'h222;
rom[50119] = 12'h222;
rom[50120] = 12'h222;
rom[50121] = 12'h111;
rom[50122] = 12'h111;
rom[50123] = 12'h111;
rom[50124] = 12'h111;
rom[50125] = 12'h111;
rom[50126] = 12'h  0;
rom[50127] = 12'h  0;
rom[50128] = 12'h  0;
rom[50129] = 12'h  0;
rom[50130] = 12'h  0;
rom[50131] = 12'h  0;
rom[50132] = 12'h  0;
rom[50133] = 12'h  0;
rom[50134] = 12'h  0;
rom[50135] = 12'h  0;
rom[50136] = 12'h  0;
rom[50137] = 12'h  0;
rom[50138] = 12'h  0;
rom[50139] = 12'h  0;
rom[50140] = 12'h  0;
rom[50141] = 12'h  0;
rom[50142] = 12'h  0;
rom[50143] = 12'h  0;
rom[50144] = 12'h  0;
rom[50145] = 12'h  0;
rom[50146] = 12'h  0;
rom[50147] = 12'h111;
rom[50148] = 12'h111;
rom[50149] = 12'h111;
rom[50150] = 12'h111;
rom[50151] = 12'h111;
rom[50152] = 12'h111;
rom[50153] = 12'h111;
rom[50154] = 12'h111;
rom[50155] = 12'h111;
rom[50156] = 12'h111;
rom[50157] = 12'h111;
rom[50158] = 12'h111;
rom[50159] = 12'h111;
rom[50160] = 12'h111;
rom[50161] = 12'h111;
rom[50162] = 12'h111;
rom[50163] = 12'h111;
rom[50164] = 12'h111;
rom[50165] = 12'h111;
rom[50166] = 12'h111;
rom[50167] = 12'h111;
rom[50168] = 12'h111;
rom[50169] = 12'h111;
rom[50170] = 12'h111;
rom[50171] = 12'h111;
rom[50172] = 12'h111;
rom[50173] = 12'h111;
rom[50174] = 12'h111;
rom[50175] = 12'h111;
rom[50176] = 12'h111;
rom[50177] = 12'h111;
rom[50178] = 12'h111;
rom[50179] = 12'h111;
rom[50180] = 12'h111;
rom[50181] = 12'h111;
rom[50182] = 12'h111;
rom[50183] = 12'h  0;
rom[50184] = 12'h  0;
rom[50185] = 12'h  0;
rom[50186] = 12'h  0;
rom[50187] = 12'h  0;
rom[50188] = 12'h  0;
rom[50189] = 12'h  0;
rom[50190] = 12'h  0;
rom[50191] = 12'h  0;
rom[50192] = 12'h  0;
rom[50193] = 12'h  0;
rom[50194] = 12'h  0;
rom[50195] = 12'h  0;
rom[50196] = 12'h  0;
rom[50197] = 12'h  0;
rom[50198] = 12'h  0;
rom[50199] = 12'h  0;
rom[50200] = 12'h  0;
rom[50201] = 12'h  0;
rom[50202] = 12'h  0;
rom[50203] = 12'h  0;
rom[50204] = 12'h  0;
rom[50205] = 12'h  0;
rom[50206] = 12'h  0;
rom[50207] = 12'h  0;
rom[50208] = 12'h111;
rom[50209] = 12'h111;
rom[50210] = 12'h111;
rom[50211] = 12'h111;
rom[50212] = 12'h  0;
rom[50213] = 12'h  0;
rom[50214] = 12'h111;
rom[50215] = 12'h111;
rom[50216] = 12'h111;
rom[50217] = 12'h111;
rom[50218] = 12'h111;
rom[50219] = 12'h111;
rom[50220] = 12'h111;
rom[50221] = 12'h111;
rom[50222] = 12'h222;
rom[50223] = 12'h222;
rom[50224] = 12'h222;
rom[50225] = 12'h222;
rom[50226] = 12'h222;
rom[50227] = 12'h222;
rom[50228] = 12'h222;
rom[50229] = 12'h111;
rom[50230] = 12'h111;
rom[50231] = 12'h111;
rom[50232] = 12'h111;
rom[50233] = 12'h111;
rom[50234] = 12'h111;
rom[50235] = 12'h  0;
rom[50236] = 12'h  0;
rom[50237] = 12'h  0;
rom[50238] = 12'h  0;
rom[50239] = 12'h  0;
rom[50240] = 12'h  0;
rom[50241] = 12'h  0;
rom[50242] = 12'h  0;
rom[50243] = 12'h  0;
rom[50244] = 12'h  0;
rom[50245] = 12'h  0;
rom[50246] = 12'h  0;
rom[50247] = 12'h  0;
rom[50248] = 12'h  0;
rom[50249] = 12'h  0;
rom[50250] = 12'h  0;
rom[50251] = 12'h  0;
rom[50252] = 12'h  0;
rom[50253] = 12'h  0;
rom[50254] = 12'h  0;
rom[50255] = 12'h  0;
rom[50256] = 12'h  0;
rom[50257] = 12'h  0;
rom[50258] = 12'h  0;
rom[50259] = 12'h  0;
rom[50260] = 12'h  0;
rom[50261] = 12'h  0;
rom[50262] = 12'h  0;
rom[50263] = 12'h  0;
rom[50264] = 12'h  0;
rom[50265] = 12'h  0;
rom[50266] = 12'h  0;
rom[50267] = 12'h  0;
rom[50268] = 12'h  0;
rom[50269] = 12'h111;
rom[50270] = 12'h111;
rom[50271] = 12'h111;
rom[50272] = 12'h111;
rom[50273] = 12'h111;
rom[50274] = 12'h222;
rom[50275] = 12'h333;
rom[50276] = 12'h444;
rom[50277] = 12'h444;
rom[50278] = 12'h444;
rom[50279] = 12'h444;
rom[50280] = 12'h333;
rom[50281] = 12'h444;
rom[50282] = 12'h444;
rom[50283] = 12'h444;
rom[50284] = 12'h555;
rom[50285] = 12'h555;
rom[50286] = 12'h666;
rom[50287] = 12'h666;
rom[50288] = 12'h777;
rom[50289] = 12'h777;
rom[50290] = 12'h777;
rom[50291] = 12'h666;
rom[50292] = 12'h666;
rom[50293] = 12'h777;
rom[50294] = 12'h788;
rom[50295] = 12'h888;
rom[50296] = 12'h788;
rom[50297] = 12'h777;
rom[50298] = 12'h666;
rom[50299] = 12'h665;
rom[50300] = 12'h555;
rom[50301] = 12'h444;
rom[50302] = 12'h333;
rom[50303] = 12'h222;
rom[50304] = 12'h211;
rom[50305] = 12'h111;
rom[50306] = 12'h100;
rom[50307] = 12'h100;
rom[50308] = 12'h  0;
rom[50309] = 12'h  0;
rom[50310] = 12'h  0;
rom[50311] = 12'h  0;
rom[50312] = 12'h100;
rom[50313] = 12'h100;
rom[50314] = 12'h100;
rom[50315] = 12'h100;
rom[50316] = 12'h100;
rom[50317] = 12'h100;
rom[50318] = 12'h100;
rom[50319] = 12'h100;
rom[50320] = 12'h100;
rom[50321] = 12'h100;
rom[50322] = 12'h100;
rom[50323] = 12'h100;
rom[50324] = 12'h100;
rom[50325] = 12'h100;
rom[50326] = 12'h100;
rom[50327] = 12'h100;
rom[50328] = 12'h100;
rom[50329] = 12'h100;
rom[50330] = 12'h100;
rom[50331] = 12'h100;
rom[50332] = 12'h100;
rom[50333] = 12'h100;
rom[50334] = 12'h100;
rom[50335] = 12'h111;
rom[50336] = 12'h211;
rom[50337] = 12'h211;
rom[50338] = 12'h322;
rom[50339] = 12'h333;
rom[50340] = 12'h433;
rom[50341] = 12'h443;
rom[50342] = 12'h544;
rom[50343] = 12'h544;
rom[50344] = 12'h544;
rom[50345] = 12'h544;
rom[50346] = 12'h544;
rom[50347] = 12'h544;
rom[50348] = 12'h544;
rom[50349] = 12'h554;
rom[50350] = 12'h555;
rom[50351] = 12'h555;
rom[50352] = 12'h555;
rom[50353] = 12'h555;
rom[50354] = 12'h555;
rom[50355] = 12'h555;
rom[50356] = 12'h666;
rom[50357] = 12'h666;
rom[50358] = 12'h666;
rom[50359] = 12'h666;
rom[50360] = 12'h777;
rom[50361] = 12'h777;
rom[50362] = 12'h777;
rom[50363] = 12'h777;
rom[50364] = 12'h888;
rom[50365] = 12'h888;
rom[50366] = 12'h989;
rom[50367] = 12'h999;
rom[50368] = 12'h99a;
rom[50369] = 12'haaa;
rom[50370] = 12'haab;
rom[50371] = 12'hbbb;
rom[50372] = 12'hbbc;
rom[50373] = 12'hccc;
rom[50374] = 12'hddd;
rom[50375] = 12'hddd;
rom[50376] = 12'hddd;
rom[50377] = 12'hccc;
rom[50378] = 12'hccc;
rom[50379] = 12'hccb;
rom[50380] = 12'hccb;
rom[50381] = 12'hbcb;
rom[50382] = 12'hbbb;
rom[50383] = 12'hbbb;
rom[50384] = 12'hbbb;
rom[50385] = 12'hbbb;
rom[50386] = 12'hbbb;
rom[50387] = 12'hbbb;
rom[50388] = 12'hbbb;
rom[50389] = 12'hbbb;
rom[50390] = 12'hbbb;
rom[50391] = 12'hbbb;
rom[50392] = 12'hbbb;
rom[50393] = 12'hbbb;
rom[50394] = 12'hbbb;
rom[50395] = 12'hbbb;
rom[50396] = 12'hbbb;
rom[50397] = 12'hbbb;
rom[50398] = 12'hbbb;
rom[50399] = 12'hbbb;
rom[50400] = 12'hbbb;
rom[50401] = 12'hbbb;
rom[50402] = 12'haaa;
rom[50403] = 12'haaa;
rom[50404] = 12'haaa;
rom[50405] = 12'h999;
rom[50406] = 12'h999;
rom[50407] = 12'h999;
rom[50408] = 12'h888;
rom[50409] = 12'h888;
rom[50410] = 12'h888;
rom[50411] = 12'h888;
rom[50412] = 12'h888;
rom[50413] = 12'h888;
rom[50414] = 12'h888;
rom[50415] = 12'h888;
rom[50416] = 12'h888;
rom[50417] = 12'h888;
rom[50418] = 12'h888;
rom[50419] = 12'h888;
rom[50420] = 12'h888;
rom[50421] = 12'h888;
rom[50422] = 12'h888;
rom[50423] = 12'h888;
rom[50424] = 12'h888;
rom[50425] = 12'h999;
rom[50426] = 12'h999;
rom[50427] = 12'h999;
rom[50428] = 12'h999;
rom[50429] = 12'h999;
rom[50430] = 12'h888;
rom[50431] = 12'h888;
rom[50432] = 12'h888;
rom[50433] = 12'h888;
rom[50434] = 12'h888;
rom[50435] = 12'h888;
rom[50436] = 12'h888;
rom[50437] = 12'h888;
rom[50438] = 12'h888;
rom[50439] = 12'h888;
rom[50440] = 12'h888;
rom[50441] = 12'h888;
rom[50442] = 12'h888;
rom[50443] = 12'h888;
rom[50444] = 12'h888;
rom[50445] = 12'h888;
rom[50446] = 12'h888;
rom[50447] = 12'h888;
rom[50448] = 12'h888;
rom[50449] = 12'h888;
rom[50450] = 12'h888;
rom[50451] = 12'h999;
rom[50452] = 12'h999;
rom[50453] = 12'h999;
rom[50454] = 12'h999;
rom[50455] = 12'h999;
rom[50456] = 12'h999;
rom[50457] = 12'h999;
rom[50458] = 12'h999;
rom[50459] = 12'h999;
rom[50460] = 12'haaa;
rom[50461] = 12'haaa;
rom[50462] = 12'haaa;
rom[50463] = 12'haaa;
rom[50464] = 12'hbbb;
rom[50465] = 12'hbbb;
rom[50466] = 12'hbbb;
rom[50467] = 12'hbbb;
rom[50468] = 12'hbbb;
rom[50469] = 12'hbbb;
rom[50470] = 12'hbbb;
rom[50471] = 12'hbbb;
rom[50472] = 12'haaa;
rom[50473] = 12'haaa;
rom[50474] = 12'h999;
rom[50475] = 12'h999;
rom[50476] = 12'h888;
rom[50477] = 12'h888;
rom[50478] = 12'h888;
rom[50479] = 12'h888;
rom[50480] = 12'h888;
rom[50481] = 12'h888;
rom[50482] = 12'h777;
rom[50483] = 12'h777;
rom[50484] = 12'h888;
rom[50485] = 12'h888;
rom[50486] = 12'h888;
rom[50487] = 12'h888;
rom[50488] = 12'h888;
rom[50489] = 12'h888;
rom[50490] = 12'h777;
rom[50491] = 12'h777;
rom[50492] = 12'h777;
rom[50493] = 12'h777;
rom[50494] = 12'h777;
rom[50495] = 12'h777;
rom[50496] = 12'h777;
rom[50497] = 12'h777;
rom[50498] = 12'h666;
rom[50499] = 12'h666;
rom[50500] = 12'h666;
rom[50501] = 12'h666;
rom[50502] = 12'h666;
rom[50503] = 12'h666;
rom[50504] = 12'h666;
rom[50505] = 12'h666;
rom[50506] = 12'h666;
rom[50507] = 12'h555;
rom[50508] = 12'h555;
rom[50509] = 12'h555;
rom[50510] = 12'h444;
rom[50511] = 12'h444;
rom[50512] = 12'h444;
rom[50513] = 12'h444;
rom[50514] = 12'h444;
rom[50515] = 12'h444;
rom[50516] = 12'h444;
rom[50517] = 12'h444;
rom[50518] = 12'h333;
rom[50519] = 12'h333;
rom[50520] = 12'h222;
rom[50521] = 12'h222;
rom[50522] = 12'h111;
rom[50523] = 12'h111;
rom[50524] = 12'h111;
rom[50525] = 12'h111;
rom[50526] = 12'h111;
rom[50527] = 12'h111;
rom[50528] = 12'h111;
rom[50529] = 12'h111;
rom[50530] = 12'h111;
rom[50531] = 12'h111;
rom[50532] = 12'h111;
rom[50533] = 12'h111;
rom[50534] = 12'h  0;
rom[50535] = 12'h  0;
rom[50536] = 12'h  0;
rom[50537] = 12'h  0;
rom[50538] = 12'h  0;
rom[50539] = 12'h  0;
rom[50540] = 12'h  0;
rom[50541] = 12'h  0;
rom[50542] = 12'h  0;
rom[50543] = 12'h  0;
rom[50544] = 12'h111;
rom[50545] = 12'h111;
rom[50546] = 12'h111;
rom[50547] = 12'h111;
rom[50548] = 12'h111;
rom[50549] = 12'h111;
rom[50550] = 12'h111;
rom[50551] = 12'h111;
rom[50552] = 12'h111;
rom[50553] = 12'h111;
rom[50554] = 12'h111;
rom[50555] = 12'h111;
rom[50556] = 12'h111;
rom[50557] = 12'h111;
rom[50558] = 12'h111;
rom[50559] = 12'h111;
rom[50560] = 12'h111;
rom[50561] = 12'h111;
rom[50562] = 12'h111;
rom[50563] = 12'h111;
rom[50564] = 12'h111;
rom[50565] = 12'h111;
rom[50566] = 12'h111;
rom[50567] = 12'h222;
rom[50568] = 12'h222;
rom[50569] = 12'h111;
rom[50570] = 12'h111;
rom[50571] = 12'h111;
rom[50572] = 12'h111;
rom[50573] = 12'h111;
rom[50574] = 12'h111;
rom[50575] = 12'h111;
rom[50576] = 12'h111;
rom[50577] = 12'h111;
rom[50578] = 12'h111;
rom[50579] = 12'h111;
rom[50580] = 12'h111;
rom[50581] = 12'h  0;
rom[50582] = 12'h  0;
rom[50583] = 12'h  0;
rom[50584] = 12'h  0;
rom[50585] = 12'h  0;
rom[50586] = 12'h  0;
rom[50587] = 12'h  0;
rom[50588] = 12'h  0;
rom[50589] = 12'h  0;
rom[50590] = 12'h  0;
rom[50591] = 12'h  0;
rom[50592] = 12'h  0;
rom[50593] = 12'h  0;
rom[50594] = 12'h  0;
rom[50595] = 12'h  0;
rom[50596] = 12'h  0;
rom[50597] = 12'h  0;
rom[50598] = 12'h  0;
rom[50599] = 12'h  0;
rom[50600] = 12'h  0;
rom[50601] = 12'h  0;
rom[50602] = 12'h  0;
rom[50603] = 12'h  0;
rom[50604] = 12'h  0;
rom[50605] = 12'h  0;
rom[50606] = 12'h  0;
rom[50607] = 12'h  0;
rom[50608] = 12'h111;
rom[50609] = 12'h111;
rom[50610] = 12'h111;
rom[50611] = 12'h  0;
rom[50612] = 12'h  0;
rom[50613] = 12'h  0;
rom[50614] = 12'h111;
rom[50615] = 12'h111;
rom[50616] = 12'h111;
rom[50617] = 12'h111;
rom[50618] = 12'h111;
rom[50619] = 12'h111;
rom[50620] = 12'h111;
rom[50621] = 12'h111;
rom[50622] = 12'h222;
rom[50623] = 12'h222;
rom[50624] = 12'h222;
rom[50625] = 12'h222;
rom[50626] = 12'h222;
rom[50627] = 12'h222;
rom[50628] = 12'h222;
rom[50629] = 12'h111;
rom[50630] = 12'h111;
rom[50631] = 12'h111;
rom[50632] = 12'h111;
rom[50633] = 12'h111;
rom[50634] = 12'h  0;
rom[50635] = 12'h  0;
rom[50636] = 12'h  0;
rom[50637] = 12'h  0;
rom[50638] = 12'h  0;
rom[50639] = 12'h  0;
rom[50640] = 12'h  0;
rom[50641] = 12'h  0;
rom[50642] = 12'h  0;
rom[50643] = 12'h  0;
rom[50644] = 12'h  0;
rom[50645] = 12'h  0;
rom[50646] = 12'h  0;
rom[50647] = 12'h  0;
rom[50648] = 12'h  0;
rom[50649] = 12'h  0;
rom[50650] = 12'h  0;
rom[50651] = 12'h  0;
rom[50652] = 12'h  0;
rom[50653] = 12'h  0;
rom[50654] = 12'h  0;
rom[50655] = 12'h  0;
rom[50656] = 12'h  0;
rom[50657] = 12'h  0;
rom[50658] = 12'h  0;
rom[50659] = 12'h  0;
rom[50660] = 12'h  0;
rom[50661] = 12'h  0;
rom[50662] = 12'h  0;
rom[50663] = 12'h  0;
rom[50664] = 12'h  0;
rom[50665] = 12'h  0;
rom[50666] = 12'h  0;
rom[50667] = 12'h  0;
rom[50668] = 12'h  0;
rom[50669] = 12'h111;
rom[50670] = 12'h111;
rom[50671] = 12'h111;
rom[50672] = 12'h111;
rom[50673] = 12'h111;
rom[50674] = 12'h222;
rom[50675] = 12'h333;
rom[50676] = 12'h444;
rom[50677] = 12'h444;
rom[50678] = 12'h444;
rom[50679] = 12'h444;
rom[50680] = 12'h444;
rom[50681] = 12'h444;
rom[50682] = 12'h444;
rom[50683] = 12'h444;
rom[50684] = 12'h555;
rom[50685] = 12'h555;
rom[50686] = 12'h666;
rom[50687] = 12'h666;
rom[50688] = 12'h777;
rom[50689] = 12'h777;
rom[50690] = 12'h666;
rom[50691] = 12'h666;
rom[50692] = 12'h666;
rom[50693] = 12'h777;
rom[50694] = 12'h787;
rom[50695] = 12'h787;
rom[50696] = 12'h777;
rom[50697] = 12'h777;
rom[50698] = 12'h677;
rom[50699] = 12'h666;
rom[50700] = 12'h655;
rom[50701] = 12'h555;
rom[50702] = 12'h444;
rom[50703] = 12'h333;
rom[50704] = 12'h222;
rom[50705] = 12'h222;
rom[50706] = 12'h111;
rom[50707] = 12'h100;
rom[50708] = 12'h  0;
rom[50709] = 12'h  0;
rom[50710] = 12'h  0;
rom[50711] = 12'h  0;
rom[50712] = 12'h  0;
rom[50713] = 12'h  0;
rom[50714] = 12'h  0;
rom[50715] = 12'h  0;
rom[50716] = 12'h  0;
rom[50717] = 12'h100;
rom[50718] = 12'h100;
rom[50719] = 12'h100;
rom[50720] = 12'h100;
rom[50721] = 12'h100;
rom[50722] = 12'h100;
rom[50723] = 12'h100;
rom[50724] = 12'h100;
rom[50725] = 12'h100;
rom[50726] = 12'h100;
rom[50727] = 12'h100;
rom[50728] = 12'h100;
rom[50729] = 12'h100;
rom[50730] = 12'h100;
rom[50731] = 12'h100;
rom[50732] = 12'h111;
rom[50733] = 12'h111;
rom[50734] = 12'h211;
rom[50735] = 12'h222;
rom[50736] = 12'h322;
rom[50737] = 12'h323;
rom[50738] = 12'h433;
rom[50739] = 12'h433;
rom[50740] = 12'h444;
rom[50741] = 12'h444;
rom[50742] = 12'h544;
rom[50743] = 12'h544;
rom[50744] = 12'h544;
rom[50745] = 12'h554;
rom[50746] = 12'h554;
rom[50747] = 12'h554;
rom[50748] = 12'h554;
rom[50749] = 12'h555;
rom[50750] = 12'h555;
rom[50751] = 12'h555;
rom[50752] = 12'h555;
rom[50753] = 12'h655;
rom[50754] = 12'h665;
rom[50755] = 12'h666;
rom[50756] = 12'h666;
rom[50757] = 12'h666;
rom[50758] = 12'h676;
rom[50759] = 12'h777;
rom[50760] = 12'h777;
rom[50761] = 12'h787;
rom[50762] = 12'h888;
rom[50763] = 12'h888;
rom[50764] = 12'h888;
rom[50765] = 12'h999;
rom[50766] = 12'ha99;
rom[50767] = 12'haaa;
rom[50768] = 12'haaa;
rom[50769] = 12'haab;
rom[50770] = 12'hbbb;
rom[50771] = 12'hbbc;
rom[50772] = 12'hccc;
rom[50773] = 12'hddd;
rom[50774] = 12'hddd;
rom[50775] = 12'hddd;
rom[50776] = 12'hcdd;
rom[50777] = 12'hccc;
rom[50778] = 12'hccc;
rom[50779] = 12'hccb;
rom[50780] = 12'hccb;
rom[50781] = 12'hccb;
rom[50782] = 12'hbcb;
rom[50783] = 12'hbcb;
rom[50784] = 12'hccb;
rom[50785] = 12'hccc;
rom[50786] = 12'hccc;
rom[50787] = 12'hccc;
rom[50788] = 12'hccc;
rom[50789] = 12'hccc;
rom[50790] = 12'hccc;
rom[50791] = 12'hccc;
rom[50792] = 12'hbbb;
rom[50793] = 12'hbbb;
rom[50794] = 12'hbbb;
rom[50795] = 12'hbbb;
rom[50796] = 12'hbbb;
rom[50797] = 12'hbbb;
rom[50798] = 12'hbbb;
rom[50799] = 12'hbbb;
rom[50800] = 12'hbbb;
rom[50801] = 12'hbbb;
rom[50802] = 12'hbbb;
rom[50803] = 12'haaa;
rom[50804] = 12'haaa;
rom[50805] = 12'haaa;
rom[50806] = 12'h999;
rom[50807] = 12'h999;
rom[50808] = 12'h999;
rom[50809] = 12'h888;
rom[50810] = 12'h888;
rom[50811] = 12'h888;
rom[50812] = 12'h888;
rom[50813] = 12'h888;
rom[50814] = 12'h888;
rom[50815] = 12'h888;
rom[50816] = 12'h888;
rom[50817] = 12'h888;
rom[50818] = 12'h888;
rom[50819] = 12'h888;
rom[50820] = 12'h888;
rom[50821] = 12'h888;
rom[50822] = 12'h888;
rom[50823] = 12'h888;
rom[50824] = 12'h999;
rom[50825] = 12'h999;
rom[50826] = 12'h999;
rom[50827] = 12'h999;
rom[50828] = 12'h999;
rom[50829] = 12'h999;
rom[50830] = 12'h888;
rom[50831] = 12'h888;
rom[50832] = 12'h888;
rom[50833] = 12'h888;
rom[50834] = 12'h888;
rom[50835] = 12'h888;
rom[50836] = 12'h888;
rom[50837] = 12'h888;
rom[50838] = 12'h999;
rom[50839] = 12'h999;
rom[50840] = 12'h888;
rom[50841] = 12'h888;
rom[50842] = 12'h888;
rom[50843] = 12'h888;
rom[50844] = 12'h888;
rom[50845] = 12'h888;
rom[50846] = 12'h888;
rom[50847] = 12'h888;
rom[50848] = 12'h888;
rom[50849] = 12'h888;
rom[50850] = 12'h999;
rom[50851] = 12'h999;
rom[50852] = 12'h999;
rom[50853] = 12'h999;
rom[50854] = 12'h999;
rom[50855] = 12'h999;
rom[50856] = 12'h999;
rom[50857] = 12'h999;
rom[50858] = 12'h999;
rom[50859] = 12'h999;
rom[50860] = 12'haaa;
rom[50861] = 12'haaa;
rom[50862] = 12'haaa;
rom[50863] = 12'haaa;
rom[50864] = 12'hbbb;
rom[50865] = 12'hbbb;
rom[50866] = 12'hbbb;
rom[50867] = 12'hbbb;
rom[50868] = 12'hbbb;
rom[50869] = 12'hbbb;
rom[50870] = 12'hbbb;
rom[50871] = 12'hbbb;
rom[50872] = 12'haaa;
rom[50873] = 12'haaa;
rom[50874] = 12'h999;
rom[50875] = 12'h999;
rom[50876] = 12'h999;
rom[50877] = 12'h999;
rom[50878] = 12'h888;
rom[50879] = 12'h888;
rom[50880] = 12'h888;
rom[50881] = 12'h777;
rom[50882] = 12'h777;
rom[50883] = 12'h777;
rom[50884] = 12'h777;
rom[50885] = 12'h777;
rom[50886] = 12'h777;
rom[50887] = 12'h777;
rom[50888] = 12'h777;
rom[50889] = 12'h777;
rom[50890] = 12'h777;
rom[50891] = 12'h777;
rom[50892] = 12'h777;
rom[50893] = 12'h777;
rom[50894] = 12'h777;
rom[50895] = 12'h777;
rom[50896] = 12'h777;
rom[50897] = 12'h777;
rom[50898] = 12'h777;
rom[50899] = 12'h777;
rom[50900] = 12'h777;
rom[50901] = 12'h666;
rom[50902] = 12'h666;
rom[50903] = 12'h666;
rom[50904] = 12'h777;
rom[50905] = 12'h666;
rom[50906] = 12'h666;
rom[50907] = 12'h666;
rom[50908] = 12'h666;
rom[50909] = 12'h555;
rom[50910] = 12'h555;
rom[50911] = 12'h444;
rom[50912] = 12'h444;
rom[50913] = 12'h444;
rom[50914] = 12'h444;
rom[50915] = 12'h444;
rom[50916] = 12'h555;
rom[50917] = 12'h555;
rom[50918] = 12'h444;
rom[50919] = 12'h333;
rom[50920] = 12'h333;
rom[50921] = 12'h222;
rom[50922] = 12'h222;
rom[50923] = 12'h111;
rom[50924] = 12'h111;
rom[50925] = 12'h111;
rom[50926] = 12'h111;
rom[50927] = 12'h111;
rom[50928] = 12'h111;
rom[50929] = 12'h111;
rom[50930] = 12'h111;
rom[50931] = 12'h111;
rom[50932] = 12'h111;
rom[50933] = 12'h111;
rom[50934] = 12'h  0;
rom[50935] = 12'h  0;
rom[50936] = 12'h  0;
rom[50937] = 12'h  0;
rom[50938] = 12'h  0;
rom[50939] = 12'h  0;
rom[50940] = 12'h  0;
rom[50941] = 12'h  0;
rom[50942] = 12'h  0;
rom[50943] = 12'h  0;
rom[50944] = 12'h111;
rom[50945] = 12'h111;
rom[50946] = 12'h111;
rom[50947] = 12'h111;
rom[50948] = 12'h111;
rom[50949] = 12'h111;
rom[50950] = 12'h111;
rom[50951] = 12'h111;
rom[50952] = 12'h111;
rom[50953] = 12'h111;
rom[50954] = 12'h111;
rom[50955] = 12'h111;
rom[50956] = 12'h111;
rom[50957] = 12'h111;
rom[50958] = 12'h111;
rom[50959] = 12'h111;
rom[50960] = 12'h111;
rom[50961] = 12'h111;
rom[50962] = 12'h111;
rom[50963] = 12'h111;
rom[50964] = 12'h111;
rom[50965] = 12'h111;
rom[50966] = 12'h111;
rom[50967] = 12'h222;
rom[50968] = 12'h222;
rom[50969] = 12'h222;
rom[50970] = 12'h111;
rom[50971] = 12'h111;
rom[50972] = 12'h111;
rom[50973] = 12'h111;
rom[50974] = 12'h111;
rom[50975] = 12'h222;
rom[50976] = 12'h111;
rom[50977] = 12'h111;
rom[50978] = 12'h111;
rom[50979] = 12'h111;
rom[50980] = 12'h111;
rom[50981] = 12'h  0;
rom[50982] = 12'h  0;
rom[50983] = 12'h  0;
rom[50984] = 12'h  0;
rom[50985] = 12'h  0;
rom[50986] = 12'h  0;
rom[50987] = 12'h  0;
rom[50988] = 12'h  0;
rom[50989] = 12'h  0;
rom[50990] = 12'h  0;
rom[50991] = 12'h  0;
rom[50992] = 12'h  0;
rom[50993] = 12'h  0;
rom[50994] = 12'h  0;
rom[50995] = 12'h  0;
rom[50996] = 12'h  0;
rom[50997] = 12'h  0;
rom[50998] = 12'h  0;
rom[50999] = 12'h  0;
rom[51000] = 12'h  0;
rom[51001] = 12'h  0;
rom[51002] = 12'h  0;
rom[51003] = 12'h  0;
rom[51004] = 12'h  0;
rom[51005] = 12'h  0;
rom[51006] = 12'h  0;
rom[51007] = 12'h  0;
rom[51008] = 12'h111;
rom[51009] = 12'h111;
rom[51010] = 12'h111;
rom[51011] = 12'h  0;
rom[51012] = 12'h  0;
rom[51013] = 12'h  0;
rom[51014] = 12'h111;
rom[51015] = 12'h111;
rom[51016] = 12'h111;
rom[51017] = 12'h111;
rom[51018] = 12'h111;
rom[51019] = 12'h111;
rom[51020] = 12'h111;
rom[51021] = 12'h111;
rom[51022] = 12'h222;
rom[51023] = 12'h222;
rom[51024] = 12'h222;
rom[51025] = 12'h222;
rom[51026] = 12'h222;
rom[51027] = 12'h222;
rom[51028] = 12'h222;
rom[51029] = 12'h111;
rom[51030] = 12'h111;
rom[51031] = 12'h111;
rom[51032] = 12'h111;
rom[51033] = 12'h111;
rom[51034] = 12'h  0;
rom[51035] = 12'h  0;
rom[51036] = 12'h  0;
rom[51037] = 12'h  0;
rom[51038] = 12'h  0;
rom[51039] = 12'h  0;
rom[51040] = 12'h  0;
rom[51041] = 12'h  0;
rom[51042] = 12'h  0;
rom[51043] = 12'h  0;
rom[51044] = 12'h  0;
rom[51045] = 12'h  0;
rom[51046] = 12'h  0;
rom[51047] = 12'h  0;
rom[51048] = 12'h  0;
rom[51049] = 12'h  0;
rom[51050] = 12'h  0;
rom[51051] = 12'h  0;
rom[51052] = 12'h  0;
rom[51053] = 12'h  0;
rom[51054] = 12'h  0;
rom[51055] = 12'h  0;
rom[51056] = 12'h  0;
rom[51057] = 12'h  0;
rom[51058] = 12'h  0;
rom[51059] = 12'h  0;
rom[51060] = 12'h  0;
rom[51061] = 12'h  0;
rom[51062] = 12'h  0;
rom[51063] = 12'h  0;
rom[51064] = 12'h  0;
rom[51065] = 12'h  0;
rom[51066] = 12'h  0;
rom[51067] = 12'h  0;
rom[51068] = 12'h  0;
rom[51069] = 12'h111;
rom[51070] = 12'h111;
rom[51071] = 12'h111;
rom[51072] = 12'h111;
rom[51073] = 12'h111;
rom[51074] = 12'h222;
rom[51075] = 12'h333;
rom[51076] = 12'h444;
rom[51077] = 12'h444;
rom[51078] = 12'h444;
rom[51079] = 12'h444;
rom[51080] = 12'h444;
rom[51081] = 12'h444;
rom[51082] = 12'h444;
rom[51083] = 12'h444;
rom[51084] = 12'h444;
rom[51085] = 12'h555;
rom[51086] = 12'h666;
rom[51087] = 12'h666;
rom[51088] = 12'h777;
rom[51089] = 12'h666;
rom[51090] = 12'h666;
rom[51091] = 12'h555;
rom[51092] = 12'h666;
rom[51093] = 12'h777;
rom[51094] = 12'h777;
rom[51095] = 12'h777;
rom[51096] = 12'h777;
rom[51097] = 12'h777;
rom[51098] = 12'h777;
rom[51099] = 12'h666;
rom[51100] = 12'h666;
rom[51101] = 12'h555;
rom[51102] = 12'h544;
rom[51103] = 12'h444;
rom[51104] = 12'h333;
rom[51105] = 12'h222;
rom[51106] = 12'h221;
rom[51107] = 12'h111;
rom[51108] = 12'h  0;
rom[51109] = 12'h  0;
rom[51110] = 12'h  0;
rom[51111] = 12'h  0;
rom[51112] = 12'h  0;
rom[51113] = 12'h  0;
rom[51114] = 12'h  0;
rom[51115] = 12'h  0;
rom[51116] = 12'h  0;
rom[51117] = 12'h  0;
rom[51118] = 12'h  0;
rom[51119] = 12'h  0;
rom[51120] = 12'h100;
rom[51121] = 12'h100;
rom[51122] = 12'h100;
rom[51123] = 12'h100;
rom[51124] = 12'h100;
rom[51125] = 12'h  0;
rom[51126] = 12'h  0;
rom[51127] = 12'h  0;
rom[51128] = 12'h  0;
rom[51129] = 12'h  0;
rom[51130] = 12'h100;
rom[51131] = 12'h111;
rom[51132] = 12'h111;
rom[51133] = 12'h222;
rom[51134] = 12'h222;
rom[51135] = 12'h322;
rom[51136] = 12'h333;
rom[51137] = 12'h433;
rom[51138] = 12'h444;
rom[51139] = 12'h444;
rom[51140] = 12'h444;
rom[51141] = 12'h444;
rom[51142] = 12'h444;
rom[51143] = 12'h444;
rom[51144] = 12'h554;
rom[51145] = 12'h554;
rom[51146] = 12'h555;
rom[51147] = 12'h555;
rom[51148] = 12'h555;
rom[51149] = 12'h555;
rom[51150] = 12'h555;
rom[51151] = 12'h555;
rom[51152] = 12'h666;
rom[51153] = 12'h666;
rom[51154] = 12'h666;
rom[51155] = 12'h666;
rom[51156] = 12'h666;
rom[51157] = 12'h777;
rom[51158] = 12'h777;
rom[51159] = 12'h777;
rom[51160] = 12'h887;
rom[51161] = 12'h888;
rom[51162] = 12'h888;
rom[51163] = 12'h888;
rom[51164] = 12'h999;
rom[51165] = 12'h999;
rom[51166] = 12'haaa;
rom[51167] = 12'haaa;
rom[51168] = 12'hbbb;
rom[51169] = 12'hbbb;
rom[51170] = 12'hbbc;
rom[51171] = 12'hccc;
rom[51172] = 12'hccd;
rom[51173] = 12'hddd;
rom[51174] = 12'hddd;
rom[51175] = 12'hddd;
rom[51176] = 12'hccc;
rom[51177] = 12'hccc;
rom[51178] = 12'hccc;
rom[51179] = 12'hccc;
rom[51180] = 12'hccc;
rom[51181] = 12'hccc;
rom[51182] = 12'hccc;
rom[51183] = 12'hbcb;
rom[51184] = 12'hccc;
rom[51185] = 12'hccc;
rom[51186] = 12'hccc;
rom[51187] = 12'hccc;
rom[51188] = 12'hccc;
rom[51189] = 12'hccc;
rom[51190] = 12'hccc;
rom[51191] = 12'hccc;
rom[51192] = 12'hbbb;
rom[51193] = 12'hbbb;
rom[51194] = 12'hccc;
rom[51195] = 12'hccc;
rom[51196] = 12'hccc;
rom[51197] = 12'hccc;
rom[51198] = 12'hccc;
rom[51199] = 12'hccc;
rom[51200] = 12'hccc;
rom[51201] = 12'hccc;
rom[51202] = 12'hbbb;
rom[51203] = 12'hbbb;
rom[51204] = 12'haaa;
rom[51205] = 12'haaa;
rom[51206] = 12'haaa;
rom[51207] = 12'h999;
rom[51208] = 12'h999;
rom[51209] = 12'h999;
rom[51210] = 12'h999;
rom[51211] = 12'h999;
rom[51212] = 12'h999;
rom[51213] = 12'h999;
rom[51214] = 12'h999;
rom[51215] = 12'h999;
rom[51216] = 12'h999;
rom[51217] = 12'h999;
rom[51218] = 12'h999;
rom[51219] = 12'h999;
rom[51220] = 12'h999;
rom[51221] = 12'h999;
rom[51222] = 12'h999;
rom[51223] = 12'h999;
rom[51224] = 12'h999;
rom[51225] = 12'h999;
rom[51226] = 12'h999;
rom[51227] = 12'h999;
rom[51228] = 12'h999;
rom[51229] = 12'h999;
rom[51230] = 12'h999;
rom[51231] = 12'h999;
rom[51232] = 12'h888;
rom[51233] = 12'h888;
rom[51234] = 12'h888;
rom[51235] = 12'h999;
rom[51236] = 12'h999;
rom[51237] = 12'h999;
rom[51238] = 12'h999;
rom[51239] = 12'h999;
rom[51240] = 12'h999;
rom[51241] = 12'h999;
rom[51242] = 12'h999;
rom[51243] = 12'h999;
rom[51244] = 12'h999;
rom[51245] = 12'h999;
rom[51246] = 12'h999;
rom[51247] = 12'h999;
rom[51248] = 12'h999;
rom[51249] = 12'h999;
rom[51250] = 12'h999;
rom[51251] = 12'h999;
rom[51252] = 12'h999;
rom[51253] = 12'h999;
rom[51254] = 12'h999;
rom[51255] = 12'h999;
rom[51256] = 12'h999;
rom[51257] = 12'haaa;
rom[51258] = 12'haaa;
rom[51259] = 12'haaa;
rom[51260] = 12'haaa;
rom[51261] = 12'haaa;
rom[51262] = 12'haaa;
rom[51263] = 12'haaa;
rom[51264] = 12'hbbb;
rom[51265] = 12'hbbb;
rom[51266] = 12'hbbb;
rom[51267] = 12'hbbb;
rom[51268] = 12'hbbb;
rom[51269] = 12'hbbb;
rom[51270] = 12'hbbb;
rom[51271] = 12'hccc;
rom[51272] = 12'hbbb;
rom[51273] = 12'haaa;
rom[51274] = 12'haaa;
rom[51275] = 12'haaa;
rom[51276] = 12'h999;
rom[51277] = 12'h999;
rom[51278] = 12'h999;
rom[51279] = 12'h888;
rom[51280] = 12'h888;
rom[51281] = 12'h777;
rom[51282] = 12'h777;
rom[51283] = 12'h777;
rom[51284] = 12'h777;
rom[51285] = 12'h777;
rom[51286] = 12'h777;
rom[51287] = 12'h777;
rom[51288] = 12'h777;
rom[51289] = 12'h777;
rom[51290] = 12'h777;
rom[51291] = 12'h777;
rom[51292] = 12'h777;
rom[51293] = 12'h777;
rom[51294] = 12'h777;
rom[51295] = 12'h777;
rom[51296] = 12'h777;
rom[51297] = 12'h777;
rom[51298] = 12'h777;
rom[51299] = 12'h777;
rom[51300] = 12'h777;
rom[51301] = 12'h777;
rom[51302] = 12'h777;
rom[51303] = 12'h777;
rom[51304] = 12'h777;
rom[51305] = 12'h777;
rom[51306] = 12'h777;
rom[51307] = 12'h666;
rom[51308] = 12'h666;
rom[51309] = 12'h666;
rom[51310] = 12'h555;
rom[51311] = 12'h555;
rom[51312] = 12'h555;
rom[51313] = 12'h444;
rom[51314] = 12'h444;
rom[51315] = 12'h444;
rom[51316] = 12'h444;
rom[51317] = 12'h444;
rom[51318] = 12'h444;
rom[51319] = 12'h444;
rom[51320] = 12'h444;
rom[51321] = 12'h333;
rom[51322] = 12'h222;
rom[51323] = 12'h222;
rom[51324] = 12'h111;
rom[51325] = 12'h111;
rom[51326] = 12'h222;
rom[51327] = 12'h222;
rom[51328] = 12'h111;
rom[51329] = 12'h111;
rom[51330] = 12'h111;
rom[51331] = 12'h111;
rom[51332] = 12'h111;
rom[51333] = 12'h111;
rom[51334] = 12'h111;
rom[51335] = 12'h111;
rom[51336] = 12'h111;
rom[51337] = 12'h111;
rom[51338] = 12'h  0;
rom[51339] = 12'h  0;
rom[51340] = 12'h  0;
rom[51341] = 12'h111;
rom[51342] = 12'h111;
rom[51343] = 12'h111;
rom[51344] = 12'h111;
rom[51345] = 12'h111;
rom[51346] = 12'h111;
rom[51347] = 12'h111;
rom[51348] = 12'h111;
rom[51349] = 12'h111;
rom[51350] = 12'h111;
rom[51351] = 12'h111;
rom[51352] = 12'h111;
rom[51353] = 12'h111;
rom[51354] = 12'h111;
rom[51355] = 12'h111;
rom[51356] = 12'h111;
rom[51357] = 12'h111;
rom[51358] = 12'h111;
rom[51359] = 12'h111;
rom[51360] = 12'h111;
rom[51361] = 12'h111;
rom[51362] = 12'h111;
rom[51363] = 12'h111;
rom[51364] = 12'h111;
rom[51365] = 12'h111;
rom[51366] = 12'h111;
rom[51367] = 12'h111;
rom[51368] = 12'h222;
rom[51369] = 12'h111;
rom[51370] = 12'h111;
rom[51371] = 12'h111;
rom[51372] = 12'h111;
rom[51373] = 12'h111;
rom[51374] = 12'h111;
rom[51375] = 12'h111;
rom[51376] = 12'h111;
rom[51377] = 12'h111;
rom[51378] = 12'h111;
rom[51379] = 12'h  0;
rom[51380] = 12'h  0;
rom[51381] = 12'h  0;
rom[51382] = 12'h  0;
rom[51383] = 12'h  0;
rom[51384] = 12'h  0;
rom[51385] = 12'h  0;
rom[51386] = 12'h  0;
rom[51387] = 12'h  0;
rom[51388] = 12'h  0;
rom[51389] = 12'h  0;
rom[51390] = 12'h  0;
rom[51391] = 12'h  0;
rom[51392] = 12'h  0;
rom[51393] = 12'h  0;
rom[51394] = 12'h  0;
rom[51395] = 12'h  0;
rom[51396] = 12'h  0;
rom[51397] = 12'h  0;
rom[51398] = 12'h  0;
rom[51399] = 12'h  0;
rom[51400] = 12'h  0;
rom[51401] = 12'h  0;
rom[51402] = 12'h  0;
rom[51403] = 12'h  0;
rom[51404] = 12'h  0;
rom[51405] = 12'h  0;
rom[51406] = 12'h  0;
rom[51407] = 12'h  0;
rom[51408] = 12'h111;
rom[51409] = 12'h111;
rom[51410] = 12'h  0;
rom[51411] = 12'h  0;
rom[51412] = 12'h  0;
rom[51413] = 12'h111;
rom[51414] = 12'h111;
rom[51415] = 12'h111;
rom[51416] = 12'h111;
rom[51417] = 12'h  0;
rom[51418] = 12'h  0;
rom[51419] = 12'h111;
rom[51420] = 12'h222;
rom[51421] = 12'h111;
rom[51422] = 12'h111;
rom[51423] = 12'h222;
rom[51424] = 12'h333;
rom[51425] = 12'h222;
rom[51426] = 12'h222;
rom[51427] = 12'h222;
rom[51428] = 12'h222;
rom[51429] = 12'h222;
rom[51430] = 12'h111;
rom[51431] = 12'h111;
rom[51432] = 12'h111;
rom[51433] = 12'h111;
rom[51434] = 12'h111;
rom[51435] = 12'h  0;
rom[51436] = 12'h  0;
rom[51437] = 12'h  0;
rom[51438] = 12'h  0;
rom[51439] = 12'h  0;
rom[51440] = 12'h  0;
rom[51441] = 12'h  0;
rom[51442] = 12'h  0;
rom[51443] = 12'h  0;
rom[51444] = 12'h  0;
rom[51445] = 12'h  0;
rom[51446] = 12'h  0;
rom[51447] = 12'h  0;
rom[51448] = 12'h  0;
rom[51449] = 12'h  0;
rom[51450] = 12'h  0;
rom[51451] = 12'h  0;
rom[51452] = 12'h  0;
rom[51453] = 12'h  0;
rom[51454] = 12'h  0;
rom[51455] = 12'h  0;
rom[51456] = 12'h  0;
rom[51457] = 12'h  0;
rom[51458] = 12'h  0;
rom[51459] = 12'h  0;
rom[51460] = 12'h  0;
rom[51461] = 12'h  0;
rom[51462] = 12'h  0;
rom[51463] = 12'h  0;
rom[51464] = 12'h  0;
rom[51465] = 12'h  0;
rom[51466] = 12'h  0;
rom[51467] = 12'h  0;
rom[51468] = 12'h  0;
rom[51469] = 12'h  0;
rom[51470] = 12'h111;
rom[51471] = 12'h111;
rom[51472] = 12'h111;
rom[51473] = 12'h222;
rom[51474] = 12'h222;
rom[51475] = 12'h333;
rom[51476] = 12'h444;
rom[51477] = 12'h444;
rom[51478] = 12'h444;
rom[51479] = 12'h444;
rom[51480] = 12'h444;
rom[51481] = 12'h444;
rom[51482] = 12'h444;
rom[51483] = 12'h444;
rom[51484] = 12'h444;
rom[51485] = 12'h555;
rom[51486] = 12'h555;
rom[51487] = 12'h666;
rom[51488] = 12'h777;
rom[51489] = 12'h666;
rom[51490] = 12'h555;
rom[51491] = 12'h666;
rom[51492] = 12'h666;
rom[51493] = 12'h777;
rom[51494] = 12'h777;
rom[51495] = 12'h777;
rom[51496] = 12'h777;
rom[51497] = 12'h777;
rom[51498] = 12'h777;
rom[51499] = 12'h666;
rom[51500] = 12'h666;
rom[51501] = 12'h666;
rom[51502] = 12'h555;
rom[51503] = 12'h555;
rom[51504] = 12'h444;
rom[51505] = 12'h444;
rom[51506] = 12'h333;
rom[51507] = 12'h222;
rom[51508] = 12'h222;
rom[51509] = 12'h111;
rom[51510] = 12'h111;
rom[51511] = 12'h111;
rom[51512] = 12'h100;
rom[51513] = 12'h  0;
rom[51514] = 12'h  0;
rom[51515] = 12'h  0;
rom[51516] = 12'h  0;
rom[51517] = 12'h  0;
rom[51518] = 12'h  0;
rom[51519] = 12'h  0;
rom[51520] = 12'h  0;
rom[51521] = 12'h  0;
rom[51522] = 12'h  0;
rom[51523] = 12'h  0;
rom[51524] = 12'h  0;
rom[51525] = 12'h100;
rom[51526] = 12'h111;
rom[51527] = 12'h111;
rom[51528] = 12'h111;
rom[51529] = 12'h211;
rom[51530] = 12'h222;
rom[51531] = 12'h222;
rom[51532] = 12'h333;
rom[51533] = 12'h333;
rom[51534] = 12'h444;
rom[51535] = 12'h444;
rom[51536] = 12'h444;
rom[51537] = 12'h444;
rom[51538] = 12'h444;
rom[51539] = 12'h444;
rom[51540] = 12'h444;
rom[51541] = 12'h444;
rom[51542] = 12'h444;
rom[51543] = 12'h444;
rom[51544] = 12'h454;
rom[51545] = 12'h554;
rom[51546] = 12'h555;
rom[51547] = 12'h555;
rom[51548] = 12'h555;
rom[51549] = 12'h555;
rom[51550] = 12'h555;
rom[51551] = 12'h666;
rom[51552] = 12'h666;
rom[51553] = 12'h666;
rom[51554] = 12'h666;
rom[51555] = 12'h777;
rom[51556] = 12'h777;
rom[51557] = 12'h777;
rom[51558] = 12'h777;
rom[51559] = 12'h888;
rom[51560] = 12'h888;
rom[51561] = 12'h888;
rom[51562] = 12'h999;
rom[51563] = 12'h999;
rom[51564] = 12'h999;
rom[51565] = 12'haaa;
rom[51566] = 12'hbaa;
rom[51567] = 12'hbbb;
rom[51568] = 12'hbbb;
rom[51569] = 12'hbbb;
rom[51570] = 12'hccc;
rom[51571] = 12'hccc;
rom[51572] = 12'hddd;
rom[51573] = 12'hddd;
rom[51574] = 12'hddd;
rom[51575] = 12'hddd;
rom[51576] = 12'hccc;
rom[51577] = 12'hccc;
rom[51578] = 12'hccc;
rom[51579] = 12'hccc;
rom[51580] = 12'hccc;
rom[51581] = 12'hccc;
rom[51582] = 12'hccc;
rom[51583] = 12'hccc;
rom[51584] = 12'hccc;
rom[51585] = 12'hccc;
rom[51586] = 12'hccc;
rom[51587] = 12'hccc;
rom[51588] = 12'hccc;
rom[51589] = 12'hccc;
rom[51590] = 12'hccc;
rom[51591] = 12'hccc;
rom[51592] = 12'hccc;
rom[51593] = 12'hccc;
rom[51594] = 12'hccc;
rom[51595] = 12'hccc;
rom[51596] = 12'hccc;
rom[51597] = 12'hccc;
rom[51598] = 12'hccc;
rom[51599] = 12'hccc;
rom[51600] = 12'hddd;
rom[51601] = 12'hddd;
rom[51602] = 12'hccc;
rom[51603] = 12'hccc;
rom[51604] = 12'hbbb;
rom[51605] = 12'hbbb;
rom[51606] = 12'haaa;
rom[51607] = 12'haaa;
rom[51608] = 12'h999;
rom[51609] = 12'h999;
rom[51610] = 12'h999;
rom[51611] = 12'h999;
rom[51612] = 12'h999;
rom[51613] = 12'h999;
rom[51614] = 12'h999;
rom[51615] = 12'h999;
rom[51616] = 12'h999;
rom[51617] = 12'h999;
rom[51618] = 12'h999;
rom[51619] = 12'h999;
rom[51620] = 12'h999;
rom[51621] = 12'h999;
rom[51622] = 12'h999;
rom[51623] = 12'h999;
rom[51624] = 12'h999;
rom[51625] = 12'h999;
rom[51626] = 12'h999;
rom[51627] = 12'h999;
rom[51628] = 12'h999;
rom[51629] = 12'h999;
rom[51630] = 12'h999;
rom[51631] = 12'h999;
rom[51632] = 12'h999;
rom[51633] = 12'h999;
rom[51634] = 12'h999;
rom[51635] = 12'h999;
rom[51636] = 12'h999;
rom[51637] = 12'h999;
rom[51638] = 12'h999;
rom[51639] = 12'h999;
rom[51640] = 12'h999;
rom[51641] = 12'h999;
rom[51642] = 12'h999;
rom[51643] = 12'h999;
rom[51644] = 12'h999;
rom[51645] = 12'h999;
rom[51646] = 12'h999;
rom[51647] = 12'h999;
rom[51648] = 12'h999;
rom[51649] = 12'h999;
rom[51650] = 12'h999;
rom[51651] = 12'haaa;
rom[51652] = 12'haaa;
rom[51653] = 12'haaa;
rom[51654] = 12'haaa;
rom[51655] = 12'h999;
rom[51656] = 12'haaa;
rom[51657] = 12'haaa;
rom[51658] = 12'haaa;
rom[51659] = 12'haaa;
rom[51660] = 12'haaa;
rom[51661] = 12'haaa;
rom[51662] = 12'hbbb;
rom[51663] = 12'hbbb;
rom[51664] = 12'hbbb;
rom[51665] = 12'hbbb;
rom[51666] = 12'hbbb;
rom[51667] = 12'hbbb;
rom[51668] = 12'hbbb;
rom[51669] = 12'hccc;
rom[51670] = 12'hccc;
rom[51671] = 12'hccc;
rom[51672] = 12'hbbb;
rom[51673] = 12'hbbb;
rom[51674] = 12'haaa;
rom[51675] = 12'haaa;
rom[51676] = 12'haaa;
rom[51677] = 12'h999;
rom[51678] = 12'h999;
rom[51679] = 12'h888;
rom[51680] = 12'h888;
rom[51681] = 12'h888;
rom[51682] = 12'h888;
rom[51683] = 12'h888;
rom[51684] = 12'h888;
rom[51685] = 12'h777;
rom[51686] = 12'h777;
rom[51687] = 12'h777;
rom[51688] = 12'h777;
rom[51689] = 12'h777;
rom[51690] = 12'h777;
rom[51691] = 12'h777;
rom[51692] = 12'h777;
rom[51693] = 12'h777;
rom[51694] = 12'h777;
rom[51695] = 12'h777;
rom[51696] = 12'h777;
rom[51697] = 12'h777;
rom[51698] = 12'h777;
rom[51699] = 12'h777;
rom[51700] = 12'h777;
rom[51701] = 12'h777;
rom[51702] = 12'h888;
rom[51703] = 12'h888;
rom[51704] = 12'h777;
rom[51705] = 12'h777;
rom[51706] = 12'h777;
rom[51707] = 12'h777;
rom[51708] = 12'h777;
rom[51709] = 12'h666;
rom[51710] = 12'h666;
rom[51711] = 12'h666;
rom[51712] = 12'h555;
rom[51713] = 12'h444;
rom[51714] = 12'h444;
rom[51715] = 12'h444;
rom[51716] = 12'h444;
rom[51717] = 12'h444;
rom[51718] = 12'h444;
rom[51719] = 12'h444;
rom[51720] = 12'h444;
rom[51721] = 12'h333;
rom[51722] = 12'h333;
rom[51723] = 12'h333;
rom[51724] = 12'h333;
rom[51725] = 12'h222;
rom[51726] = 12'h222;
rom[51727] = 12'h111;
rom[51728] = 12'h111;
rom[51729] = 12'h111;
rom[51730] = 12'h111;
rom[51731] = 12'h111;
rom[51732] = 12'h111;
rom[51733] = 12'h111;
rom[51734] = 12'h111;
rom[51735] = 12'h111;
rom[51736] = 12'h111;
rom[51737] = 12'h111;
rom[51738] = 12'h111;
rom[51739] = 12'h111;
rom[51740] = 12'h111;
rom[51741] = 12'h111;
rom[51742] = 12'h111;
rom[51743] = 12'h111;
rom[51744] = 12'h111;
rom[51745] = 12'h111;
rom[51746] = 12'h111;
rom[51747] = 12'h111;
rom[51748] = 12'h111;
rom[51749] = 12'h111;
rom[51750] = 12'h111;
rom[51751] = 12'h111;
rom[51752] = 12'h111;
rom[51753] = 12'h111;
rom[51754] = 12'h111;
rom[51755] = 12'h111;
rom[51756] = 12'h111;
rom[51757] = 12'h111;
rom[51758] = 12'h111;
rom[51759] = 12'h111;
rom[51760] = 12'h111;
rom[51761] = 12'h111;
rom[51762] = 12'h111;
rom[51763] = 12'h111;
rom[51764] = 12'h111;
rom[51765] = 12'h111;
rom[51766] = 12'h111;
rom[51767] = 12'h111;
rom[51768] = 12'h111;
rom[51769] = 12'h111;
rom[51770] = 12'h111;
rom[51771] = 12'h111;
rom[51772] = 12'h111;
rom[51773] = 12'h111;
rom[51774] = 12'h111;
rom[51775] = 12'h111;
rom[51776] = 12'h111;
rom[51777] = 12'h111;
rom[51778] = 12'h111;
rom[51779] = 12'h  0;
rom[51780] = 12'h  0;
rom[51781] = 12'h  0;
rom[51782] = 12'h  0;
rom[51783] = 12'h  0;
rom[51784] = 12'h  0;
rom[51785] = 12'h  0;
rom[51786] = 12'h  0;
rom[51787] = 12'h  0;
rom[51788] = 12'h  0;
rom[51789] = 12'h  0;
rom[51790] = 12'h  0;
rom[51791] = 12'h  0;
rom[51792] = 12'h  0;
rom[51793] = 12'h  0;
rom[51794] = 12'h  0;
rom[51795] = 12'h  0;
rom[51796] = 12'h  0;
rom[51797] = 12'h  0;
rom[51798] = 12'h  0;
rom[51799] = 12'h  0;
rom[51800] = 12'h  0;
rom[51801] = 12'h  0;
rom[51802] = 12'h  0;
rom[51803] = 12'h  0;
rom[51804] = 12'h  0;
rom[51805] = 12'h  0;
rom[51806] = 12'h  0;
rom[51807] = 12'h  0;
rom[51808] = 12'h111;
rom[51809] = 12'h111;
rom[51810] = 12'h  0;
rom[51811] = 12'h  0;
rom[51812] = 12'h  0;
rom[51813] = 12'h111;
rom[51814] = 12'h111;
rom[51815] = 12'h111;
rom[51816] = 12'h111;
rom[51817] = 12'h  0;
rom[51818] = 12'h  0;
rom[51819] = 12'h111;
rom[51820] = 12'h111;
rom[51821] = 12'h111;
rom[51822] = 12'h111;
rom[51823] = 12'h222;
rom[51824] = 12'h333;
rom[51825] = 12'h222;
rom[51826] = 12'h222;
rom[51827] = 12'h222;
rom[51828] = 12'h222;
rom[51829] = 12'h222;
rom[51830] = 12'h111;
rom[51831] = 12'h111;
rom[51832] = 12'h111;
rom[51833] = 12'h111;
rom[51834] = 12'h111;
rom[51835] = 12'h  0;
rom[51836] = 12'h  0;
rom[51837] = 12'h  0;
rom[51838] = 12'h  0;
rom[51839] = 12'h  0;
rom[51840] = 12'h  0;
rom[51841] = 12'h  0;
rom[51842] = 12'h  0;
rom[51843] = 12'h  0;
rom[51844] = 12'h  0;
rom[51845] = 12'h  0;
rom[51846] = 12'h  0;
rom[51847] = 12'h  0;
rom[51848] = 12'h  0;
rom[51849] = 12'h  0;
rom[51850] = 12'h  0;
rom[51851] = 12'h  0;
rom[51852] = 12'h  0;
rom[51853] = 12'h  0;
rom[51854] = 12'h  0;
rom[51855] = 12'h  0;
rom[51856] = 12'h  0;
rom[51857] = 12'h  0;
rom[51858] = 12'h  0;
rom[51859] = 12'h  0;
rom[51860] = 12'h  0;
rom[51861] = 12'h  0;
rom[51862] = 12'h  0;
rom[51863] = 12'h  0;
rom[51864] = 12'h  0;
rom[51865] = 12'h  0;
rom[51866] = 12'h  0;
rom[51867] = 12'h  0;
rom[51868] = 12'h  0;
rom[51869] = 12'h  0;
rom[51870] = 12'h111;
rom[51871] = 12'h111;
rom[51872] = 12'h111;
rom[51873] = 12'h222;
rom[51874] = 12'h222;
rom[51875] = 12'h333;
rom[51876] = 12'h444;
rom[51877] = 12'h444;
rom[51878] = 12'h333;
rom[51879] = 12'h444;
rom[51880] = 12'h444;
rom[51881] = 12'h444;
rom[51882] = 12'h444;
rom[51883] = 12'h444;
rom[51884] = 12'h444;
rom[51885] = 12'h555;
rom[51886] = 12'h666;
rom[51887] = 12'h666;
rom[51888] = 12'h666;
rom[51889] = 12'h666;
rom[51890] = 12'h555;
rom[51891] = 12'h555;
rom[51892] = 12'h666;
rom[51893] = 12'h777;
rom[51894] = 12'h777;
rom[51895] = 12'h777;
rom[51896] = 12'h777;
rom[51897] = 12'h777;
rom[51898] = 12'h777;
rom[51899] = 12'h666;
rom[51900] = 12'h666;
rom[51901] = 12'h666;
rom[51902] = 12'h666;
rom[51903] = 12'h555;
rom[51904] = 12'h555;
rom[51905] = 12'h444;
rom[51906] = 12'h444;
rom[51907] = 12'h333;
rom[51908] = 12'h333;
rom[51909] = 12'h222;
rom[51910] = 12'h222;
rom[51911] = 12'h222;
rom[51912] = 12'h111;
rom[51913] = 12'h111;
rom[51914] = 12'h111;
rom[51915] = 12'h111;
rom[51916] = 12'h111;
rom[51917] = 12'h111;
rom[51918] = 12'h111;
rom[51919] = 12'h111;
rom[51920] = 12'h111;
rom[51921] = 12'h111;
rom[51922] = 12'h111;
rom[51923] = 12'h111;
rom[51924] = 12'h111;
rom[51925] = 12'h111;
rom[51926] = 12'h222;
rom[51927] = 12'h222;
rom[51928] = 12'h222;
rom[51929] = 12'h222;
rom[51930] = 12'h333;
rom[51931] = 12'h333;
rom[51932] = 12'h333;
rom[51933] = 12'h444;
rom[51934] = 12'h444;
rom[51935] = 12'h444;
rom[51936] = 12'h444;
rom[51937] = 12'h444;
rom[51938] = 12'h444;
rom[51939] = 12'h444;
rom[51940] = 12'h444;
rom[51941] = 12'h555;
rom[51942] = 12'h555;
rom[51943] = 12'h555;
rom[51944] = 12'h555;
rom[51945] = 12'h555;
rom[51946] = 12'h555;
rom[51947] = 12'h555;
rom[51948] = 12'h555;
rom[51949] = 12'h666;
rom[51950] = 12'h666;
rom[51951] = 12'h666;
rom[51952] = 12'h666;
rom[51953] = 12'h666;
rom[51954] = 12'h777;
rom[51955] = 12'h777;
rom[51956] = 12'h777;
rom[51957] = 12'h777;
rom[51958] = 12'h888;
rom[51959] = 12'h888;
rom[51960] = 12'h888;
rom[51961] = 12'h888;
rom[51962] = 12'h999;
rom[51963] = 12'h999;
rom[51964] = 12'haaa;
rom[51965] = 12'haaa;
rom[51966] = 12'hbbb;
rom[51967] = 12'hbbb;
rom[51968] = 12'hbbb;
rom[51969] = 12'hccc;
rom[51970] = 12'hccc;
rom[51971] = 12'hddd;
rom[51972] = 12'hddd;
rom[51973] = 12'hddd;
rom[51974] = 12'hddd;
rom[51975] = 12'hddd;
rom[51976] = 12'hccc;
rom[51977] = 12'hccc;
rom[51978] = 12'hccc;
rom[51979] = 12'hccc;
rom[51980] = 12'hccc;
rom[51981] = 12'hccc;
rom[51982] = 12'hccc;
rom[51983] = 12'hccc;
rom[51984] = 12'hccc;
rom[51985] = 12'hccc;
rom[51986] = 12'hccc;
rom[51987] = 12'hccc;
rom[51988] = 12'hccc;
rom[51989] = 12'hccc;
rom[51990] = 12'hddd;
rom[51991] = 12'hddd;
rom[51992] = 12'hccc;
rom[51993] = 12'hccc;
rom[51994] = 12'hccc;
rom[51995] = 12'hccc;
rom[51996] = 12'hccc;
rom[51997] = 12'hccc;
rom[51998] = 12'hccc;
rom[51999] = 12'hccc;
rom[52000] = 12'heee;
rom[52001] = 12'heee;
rom[52002] = 12'hddd;
rom[52003] = 12'hddd;
rom[52004] = 12'hccc;
rom[52005] = 12'hbbb;
rom[52006] = 12'hbbb;
rom[52007] = 12'hbbb;
rom[52008] = 12'haaa;
rom[52009] = 12'haaa;
rom[52010] = 12'haaa;
rom[52011] = 12'haaa;
rom[52012] = 12'haaa;
rom[52013] = 12'haaa;
rom[52014] = 12'haaa;
rom[52015] = 12'haaa;
rom[52016] = 12'haaa;
rom[52017] = 12'haaa;
rom[52018] = 12'haaa;
rom[52019] = 12'haaa;
rom[52020] = 12'haaa;
rom[52021] = 12'h999;
rom[52022] = 12'h999;
rom[52023] = 12'h999;
rom[52024] = 12'haaa;
rom[52025] = 12'haaa;
rom[52026] = 12'haaa;
rom[52027] = 12'haaa;
rom[52028] = 12'h999;
rom[52029] = 12'h999;
rom[52030] = 12'h999;
rom[52031] = 12'h999;
rom[52032] = 12'h999;
rom[52033] = 12'h999;
rom[52034] = 12'h999;
rom[52035] = 12'h999;
rom[52036] = 12'h999;
rom[52037] = 12'h999;
rom[52038] = 12'haaa;
rom[52039] = 12'haaa;
rom[52040] = 12'h999;
rom[52041] = 12'h999;
rom[52042] = 12'h999;
rom[52043] = 12'h999;
rom[52044] = 12'h999;
rom[52045] = 12'h999;
rom[52046] = 12'haaa;
rom[52047] = 12'haaa;
rom[52048] = 12'haaa;
rom[52049] = 12'haaa;
rom[52050] = 12'haaa;
rom[52051] = 12'haaa;
rom[52052] = 12'haaa;
rom[52053] = 12'haaa;
rom[52054] = 12'haaa;
rom[52055] = 12'haaa;
rom[52056] = 12'haaa;
rom[52057] = 12'haaa;
rom[52058] = 12'haaa;
rom[52059] = 12'haaa;
rom[52060] = 12'hbbb;
rom[52061] = 12'hbbb;
rom[52062] = 12'hbbb;
rom[52063] = 12'hbbb;
rom[52064] = 12'hbbb;
rom[52065] = 12'hbbb;
rom[52066] = 12'hccc;
rom[52067] = 12'hccc;
rom[52068] = 12'hccc;
rom[52069] = 12'hccc;
rom[52070] = 12'hccc;
rom[52071] = 12'hccc;
rom[52072] = 12'hccc;
rom[52073] = 12'hbbb;
rom[52074] = 12'hbbb;
rom[52075] = 12'haaa;
rom[52076] = 12'haaa;
rom[52077] = 12'haaa;
rom[52078] = 12'h999;
rom[52079] = 12'h999;
rom[52080] = 12'h999;
rom[52081] = 12'h888;
rom[52082] = 12'h888;
rom[52083] = 12'h888;
rom[52084] = 12'h888;
rom[52085] = 12'h888;
rom[52086] = 12'h888;
rom[52087] = 12'h888;
rom[52088] = 12'h777;
rom[52089] = 12'h777;
rom[52090] = 12'h777;
rom[52091] = 12'h777;
rom[52092] = 12'h777;
rom[52093] = 12'h777;
rom[52094] = 12'h777;
rom[52095] = 12'h777;
rom[52096] = 12'h777;
rom[52097] = 12'h777;
rom[52098] = 12'h777;
rom[52099] = 12'h777;
rom[52100] = 12'h777;
rom[52101] = 12'h777;
rom[52102] = 12'h777;
rom[52103] = 12'h888;
rom[52104] = 12'h888;
rom[52105] = 12'h888;
rom[52106] = 12'h888;
rom[52107] = 12'h888;
rom[52108] = 12'h777;
rom[52109] = 12'h777;
rom[52110] = 12'h777;
rom[52111] = 12'h666;
rom[52112] = 12'h666;
rom[52113] = 12'h555;
rom[52114] = 12'h555;
rom[52115] = 12'h444;
rom[52116] = 12'h444;
rom[52117] = 12'h444;
rom[52118] = 12'h444;
rom[52119] = 12'h444;
rom[52120] = 12'h444;
rom[52121] = 12'h444;
rom[52122] = 12'h444;
rom[52123] = 12'h444;
rom[52124] = 12'h444;
rom[52125] = 12'h333;
rom[52126] = 12'h222;
rom[52127] = 12'h111;
rom[52128] = 12'h222;
rom[52129] = 12'h222;
rom[52130] = 12'h111;
rom[52131] = 12'h111;
rom[52132] = 12'h111;
rom[52133] = 12'h111;
rom[52134] = 12'h111;
rom[52135] = 12'h111;
rom[52136] = 12'h111;
rom[52137] = 12'h111;
rom[52138] = 12'h111;
rom[52139] = 12'h111;
rom[52140] = 12'h111;
rom[52141] = 12'h111;
rom[52142] = 12'h111;
rom[52143] = 12'h111;
rom[52144] = 12'h111;
rom[52145] = 12'h111;
rom[52146] = 12'h111;
rom[52147] = 12'h111;
rom[52148] = 12'h111;
rom[52149] = 12'h111;
rom[52150] = 12'h111;
rom[52151] = 12'h111;
rom[52152] = 12'h111;
rom[52153] = 12'h111;
rom[52154] = 12'h111;
rom[52155] = 12'h111;
rom[52156] = 12'h111;
rom[52157] = 12'h111;
rom[52158] = 12'h111;
rom[52159] = 12'h111;
rom[52160] = 12'h111;
rom[52161] = 12'h111;
rom[52162] = 12'h111;
rom[52163] = 12'h222;
rom[52164] = 12'h222;
rom[52165] = 12'h222;
rom[52166] = 12'h222;
rom[52167] = 12'h222;
rom[52168] = 12'h111;
rom[52169] = 12'h111;
rom[52170] = 12'h111;
rom[52171] = 12'h111;
rom[52172] = 12'h111;
rom[52173] = 12'h111;
rom[52174] = 12'h111;
rom[52175] = 12'h111;
rom[52176] = 12'h111;
rom[52177] = 12'h111;
rom[52178] = 12'h  0;
rom[52179] = 12'h  0;
rom[52180] = 12'h  0;
rom[52181] = 12'h  0;
rom[52182] = 12'h  0;
rom[52183] = 12'h  0;
rom[52184] = 12'h  0;
rom[52185] = 12'h  0;
rom[52186] = 12'h  0;
rom[52187] = 12'h  0;
rom[52188] = 12'h  0;
rom[52189] = 12'h  0;
rom[52190] = 12'h  0;
rom[52191] = 12'h  0;
rom[52192] = 12'h  0;
rom[52193] = 12'h  0;
rom[52194] = 12'h  0;
rom[52195] = 12'h  0;
rom[52196] = 12'h  0;
rom[52197] = 12'h  0;
rom[52198] = 12'h  0;
rom[52199] = 12'h  0;
rom[52200] = 12'h  0;
rom[52201] = 12'h  0;
rom[52202] = 12'h  0;
rom[52203] = 12'h  0;
rom[52204] = 12'h  0;
rom[52205] = 12'h  0;
rom[52206] = 12'h  0;
rom[52207] = 12'h  0;
rom[52208] = 12'h111;
rom[52209] = 12'h111;
rom[52210] = 12'h  0;
rom[52211] = 12'h  0;
rom[52212] = 12'h  0;
rom[52213] = 12'h111;
rom[52214] = 12'h111;
rom[52215] = 12'h111;
rom[52216] = 12'h111;
rom[52217] = 12'h  0;
rom[52218] = 12'h111;
rom[52219] = 12'h111;
rom[52220] = 12'h111;
rom[52221] = 12'h111;
rom[52222] = 12'h222;
rom[52223] = 12'h222;
rom[52224] = 12'h333;
rom[52225] = 12'h222;
rom[52226] = 12'h222;
rom[52227] = 12'h222;
rom[52228] = 12'h111;
rom[52229] = 12'h111;
rom[52230] = 12'h111;
rom[52231] = 12'h111;
rom[52232] = 12'h111;
rom[52233] = 12'h111;
rom[52234] = 12'h111;
rom[52235] = 12'h  0;
rom[52236] = 12'h  0;
rom[52237] = 12'h  0;
rom[52238] = 12'h  0;
rom[52239] = 12'h  0;
rom[52240] = 12'h  0;
rom[52241] = 12'h  0;
rom[52242] = 12'h  0;
rom[52243] = 12'h  0;
rom[52244] = 12'h  0;
rom[52245] = 12'h  0;
rom[52246] = 12'h  0;
rom[52247] = 12'h  0;
rom[52248] = 12'h  0;
rom[52249] = 12'h  0;
rom[52250] = 12'h  0;
rom[52251] = 12'h  0;
rom[52252] = 12'h  0;
rom[52253] = 12'h  0;
rom[52254] = 12'h  0;
rom[52255] = 12'h  0;
rom[52256] = 12'h  0;
rom[52257] = 12'h  0;
rom[52258] = 12'h  0;
rom[52259] = 12'h  0;
rom[52260] = 12'h  0;
rom[52261] = 12'h  0;
rom[52262] = 12'h  0;
rom[52263] = 12'h  0;
rom[52264] = 12'h  0;
rom[52265] = 12'h  0;
rom[52266] = 12'h  0;
rom[52267] = 12'h  0;
rom[52268] = 12'h  0;
rom[52269] = 12'h  0;
rom[52270] = 12'h111;
rom[52271] = 12'h111;
rom[52272] = 12'h111;
rom[52273] = 12'h222;
rom[52274] = 12'h222;
rom[52275] = 12'h333;
rom[52276] = 12'h444;
rom[52277] = 12'h444;
rom[52278] = 12'h333;
rom[52279] = 12'h444;
rom[52280] = 12'h444;
rom[52281] = 12'h444;
rom[52282] = 12'h444;
rom[52283] = 12'h444;
rom[52284] = 12'h444;
rom[52285] = 12'h555;
rom[52286] = 12'h666;
rom[52287] = 12'h777;
rom[52288] = 12'h666;
rom[52289] = 12'h555;
rom[52290] = 12'h555;
rom[52291] = 12'h555;
rom[52292] = 12'h666;
rom[52293] = 12'h666;
rom[52294] = 12'h666;
rom[52295] = 12'h777;
rom[52296] = 12'h777;
rom[52297] = 12'h777;
rom[52298] = 12'h777;
rom[52299] = 12'h777;
rom[52300] = 12'h666;
rom[52301] = 12'h666;
rom[52302] = 12'h666;
rom[52303] = 12'h666;
rom[52304] = 12'h666;
rom[52305] = 12'h555;
rom[52306] = 12'h555;
rom[52307] = 12'h444;
rom[52308] = 12'h444;
rom[52309] = 12'h333;
rom[52310] = 12'h333;
rom[52311] = 12'h333;
rom[52312] = 12'h333;
rom[52313] = 12'h222;
rom[52314] = 12'h222;
rom[52315] = 12'h222;
rom[52316] = 12'h222;
rom[52317] = 12'h222;
rom[52318] = 12'h222;
rom[52319] = 12'h222;
rom[52320] = 12'h222;
rom[52321] = 12'h222;
rom[52322] = 12'h222;
rom[52323] = 12'h222;
rom[52324] = 12'h333;
rom[52325] = 12'h333;
rom[52326] = 12'h333;
rom[52327] = 12'h333;
rom[52328] = 12'h333;
rom[52329] = 12'h444;
rom[52330] = 12'h444;
rom[52331] = 12'h444;
rom[52332] = 12'h444;
rom[52333] = 12'h444;
rom[52334] = 12'h444;
rom[52335] = 12'h444;
rom[52336] = 12'h555;
rom[52337] = 12'h555;
rom[52338] = 12'h555;
rom[52339] = 12'h555;
rom[52340] = 12'h555;
rom[52341] = 12'h555;
rom[52342] = 12'h555;
rom[52343] = 12'h555;
rom[52344] = 12'h555;
rom[52345] = 12'h555;
rom[52346] = 12'h555;
rom[52347] = 12'h666;
rom[52348] = 12'h666;
rom[52349] = 12'h666;
rom[52350] = 12'h666;
rom[52351] = 12'h666;
rom[52352] = 12'h666;
rom[52353] = 12'h777;
rom[52354] = 12'h777;
rom[52355] = 12'h777;
rom[52356] = 12'h777;
rom[52357] = 12'h888;
rom[52358] = 12'h888;
rom[52359] = 12'h888;
rom[52360] = 12'h999;
rom[52361] = 12'h999;
rom[52362] = 12'h999;
rom[52363] = 12'haaa;
rom[52364] = 12'haaa;
rom[52365] = 12'haaa;
rom[52366] = 12'hbbb;
rom[52367] = 12'hbbb;
rom[52368] = 12'hccc;
rom[52369] = 12'hccc;
rom[52370] = 12'hddd;
rom[52371] = 12'hddd;
rom[52372] = 12'hddd;
rom[52373] = 12'hddd;
rom[52374] = 12'hddd;
rom[52375] = 12'hccc;
rom[52376] = 12'hccc;
rom[52377] = 12'hccc;
rom[52378] = 12'hccc;
rom[52379] = 12'hccc;
rom[52380] = 12'hccc;
rom[52381] = 12'hddd;
rom[52382] = 12'hddd;
rom[52383] = 12'hccc;
rom[52384] = 12'hddd;
rom[52385] = 12'hddd;
rom[52386] = 12'hddd;
rom[52387] = 12'hddd;
rom[52388] = 12'hddd;
rom[52389] = 12'hddd;
rom[52390] = 12'hddd;
rom[52391] = 12'hddd;
rom[52392] = 12'hddd;
rom[52393] = 12'hddd;
rom[52394] = 12'hddd;
rom[52395] = 12'hccc;
rom[52396] = 12'hccc;
rom[52397] = 12'hddd;
rom[52398] = 12'hddd;
rom[52399] = 12'hddd;
rom[52400] = 12'hfff;
rom[52401] = 12'hfff;
rom[52402] = 12'heee;
rom[52403] = 12'heee;
rom[52404] = 12'hddd;
rom[52405] = 12'hccc;
rom[52406] = 12'hccc;
rom[52407] = 12'hbbb;
rom[52408] = 12'hbbb;
rom[52409] = 12'hbbb;
rom[52410] = 12'hbbb;
rom[52411] = 12'hbbb;
rom[52412] = 12'hbbb;
rom[52413] = 12'hbbb;
rom[52414] = 12'hbbb;
rom[52415] = 12'hbbb;
rom[52416] = 12'hbbb;
rom[52417] = 12'hbbb;
rom[52418] = 12'haaa;
rom[52419] = 12'haaa;
rom[52420] = 12'haaa;
rom[52421] = 12'haaa;
rom[52422] = 12'haaa;
rom[52423] = 12'haaa;
rom[52424] = 12'haaa;
rom[52425] = 12'haaa;
rom[52426] = 12'haaa;
rom[52427] = 12'haaa;
rom[52428] = 12'haaa;
rom[52429] = 12'haaa;
rom[52430] = 12'haaa;
rom[52431] = 12'haaa;
rom[52432] = 12'h999;
rom[52433] = 12'h999;
rom[52434] = 12'h999;
rom[52435] = 12'h999;
rom[52436] = 12'h999;
rom[52437] = 12'haaa;
rom[52438] = 12'haaa;
rom[52439] = 12'haaa;
rom[52440] = 12'haaa;
rom[52441] = 12'haaa;
rom[52442] = 12'haaa;
rom[52443] = 12'haaa;
rom[52444] = 12'haaa;
rom[52445] = 12'haaa;
rom[52446] = 12'haaa;
rom[52447] = 12'haaa;
rom[52448] = 12'haaa;
rom[52449] = 12'haaa;
rom[52450] = 12'haaa;
rom[52451] = 12'haaa;
rom[52452] = 12'haaa;
rom[52453] = 12'haaa;
rom[52454] = 12'haaa;
rom[52455] = 12'haaa;
rom[52456] = 12'haaa;
rom[52457] = 12'haaa;
rom[52458] = 12'haaa;
rom[52459] = 12'hbbb;
rom[52460] = 12'hbbb;
rom[52461] = 12'hbbb;
rom[52462] = 12'hbbb;
rom[52463] = 12'hbbb;
rom[52464] = 12'hbbb;
rom[52465] = 12'hccc;
rom[52466] = 12'hccc;
rom[52467] = 12'hccc;
rom[52468] = 12'hccc;
rom[52469] = 12'hccc;
rom[52470] = 12'hccc;
rom[52471] = 12'hccc;
rom[52472] = 12'hccc;
rom[52473] = 12'hccc;
rom[52474] = 12'hbbb;
rom[52475] = 12'hbbb;
rom[52476] = 12'haaa;
rom[52477] = 12'haaa;
rom[52478] = 12'h999;
rom[52479] = 12'h999;
rom[52480] = 12'h999;
rom[52481] = 12'h999;
rom[52482] = 12'h888;
rom[52483] = 12'h888;
rom[52484] = 12'h888;
rom[52485] = 12'h888;
rom[52486] = 12'h888;
rom[52487] = 12'h888;
rom[52488] = 12'h777;
rom[52489] = 12'h777;
rom[52490] = 12'h777;
rom[52491] = 12'h777;
rom[52492] = 12'h777;
rom[52493] = 12'h777;
rom[52494] = 12'h777;
rom[52495] = 12'h777;
rom[52496] = 12'h777;
rom[52497] = 12'h777;
rom[52498] = 12'h777;
rom[52499] = 12'h777;
rom[52500] = 12'h777;
rom[52501] = 12'h777;
rom[52502] = 12'h777;
rom[52503] = 12'h777;
rom[52504] = 12'h888;
rom[52505] = 12'h888;
rom[52506] = 12'h999;
rom[52507] = 12'h999;
rom[52508] = 12'h999;
rom[52509] = 12'h888;
rom[52510] = 12'h777;
rom[52511] = 12'h777;
rom[52512] = 12'h777;
rom[52513] = 12'h666;
rom[52514] = 12'h666;
rom[52515] = 12'h555;
rom[52516] = 12'h555;
rom[52517] = 12'h555;
rom[52518] = 12'h444;
rom[52519] = 12'h444;
rom[52520] = 12'h555;
rom[52521] = 12'h444;
rom[52522] = 12'h444;
rom[52523] = 12'h444;
rom[52524] = 12'h444;
rom[52525] = 12'h333;
rom[52526] = 12'h333;
rom[52527] = 12'h333;
rom[52528] = 12'h222;
rom[52529] = 12'h222;
rom[52530] = 12'h222;
rom[52531] = 12'h111;
rom[52532] = 12'h111;
rom[52533] = 12'h111;
rom[52534] = 12'h111;
rom[52535] = 12'h111;
rom[52536] = 12'h111;
rom[52537] = 12'h111;
rom[52538] = 12'h111;
rom[52539] = 12'h111;
rom[52540] = 12'h111;
rom[52541] = 12'h111;
rom[52542] = 12'h111;
rom[52543] = 12'h111;
rom[52544] = 12'h111;
rom[52545] = 12'h111;
rom[52546] = 12'h111;
rom[52547] = 12'h111;
rom[52548] = 12'h111;
rom[52549] = 12'h111;
rom[52550] = 12'h111;
rom[52551] = 12'h111;
rom[52552] = 12'h111;
rom[52553] = 12'h111;
rom[52554] = 12'h111;
rom[52555] = 12'h111;
rom[52556] = 12'h111;
rom[52557] = 12'h111;
rom[52558] = 12'h111;
rom[52559] = 12'h111;
rom[52560] = 12'h222;
rom[52561] = 12'h222;
rom[52562] = 12'h222;
rom[52563] = 12'h222;
rom[52564] = 12'h222;
rom[52565] = 12'h222;
rom[52566] = 12'h222;
rom[52567] = 12'h222;
rom[52568] = 12'h111;
rom[52569] = 12'h111;
rom[52570] = 12'h111;
rom[52571] = 12'h111;
rom[52572] = 12'h111;
rom[52573] = 12'h111;
rom[52574] = 12'h111;
rom[52575] = 12'h111;
rom[52576] = 12'h111;
rom[52577] = 12'h  0;
rom[52578] = 12'h  0;
rom[52579] = 12'h  0;
rom[52580] = 12'h  0;
rom[52581] = 12'h  0;
rom[52582] = 12'h  0;
rom[52583] = 12'h  0;
rom[52584] = 12'h  0;
rom[52585] = 12'h  0;
rom[52586] = 12'h  0;
rom[52587] = 12'h  0;
rom[52588] = 12'h  0;
rom[52589] = 12'h  0;
rom[52590] = 12'h  0;
rom[52591] = 12'h  0;
rom[52592] = 12'h  0;
rom[52593] = 12'h  0;
rom[52594] = 12'h  0;
rom[52595] = 12'h  0;
rom[52596] = 12'h  0;
rom[52597] = 12'h  0;
rom[52598] = 12'h  0;
rom[52599] = 12'h  0;
rom[52600] = 12'h  0;
rom[52601] = 12'h  0;
rom[52602] = 12'h  0;
rom[52603] = 12'h  0;
rom[52604] = 12'h  0;
rom[52605] = 12'h  0;
rom[52606] = 12'h  0;
rom[52607] = 12'h  0;
rom[52608] = 12'h111;
rom[52609] = 12'h111;
rom[52610] = 12'h  0;
rom[52611] = 12'h  0;
rom[52612] = 12'h  0;
rom[52613] = 12'h111;
rom[52614] = 12'h111;
rom[52615] = 12'h111;
rom[52616] = 12'h  0;
rom[52617] = 12'h  0;
rom[52618] = 12'h111;
rom[52619] = 12'h111;
rom[52620] = 12'h111;
rom[52621] = 12'h111;
rom[52622] = 12'h222;
rom[52623] = 12'h333;
rom[52624] = 12'h333;
rom[52625] = 12'h222;
rom[52626] = 12'h222;
rom[52627] = 12'h111;
rom[52628] = 12'h111;
rom[52629] = 12'h111;
rom[52630] = 12'h111;
rom[52631] = 12'h111;
rom[52632] = 12'h111;
rom[52633] = 12'h111;
rom[52634] = 12'h  0;
rom[52635] = 12'h  0;
rom[52636] = 12'h  0;
rom[52637] = 12'h  0;
rom[52638] = 12'h  0;
rom[52639] = 12'h  0;
rom[52640] = 12'h  0;
rom[52641] = 12'h  0;
rom[52642] = 12'h  0;
rom[52643] = 12'h  0;
rom[52644] = 12'h  0;
rom[52645] = 12'h  0;
rom[52646] = 12'h  0;
rom[52647] = 12'h  0;
rom[52648] = 12'h  0;
rom[52649] = 12'h  0;
rom[52650] = 12'h  0;
rom[52651] = 12'h  0;
rom[52652] = 12'h  0;
rom[52653] = 12'h  0;
rom[52654] = 12'h  0;
rom[52655] = 12'h  0;
rom[52656] = 12'h  0;
rom[52657] = 12'h  0;
rom[52658] = 12'h  0;
rom[52659] = 12'h  0;
rom[52660] = 12'h  0;
rom[52661] = 12'h  0;
rom[52662] = 12'h  0;
rom[52663] = 12'h  0;
rom[52664] = 12'h  0;
rom[52665] = 12'h  0;
rom[52666] = 12'h  0;
rom[52667] = 12'h  0;
rom[52668] = 12'h  0;
rom[52669] = 12'h  0;
rom[52670] = 12'h  0;
rom[52671] = 12'h111;
rom[52672] = 12'h111;
rom[52673] = 12'h111;
rom[52674] = 12'h222;
rom[52675] = 12'h222;
rom[52676] = 12'h333;
rom[52677] = 12'h333;
rom[52678] = 12'h333;
rom[52679] = 12'h444;
rom[52680] = 12'h444;
rom[52681] = 12'h444;
rom[52682] = 12'h444;
rom[52683] = 12'h444;
rom[52684] = 12'h444;
rom[52685] = 12'h555;
rom[52686] = 12'h666;
rom[52687] = 12'h666;
rom[52688] = 12'h555;
rom[52689] = 12'h555;
rom[52690] = 12'h444;
rom[52691] = 12'h555;
rom[52692] = 12'h666;
rom[52693] = 12'h666;
rom[52694] = 12'h666;
rom[52695] = 12'h666;
rom[52696] = 12'h777;
rom[52697] = 12'h777;
rom[52698] = 12'h777;
rom[52699] = 12'h777;
rom[52700] = 12'h777;
rom[52701] = 12'h777;
rom[52702] = 12'h666;
rom[52703] = 12'h666;
rom[52704] = 12'h666;
rom[52705] = 12'h666;
rom[52706] = 12'h555;
rom[52707] = 12'h555;
rom[52708] = 12'h555;
rom[52709] = 12'h555;
rom[52710] = 12'h444;
rom[52711] = 12'h444;
rom[52712] = 12'h444;
rom[52713] = 12'h444;
rom[52714] = 12'h333;
rom[52715] = 12'h333;
rom[52716] = 12'h333;
rom[52717] = 12'h333;
rom[52718] = 12'h333;
rom[52719] = 12'h333;
rom[52720] = 12'h333;
rom[52721] = 12'h333;
rom[52722] = 12'h333;
rom[52723] = 12'h444;
rom[52724] = 12'h444;
rom[52725] = 12'h444;
rom[52726] = 12'h444;
rom[52727] = 12'h444;
rom[52728] = 12'h444;
rom[52729] = 12'h444;
rom[52730] = 12'h444;
rom[52731] = 12'h444;
rom[52732] = 12'h444;
rom[52733] = 12'h555;
rom[52734] = 12'h555;
rom[52735] = 12'h555;
rom[52736] = 12'h555;
rom[52737] = 12'h555;
rom[52738] = 12'h555;
rom[52739] = 12'h555;
rom[52740] = 12'h555;
rom[52741] = 12'h555;
rom[52742] = 12'h555;
rom[52743] = 12'h555;
rom[52744] = 12'h555;
rom[52745] = 12'h555;
rom[52746] = 12'h555;
rom[52747] = 12'h666;
rom[52748] = 12'h666;
rom[52749] = 12'h666;
rom[52750] = 12'h666;
rom[52751] = 12'h666;
rom[52752] = 12'h777;
rom[52753] = 12'h777;
rom[52754] = 12'h777;
rom[52755] = 12'h777;
rom[52756] = 12'h888;
rom[52757] = 12'h888;
rom[52758] = 12'h888;
rom[52759] = 12'h888;
rom[52760] = 12'h999;
rom[52761] = 12'h999;
rom[52762] = 12'haaa;
rom[52763] = 12'haaa;
rom[52764] = 12'haaa;
rom[52765] = 12'hbbb;
rom[52766] = 12'hbbb;
rom[52767] = 12'hccc;
rom[52768] = 12'hddd;
rom[52769] = 12'hddd;
rom[52770] = 12'hddd;
rom[52771] = 12'hddd;
rom[52772] = 12'hddd;
rom[52773] = 12'hddd;
rom[52774] = 12'hccc;
rom[52775] = 12'hccc;
rom[52776] = 12'hccc;
rom[52777] = 12'hccc;
rom[52778] = 12'hccc;
rom[52779] = 12'hccc;
rom[52780] = 12'hddd;
rom[52781] = 12'hddd;
rom[52782] = 12'hddd;
rom[52783] = 12'hddd;
rom[52784] = 12'hddd;
rom[52785] = 12'hddd;
rom[52786] = 12'hddd;
rom[52787] = 12'hddd;
rom[52788] = 12'hddd;
rom[52789] = 12'hddd;
rom[52790] = 12'hddd;
rom[52791] = 12'hddd;
rom[52792] = 12'hddd;
rom[52793] = 12'hddd;
rom[52794] = 12'hddd;
rom[52795] = 12'hddd;
rom[52796] = 12'hddd;
rom[52797] = 12'hddd;
rom[52798] = 12'hddd;
rom[52799] = 12'hddd;
rom[52800] = 12'hfff;
rom[52801] = 12'hfff;
rom[52802] = 12'hfff;
rom[52803] = 12'heee;
rom[52804] = 12'heee;
rom[52805] = 12'hddd;
rom[52806] = 12'hddd;
rom[52807] = 12'hccc;
rom[52808] = 12'hccc;
rom[52809] = 12'hccc;
rom[52810] = 12'hccc;
rom[52811] = 12'hbbb;
rom[52812] = 12'hbbb;
rom[52813] = 12'hbbb;
rom[52814] = 12'hbbb;
rom[52815] = 12'hbbb;
rom[52816] = 12'hbbb;
rom[52817] = 12'hbbb;
rom[52818] = 12'hbbb;
rom[52819] = 12'haaa;
rom[52820] = 12'haaa;
rom[52821] = 12'haaa;
rom[52822] = 12'haaa;
rom[52823] = 12'hbbb;
rom[52824] = 12'haaa;
rom[52825] = 12'haaa;
rom[52826] = 12'haaa;
rom[52827] = 12'haaa;
rom[52828] = 12'haaa;
rom[52829] = 12'haaa;
rom[52830] = 12'haaa;
rom[52831] = 12'haaa;
rom[52832] = 12'haaa;
rom[52833] = 12'haaa;
rom[52834] = 12'haaa;
rom[52835] = 12'haaa;
rom[52836] = 12'haaa;
rom[52837] = 12'haaa;
rom[52838] = 12'haaa;
rom[52839] = 12'haaa;
rom[52840] = 12'haaa;
rom[52841] = 12'haaa;
rom[52842] = 12'haaa;
rom[52843] = 12'haaa;
rom[52844] = 12'haaa;
rom[52845] = 12'haaa;
rom[52846] = 12'haaa;
rom[52847] = 12'haaa;
rom[52848] = 12'haaa;
rom[52849] = 12'haaa;
rom[52850] = 12'haaa;
rom[52851] = 12'haaa;
rom[52852] = 12'haaa;
rom[52853] = 12'haaa;
rom[52854] = 12'haaa;
rom[52855] = 12'haaa;
rom[52856] = 12'haaa;
rom[52857] = 12'haaa;
rom[52858] = 12'hbbb;
rom[52859] = 12'hbbb;
rom[52860] = 12'hbbb;
rom[52861] = 12'hbbb;
rom[52862] = 12'hccc;
rom[52863] = 12'hccc;
rom[52864] = 12'hccc;
rom[52865] = 12'hccc;
rom[52866] = 12'hccc;
rom[52867] = 12'hccc;
rom[52868] = 12'hccc;
rom[52869] = 12'hccc;
rom[52870] = 12'hccc;
rom[52871] = 12'hccc;
rom[52872] = 12'hccc;
rom[52873] = 12'hccc;
rom[52874] = 12'hbbb;
rom[52875] = 12'hbbb;
rom[52876] = 12'hbbb;
rom[52877] = 12'haaa;
rom[52878] = 12'haaa;
rom[52879] = 12'haaa;
rom[52880] = 12'h999;
rom[52881] = 12'h999;
rom[52882] = 12'h999;
rom[52883] = 12'h888;
rom[52884] = 12'h888;
rom[52885] = 12'h888;
rom[52886] = 12'h888;
rom[52887] = 12'h888;
rom[52888] = 12'h888;
rom[52889] = 12'h888;
rom[52890] = 12'h888;
rom[52891] = 12'h888;
rom[52892] = 12'h888;
rom[52893] = 12'h888;
rom[52894] = 12'h888;
rom[52895] = 12'h777;
rom[52896] = 12'h777;
rom[52897] = 12'h777;
rom[52898] = 12'h777;
rom[52899] = 12'h777;
rom[52900] = 12'h777;
rom[52901] = 12'h777;
rom[52902] = 12'h777;
rom[52903] = 12'h777;
rom[52904] = 12'h777;
rom[52905] = 12'h888;
rom[52906] = 12'h999;
rom[52907] = 12'h999;
rom[52908] = 12'h999;
rom[52909] = 12'h999;
rom[52910] = 12'h888;
rom[52911] = 12'h888;
rom[52912] = 12'h888;
rom[52913] = 12'h777;
rom[52914] = 12'h666;
rom[52915] = 12'h666;
rom[52916] = 12'h555;
rom[52917] = 12'h555;
rom[52918] = 12'h555;
rom[52919] = 12'h555;
rom[52920] = 12'h555;
rom[52921] = 12'h555;
rom[52922] = 12'h444;
rom[52923] = 12'h444;
rom[52924] = 12'h444;
rom[52925] = 12'h444;
rom[52926] = 12'h444;
rom[52927] = 12'h333;
rom[52928] = 12'h222;
rom[52929] = 12'h222;
rom[52930] = 12'h222;
rom[52931] = 12'h222;
rom[52932] = 12'h222;
rom[52933] = 12'h222;
rom[52934] = 12'h111;
rom[52935] = 12'h111;
rom[52936] = 12'h222;
rom[52937] = 12'h222;
rom[52938] = 12'h222;
rom[52939] = 12'h222;
rom[52940] = 12'h111;
rom[52941] = 12'h111;
rom[52942] = 12'h111;
rom[52943] = 12'h111;
rom[52944] = 12'h111;
rom[52945] = 12'h111;
rom[52946] = 12'h111;
rom[52947] = 12'h111;
rom[52948] = 12'h111;
rom[52949] = 12'h111;
rom[52950] = 12'h111;
rom[52951] = 12'h111;
rom[52952] = 12'h111;
rom[52953] = 12'h111;
rom[52954] = 12'h111;
rom[52955] = 12'h111;
rom[52956] = 12'h111;
rom[52957] = 12'h111;
rom[52958] = 12'h111;
rom[52959] = 12'h111;
rom[52960] = 12'h222;
rom[52961] = 12'h222;
rom[52962] = 12'h222;
rom[52963] = 12'h222;
rom[52964] = 12'h222;
rom[52965] = 12'h222;
rom[52966] = 12'h222;
rom[52967] = 12'h222;
rom[52968] = 12'h111;
rom[52969] = 12'h111;
rom[52970] = 12'h111;
rom[52971] = 12'h111;
rom[52972] = 12'h111;
rom[52973] = 12'h111;
rom[52974] = 12'h111;
rom[52975] = 12'h111;
rom[52976] = 12'h111;
rom[52977] = 12'h  0;
rom[52978] = 12'h  0;
rom[52979] = 12'h  0;
rom[52980] = 12'h  0;
rom[52981] = 12'h  0;
rom[52982] = 12'h  0;
rom[52983] = 12'h  0;
rom[52984] = 12'h  0;
rom[52985] = 12'h  0;
rom[52986] = 12'h  0;
rom[52987] = 12'h  0;
rom[52988] = 12'h  0;
rom[52989] = 12'h  0;
rom[52990] = 12'h  0;
rom[52991] = 12'h  0;
rom[52992] = 12'h  0;
rom[52993] = 12'h  0;
rom[52994] = 12'h  0;
rom[52995] = 12'h  0;
rom[52996] = 12'h  0;
rom[52997] = 12'h  0;
rom[52998] = 12'h  0;
rom[52999] = 12'h  0;
rom[53000] = 12'h  0;
rom[53001] = 12'h  0;
rom[53002] = 12'h  0;
rom[53003] = 12'h  0;
rom[53004] = 12'h  0;
rom[53005] = 12'h  0;
rom[53006] = 12'h  0;
rom[53007] = 12'h  0;
rom[53008] = 12'h111;
rom[53009] = 12'h  0;
rom[53010] = 12'h  0;
rom[53011] = 12'h  0;
rom[53012] = 12'h  0;
rom[53013] = 12'h111;
rom[53014] = 12'h111;
rom[53015] = 12'h  0;
rom[53016] = 12'h  0;
rom[53017] = 12'h  0;
rom[53018] = 12'h111;
rom[53019] = 12'h111;
rom[53020] = 12'h111;
rom[53021] = 12'h111;
rom[53022] = 12'h222;
rom[53023] = 12'h333;
rom[53024] = 12'h222;
rom[53025] = 12'h222;
rom[53026] = 12'h222;
rom[53027] = 12'h111;
rom[53028] = 12'h111;
rom[53029] = 12'h111;
rom[53030] = 12'h111;
rom[53031] = 12'h111;
rom[53032] = 12'h111;
rom[53033] = 12'h  0;
rom[53034] = 12'h  0;
rom[53035] = 12'h  0;
rom[53036] = 12'h  0;
rom[53037] = 12'h  0;
rom[53038] = 12'h  0;
rom[53039] = 12'h  0;
rom[53040] = 12'h  0;
rom[53041] = 12'h  0;
rom[53042] = 12'h  0;
rom[53043] = 12'h  0;
rom[53044] = 12'h  0;
rom[53045] = 12'h  0;
rom[53046] = 12'h  0;
rom[53047] = 12'h  0;
rom[53048] = 12'h  0;
rom[53049] = 12'h  0;
rom[53050] = 12'h  0;
rom[53051] = 12'h  0;
rom[53052] = 12'h  0;
rom[53053] = 12'h  0;
rom[53054] = 12'h  0;
rom[53055] = 12'h  0;
rom[53056] = 12'h  0;
rom[53057] = 12'h  0;
rom[53058] = 12'h  0;
rom[53059] = 12'h  0;
rom[53060] = 12'h  0;
rom[53061] = 12'h  0;
rom[53062] = 12'h  0;
rom[53063] = 12'h  0;
rom[53064] = 12'h  0;
rom[53065] = 12'h  0;
rom[53066] = 12'h  0;
rom[53067] = 12'h  0;
rom[53068] = 12'h  0;
rom[53069] = 12'h  0;
rom[53070] = 12'h  0;
rom[53071] = 12'h111;
rom[53072] = 12'h111;
rom[53073] = 12'h111;
rom[53074] = 12'h222;
rom[53075] = 12'h222;
rom[53076] = 12'h333;
rom[53077] = 12'h333;
rom[53078] = 12'h333;
rom[53079] = 12'h444;
rom[53080] = 12'h444;
rom[53081] = 12'h444;
rom[53082] = 12'h333;
rom[53083] = 12'h444;
rom[53084] = 12'h444;
rom[53085] = 12'h555;
rom[53086] = 12'h666;
rom[53087] = 12'h666;
rom[53088] = 12'h555;
rom[53089] = 12'h555;
rom[53090] = 12'h444;
rom[53091] = 12'h555;
rom[53092] = 12'h666;
rom[53093] = 12'h666;
rom[53094] = 12'h666;
rom[53095] = 12'h666;
rom[53096] = 12'h777;
rom[53097] = 12'h777;
rom[53098] = 12'h666;
rom[53099] = 12'h666;
rom[53100] = 12'h666;
rom[53101] = 12'h666;
rom[53102] = 12'h666;
rom[53103] = 12'h666;
rom[53104] = 12'h666;
rom[53105] = 12'h666;
rom[53106] = 12'h666;
rom[53107] = 12'h555;
rom[53108] = 12'h555;
rom[53109] = 12'h555;
rom[53110] = 12'h555;
rom[53111] = 12'h555;
rom[53112] = 12'h555;
rom[53113] = 12'h555;
rom[53114] = 12'h444;
rom[53115] = 12'h444;
rom[53116] = 12'h444;
rom[53117] = 12'h444;
rom[53118] = 12'h444;
rom[53119] = 12'h444;
rom[53120] = 12'h444;
rom[53121] = 12'h444;
rom[53122] = 12'h444;
rom[53123] = 12'h444;
rom[53124] = 12'h444;
rom[53125] = 12'h444;
rom[53126] = 12'h444;
rom[53127] = 12'h444;
rom[53128] = 12'h444;
rom[53129] = 12'h444;
rom[53130] = 12'h555;
rom[53131] = 12'h555;
rom[53132] = 12'h555;
rom[53133] = 12'h555;
rom[53134] = 12'h555;
rom[53135] = 12'h555;
rom[53136] = 12'h555;
rom[53137] = 12'h555;
rom[53138] = 12'h555;
rom[53139] = 12'h555;
rom[53140] = 12'h555;
rom[53141] = 12'h555;
rom[53142] = 12'h555;
rom[53143] = 12'h555;
rom[53144] = 12'h666;
rom[53145] = 12'h666;
rom[53146] = 12'h666;
rom[53147] = 12'h666;
rom[53148] = 12'h666;
rom[53149] = 12'h666;
rom[53150] = 12'h666;
rom[53151] = 12'h777;
rom[53152] = 12'h777;
rom[53153] = 12'h777;
rom[53154] = 12'h777;
rom[53155] = 12'h888;
rom[53156] = 12'h888;
rom[53157] = 12'h888;
rom[53158] = 12'h999;
rom[53159] = 12'h999;
rom[53160] = 12'haaa;
rom[53161] = 12'haaa;
rom[53162] = 12'haaa;
rom[53163] = 12'hbbb;
rom[53164] = 12'hbbb;
rom[53165] = 12'hbbb;
rom[53166] = 12'hccc;
rom[53167] = 12'hccc;
rom[53168] = 12'hddd;
rom[53169] = 12'hddd;
rom[53170] = 12'hddd;
rom[53171] = 12'hddd;
rom[53172] = 12'hddd;
rom[53173] = 12'hddd;
rom[53174] = 12'hccc;
rom[53175] = 12'hccc;
rom[53176] = 12'hccc;
rom[53177] = 12'hccc;
rom[53178] = 12'hccc;
rom[53179] = 12'hddd;
rom[53180] = 12'hddd;
rom[53181] = 12'hddd;
rom[53182] = 12'hddd;
rom[53183] = 12'hddd;
rom[53184] = 12'hddd;
rom[53185] = 12'hddd;
rom[53186] = 12'hddd;
rom[53187] = 12'hddd;
rom[53188] = 12'hddd;
rom[53189] = 12'hddd;
rom[53190] = 12'hddd;
rom[53191] = 12'hddd;
rom[53192] = 12'hddd;
rom[53193] = 12'hddd;
rom[53194] = 12'hddd;
rom[53195] = 12'hddd;
rom[53196] = 12'hddd;
rom[53197] = 12'heee;
rom[53198] = 12'heee;
rom[53199] = 12'heee;
rom[53200] = 12'hfff;
rom[53201] = 12'hfff;
rom[53202] = 12'hfff;
rom[53203] = 12'hfff;
rom[53204] = 12'hfff;
rom[53205] = 12'heee;
rom[53206] = 12'heee;
rom[53207] = 12'hddd;
rom[53208] = 12'hddd;
rom[53209] = 12'hddd;
rom[53210] = 12'hccc;
rom[53211] = 12'hccc;
rom[53212] = 12'hccc;
rom[53213] = 12'hccc;
rom[53214] = 12'hbbb;
rom[53215] = 12'hbbb;
rom[53216] = 12'hbbb;
rom[53217] = 12'hbbb;
rom[53218] = 12'hbbb;
rom[53219] = 12'hbbb;
rom[53220] = 12'hbbb;
rom[53221] = 12'hbbb;
rom[53222] = 12'hbbb;
rom[53223] = 12'hbbb;
rom[53224] = 12'hbbb;
rom[53225] = 12'hbbb;
rom[53226] = 12'hbbb;
rom[53227] = 12'haaa;
rom[53228] = 12'haaa;
rom[53229] = 12'haaa;
rom[53230] = 12'haaa;
rom[53231] = 12'haaa;
rom[53232] = 12'hbbb;
rom[53233] = 12'hbbb;
rom[53234] = 12'haaa;
rom[53235] = 12'haaa;
rom[53236] = 12'hbbb;
rom[53237] = 12'hbbb;
rom[53238] = 12'hbbb;
rom[53239] = 12'hbbb;
rom[53240] = 12'hbbb;
rom[53241] = 12'hbbb;
rom[53242] = 12'hbbb;
rom[53243] = 12'hbbb;
rom[53244] = 12'hbbb;
rom[53245] = 12'hbbb;
rom[53246] = 12'hbbb;
rom[53247] = 12'hbbb;
rom[53248] = 12'haaa;
rom[53249] = 12'haaa;
rom[53250] = 12'haaa;
rom[53251] = 12'haaa;
rom[53252] = 12'haaa;
rom[53253] = 12'haaa;
rom[53254] = 12'haaa;
rom[53255] = 12'haaa;
rom[53256] = 12'hbbb;
rom[53257] = 12'hbbb;
rom[53258] = 12'hbbb;
rom[53259] = 12'hbbb;
rom[53260] = 12'hbbb;
rom[53261] = 12'hccc;
rom[53262] = 12'hccc;
rom[53263] = 12'hccc;
rom[53264] = 12'hccc;
rom[53265] = 12'hccc;
rom[53266] = 12'hccc;
rom[53267] = 12'hccc;
rom[53268] = 12'hccc;
rom[53269] = 12'hccc;
rom[53270] = 12'hddd;
rom[53271] = 12'hddd;
rom[53272] = 12'hddd;
rom[53273] = 12'hccc;
rom[53274] = 12'hccc;
rom[53275] = 12'hccc;
rom[53276] = 12'hbbb;
rom[53277] = 12'hbbb;
rom[53278] = 12'haaa;
rom[53279] = 12'haaa;
rom[53280] = 12'haaa;
rom[53281] = 12'h999;
rom[53282] = 12'h999;
rom[53283] = 12'h999;
rom[53284] = 12'h999;
rom[53285] = 12'h999;
rom[53286] = 12'h888;
rom[53287] = 12'h888;
rom[53288] = 12'h888;
rom[53289] = 12'h888;
rom[53290] = 12'h888;
rom[53291] = 12'h888;
rom[53292] = 12'h888;
rom[53293] = 12'h888;
rom[53294] = 12'h888;
rom[53295] = 12'h888;
rom[53296] = 12'h777;
rom[53297] = 12'h777;
rom[53298] = 12'h777;
rom[53299] = 12'h777;
rom[53300] = 12'h777;
rom[53301] = 12'h777;
rom[53302] = 12'h777;
rom[53303] = 12'h777;
rom[53304] = 12'h777;
rom[53305] = 12'h888;
rom[53306] = 12'h888;
rom[53307] = 12'h888;
rom[53308] = 12'h999;
rom[53309] = 12'h999;
rom[53310] = 12'haaa;
rom[53311] = 12'haaa;
rom[53312] = 12'h999;
rom[53313] = 12'h999;
rom[53314] = 12'h888;
rom[53315] = 12'h777;
rom[53316] = 12'h666;
rom[53317] = 12'h555;
rom[53318] = 12'h555;
rom[53319] = 12'h444;
rom[53320] = 12'h555;
rom[53321] = 12'h555;
rom[53322] = 12'h555;
rom[53323] = 12'h555;
rom[53324] = 12'h555;
rom[53325] = 12'h444;
rom[53326] = 12'h444;
rom[53327] = 12'h444;
rom[53328] = 12'h333;
rom[53329] = 12'h333;
rom[53330] = 12'h333;
rom[53331] = 12'h222;
rom[53332] = 12'h222;
rom[53333] = 12'h222;
rom[53334] = 12'h222;
rom[53335] = 12'h222;
rom[53336] = 12'h222;
rom[53337] = 12'h222;
rom[53338] = 12'h222;
rom[53339] = 12'h222;
rom[53340] = 12'h222;
rom[53341] = 12'h222;
rom[53342] = 12'h111;
rom[53343] = 12'h111;
rom[53344] = 12'h222;
rom[53345] = 12'h111;
rom[53346] = 12'h111;
rom[53347] = 12'h111;
rom[53348] = 12'h111;
rom[53349] = 12'h111;
rom[53350] = 12'h111;
rom[53351] = 12'h111;
rom[53352] = 12'h111;
rom[53353] = 12'h111;
rom[53354] = 12'h111;
rom[53355] = 12'h111;
rom[53356] = 12'h111;
rom[53357] = 12'h111;
rom[53358] = 12'h222;
rom[53359] = 12'h222;
rom[53360] = 12'h222;
rom[53361] = 12'h222;
rom[53362] = 12'h111;
rom[53363] = 12'h111;
rom[53364] = 12'h111;
rom[53365] = 12'h111;
rom[53366] = 12'h111;
rom[53367] = 12'h111;
rom[53368] = 12'h111;
rom[53369] = 12'h111;
rom[53370] = 12'h111;
rom[53371] = 12'h111;
rom[53372] = 12'h111;
rom[53373] = 12'h111;
rom[53374] = 12'h111;
rom[53375] = 12'h111;
rom[53376] = 12'h111;
rom[53377] = 12'h  0;
rom[53378] = 12'h  0;
rom[53379] = 12'h  0;
rom[53380] = 12'h  0;
rom[53381] = 12'h  0;
rom[53382] = 12'h  0;
rom[53383] = 12'h  0;
rom[53384] = 12'h  0;
rom[53385] = 12'h  0;
rom[53386] = 12'h  0;
rom[53387] = 12'h  0;
rom[53388] = 12'h  0;
rom[53389] = 12'h  0;
rom[53390] = 12'h  0;
rom[53391] = 12'h  0;
rom[53392] = 12'h  0;
rom[53393] = 12'h  0;
rom[53394] = 12'h  0;
rom[53395] = 12'h  0;
rom[53396] = 12'h  0;
rom[53397] = 12'h  0;
rom[53398] = 12'h  0;
rom[53399] = 12'h  0;
rom[53400] = 12'h  0;
rom[53401] = 12'h  0;
rom[53402] = 12'h  0;
rom[53403] = 12'h  0;
rom[53404] = 12'h  0;
rom[53405] = 12'h  0;
rom[53406] = 12'h111;
rom[53407] = 12'h111;
rom[53408] = 12'h111;
rom[53409] = 12'h  0;
rom[53410] = 12'h  0;
rom[53411] = 12'h  0;
rom[53412] = 12'h111;
rom[53413] = 12'h111;
rom[53414] = 12'h111;
rom[53415] = 12'h  0;
rom[53416] = 12'h  0;
rom[53417] = 12'h  0;
rom[53418] = 12'h111;
rom[53419] = 12'h111;
rom[53420] = 12'h111;
rom[53421] = 12'h222;
rom[53422] = 12'h222;
rom[53423] = 12'h333;
rom[53424] = 12'h222;
rom[53425] = 12'h222;
rom[53426] = 12'h111;
rom[53427] = 12'h111;
rom[53428] = 12'h111;
rom[53429] = 12'h111;
rom[53430] = 12'h111;
rom[53431] = 12'h111;
rom[53432] = 12'h  0;
rom[53433] = 12'h  0;
rom[53434] = 12'h  0;
rom[53435] = 12'h  0;
rom[53436] = 12'h  0;
rom[53437] = 12'h  0;
rom[53438] = 12'h  0;
rom[53439] = 12'h  0;
rom[53440] = 12'h  0;
rom[53441] = 12'h  0;
rom[53442] = 12'h  0;
rom[53443] = 12'h  0;
rom[53444] = 12'h  0;
rom[53445] = 12'h  0;
rom[53446] = 12'h  0;
rom[53447] = 12'h  0;
rom[53448] = 12'h  0;
rom[53449] = 12'h  0;
rom[53450] = 12'h  0;
rom[53451] = 12'h  0;
rom[53452] = 12'h  0;
rom[53453] = 12'h  0;
rom[53454] = 12'h  0;
rom[53455] = 12'h  0;
rom[53456] = 12'h  0;
rom[53457] = 12'h  0;
rom[53458] = 12'h  0;
rom[53459] = 12'h  0;
rom[53460] = 12'h  0;
rom[53461] = 12'h  0;
rom[53462] = 12'h  0;
rom[53463] = 12'h  0;
rom[53464] = 12'h  0;
rom[53465] = 12'h  0;
rom[53466] = 12'h  0;
rom[53467] = 12'h  0;
rom[53468] = 12'h  0;
rom[53469] = 12'h  0;
rom[53470] = 12'h  0;
rom[53471] = 12'h  0;
rom[53472] = 12'h111;
rom[53473] = 12'h111;
rom[53474] = 12'h222;
rom[53475] = 12'h222;
rom[53476] = 12'h333;
rom[53477] = 12'h333;
rom[53478] = 12'h333;
rom[53479] = 12'h333;
rom[53480] = 12'h444;
rom[53481] = 12'h333;
rom[53482] = 12'h333;
rom[53483] = 12'h333;
rom[53484] = 12'h444;
rom[53485] = 12'h555;
rom[53486] = 12'h666;
rom[53487] = 12'h666;
rom[53488] = 12'h555;
rom[53489] = 12'h444;
rom[53490] = 12'h444;
rom[53491] = 12'h555;
rom[53492] = 12'h555;
rom[53493] = 12'h666;
rom[53494] = 12'h666;
rom[53495] = 12'h666;
rom[53496] = 12'h777;
rom[53497] = 12'h777;
rom[53498] = 12'h666;
rom[53499] = 12'h666;
rom[53500] = 12'h666;
rom[53501] = 12'h666;
rom[53502] = 12'h666;
rom[53503] = 12'h666;
rom[53504] = 12'h666;
rom[53505] = 12'h666;
rom[53506] = 12'h666;
rom[53507] = 12'h666;
rom[53508] = 12'h666;
rom[53509] = 12'h666;
rom[53510] = 12'h666;
rom[53511] = 12'h666;
rom[53512] = 12'h555;
rom[53513] = 12'h555;
rom[53514] = 12'h555;
rom[53515] = 12'h555;
rom[53516] = 12'h555;
rom[53517] = 12'h555;
rom[53518] = 12'h555;
rom[53519] = 12'h555;
rom[53520] = 12'h555;
rom[53521] = 12'h555;
rom[53522] = 12'h555;
rom[53523] = 12'h555;
rom[53524] = 12'h555;
rom[53525] = 12'h555;
rom[53526] = 12'h555;
rom[53527] = 12'h555;
rom[53528] = 12'h444;
rom[53529] = 12'h555;
rom[53530] = 12'h555;
rom[53531] = 12'h555;
rom[53532] = 12'h555;
rom[53533] = 12'h555;
rom[53534] = 12'h555;
rom[53535] = 12'h555;
rom[53536] = 12'h555;
rom[53537] = 12'h555;
rom[53538] = 12'h555;
rom[53539] = 12'h555;
rom[53540] = 12'h555;
rom[53541] = 12'h555;
rom[53542] = 12'h555;
rom[53543] = 12'h666;
rom[53544] = 12'h666;
rom[53545] = 12'h666;
rom[53546] = 12'h666;
rom[53547] = 12'h666;
rom[53548] = 12'h666;
rom[53549] = 12'h777;
rom[53550] = 12'h777;
rom[53551] = 12'h777;
rom[53552] = 12'h777;
rom[53553] = 12'h888;
rom[53554] = 12'h888;
rom[53555] = 12'h888;
rom[53556] = 12'h888;
rom[53557] = 12'h999;
rom[53558] = 12'h999;
rom[53559] = 12'h999;
rom[53560] = 12'haaa;
rom[53561] = 12'haaa;
rom[53562] = 12'hbbb;
rom[53563] = 12'hbbb;
rom[53564] = 12'hbbb;
rom[53565] = 12'hccc;
rom[53566] = 12'hccc;
rom[53567] = 12'hddd;
rom[53568] = 12'hddd;
rom[53569] = 12'hddd;
rom[53570] = 12'hddd;
rom[53571] = 12'hddd;
rom[53572] = 12'hddd;
rom[53573] = 12'hccc;
rom[53574] = 12'hccc;
rom[53575] = 12'hccc;
rom[53576] = 12'hccc;
rom[53577] = 12'hccc;
rom[53578] = 12'hccc;
rom[53579] = 12'hddd;
rom[53580] = 12'hddd;
rom[53581] = 12'hddd;
rom[53582] = 12'hddd;
rom[53583] = 12'hccc;
rom[53584] = 12'hddd;
rom[53585] = 12'hddd;
rom[53586] = 12'hddd;
rom[53587] = 12'hddd;
rom[53588] = 12'hddd;
rom[53589] = 12'hddd;
rom[53590] = 12'hddd;
rom[53591] = 12'hddd;
rom[53592] = 12'hddd;
rom[53593] = 12'hddd;
rom[53594] = 12'hddd;
rom[53595] = 12'hddd;
rom[53596] = 12'hddd;
rom[53597] = 12'heee;
rom[53598] = 12'heee;
rom[53599] = 12'heee;
rom[53600] = 12'hfff;
rom[53601] = 12'hfff;
rom[53602] = 12'hfff;
rom[53603] = 12'hfff;
rom[53604] = 12'hfff;
rom[53605] = 12'hfff;
rom[53606] = 12'hfff;
rom[53607] = 12'heee;
rom[53608] = 12'heee;
rom[53609] = 12'hddd;
rom[53610] = 12'hddd;
rom[53611] = 12'hddd;
rom[53612] = 12'hccc;
rom[53613] = 12'hccc;
rom[53614] = 12'hccc;
rom[53615] = 12'hbbb;
rom[53616] = 12'hbbb;
rom[53617] = 12'hbbb;
rom[53618] = 12'hbbb;
rom[53619] = 12'hbbb;
rom[53620] = 12'hbbb;
rom[53621] = 12'hbbb;
rom[53622] = 12'hbbb;
rom[53623] = 12'hbbb;
rom[53624] = 12'hbbb;
rom[53625] = 12'hbbb;
rom[53626] = 12'hbbb;
rom[53627] = 12'hbbb;
rom[53628] = 12'hbbb;
rom[53629] = 12'hbbb;
rom[53630] = 12'hbbb;
rom[53631] = 12'hbbb;
rom[53632] = 12'hbbb;
rom[53633] = 12'hbbb;
rom[53634] = 12'hbbb;
rom[53635] = 12'hbbb;
rom[53636] = 12'hbbb;
rom[53637] = 12'hbbb;
rom[53638] = 12'hbbb;
rom[53639] = 12'hbbb;
rom[53640] = 12'hbbb;
rom[53641] = 12'hbbb;
rom[53642] = 12'hbbb;
rom[53643] = 12'hbbb;
rom[53644] = 12'hbbb;
rom[53645] = 12'hbbb;
rom[53646] = 12'hbbb;
rom[53647] = 12'hbbb;
rom[53648] = 12'hbbb;
rom[53649] = 12'hbbb;
rom[53650] = 12'hbbb;
rom[53651] = 12'hbbb;
rom[53652] = 12'hbbb;
rom[53653] = 12'hbbb;
rom[53654] = 12'hbbb;
rom[53655] = 12'hbbb;
rom[53656] = 12'hbbb;
rom[53657] = 12'hbbb;
rom[53658] = 12'hbbb;
rom[53659] = 12'hccc;
rom[53660] = 12'hccc;
rom[53661] = 12'hccc;
rom[53662] = 12'hccc;
rom[53663] = 12'hccc;
rom[53664] = 12'hccc;
rom[53665] = 12'hccc;
rom[53666] = 12'hddd;
rom[53667] = 12'hddd;
rom[53668] = 12'hccc;
rom[53669] = 12'hddd;
rom[53670] = 12'hddd;
rom[53671] = 12'hddd;
rom[53672] = 12'hddd;
rom[53673] = 12'hddd;
rom[53674] = 12'hccc;
rom[53675] = 12'hccc;
rom[53676] = 12'hccc;
rom[53677] = 12'hccc;
rom[53678] = 12'hbbb;
rom[53679] = 12'hbbb;
rom[53680] = 12'haaa;
rom[53681] = 12'haaa;
rom[53682] = 12'haaa;
rom[53683] = 12'h999;
rom[53684] = 12'h999;
rom[53685] = 12'h999;
rom[53686] = 12'h999;
rom[53687] = 12'h999;
rom[53688] = 12'h999;
rom[53689] = 12'h999;
rom[53690] = 12'h999;
rom[53691] = 12'h999;
rom[53692] = 12'h999;
rom[53693] = 12'h999;
rom[53694] = 12'h999;
rom[53695] = 12'h888;
rom[53696] = 12'h888;
rom[53697] = 12'h888;
rom[53698] = 12'h888;
rom[53699] = 12'h888;
rom[53700] = 12'h777;
rom[53701] = 12'h777;
rom[53702] = 12'h777;
rom[53703] = 12'h777;
rom[53704] = 12'h777;
rom[53705] = 12'h888;
rom[53706] = 12'h888;
rom[53707] = 12'h888;
rom[53708] = 12'h888;
rom[53709] = 12'h888;
rom[53710] = 12'h999;
rom[53711] = 12'haaa;
rom[53712] = 12'haaa;
rom[53713] = 12'haaa;
rom[53714] = 12'haaa;
rom[53715] = 12'h999;
rom[53716] = 12'h888;
rom[53717] = 12'h777;
rom[53718] = 12'h666;
rom[53719] = 12'h555;
rom[53720] = 12'h555;
rom[53721] = 12'h555;
rom[53722] = 12'h555;
rom[53723] = 12'h555;
rom[53724] = 12'h555;
rom[53725] = 12'h555;
rom[53726] = 12'h444;
rom[53727] = 12'h444;
rom[53728] = 12'h444;
rom[53729] = 12'h444;
rom[53730] = 12'h333;
rom[53731] = 12'h333;
rom[53732] = 12'h333;
rom[53733] = 12'h222;
rom[53734] = 12'h222;
rom[53735] = 12'h222;
rom[53736] = 12'h222;
rom[53737] = 12'h222;
rom[53738] = 12'h222;
rom[53739] = 12'h222;
rom[53740] = 12'h222;
rom[53741] = 12'h222;
rom[53742] = 12'h222;
rom[53743] = 12'h222;
rom[53744] = 12'h222;
rom[53745] = 12'h111;
rom[53746] = 12'h111;
rom[53747] = 12'h111;
rom[53748] = 12'h111;
rom[53749] = 12'h111;
rom[53750] = 12'h111;
rom[53751] = 12'h111;
rom[53752] = 12'h111;
rom[53753] = 12'h111;
rom[53754] = 12'h111;
rom[53755] = 12'h222;
rom[53756] = 12'h222;
rom[53757] = 12'h222;
rom[53758] = 12'h222;
rom[53759] = 12'h222;
rom[53760] = 12'h222;
rom[53761] = 12'h111;
rom[53762] = 12'h111;
rom[53763] = 12'h111;
rom[53764] = 12'h111;
rom[53765] = 12'h111;
rom[53766] = 12'h111;
rom[53767] = 12'h111;
rom[53768] = 12'h111;
rom[53769] = 12'h111;
rom[53770] = 12'h111;
rom[53771] = 12'h111;
rom[53772] = 12'h111;
rom[53773] = 12'h111;
rom[53774] = 12'h111;
rom[53775] = 12'h111;
rom[53776] = 12'h111;
rom[53777] = 12'h  0;
rom[53778] = 12'h  0;
rom[53779] = 12'h  0;
rom[53780] = 12'h  0;
rom[53781] = 12'h  0;
rom[53782] = 12'h  0;
rom[53783] = 12'h  0;
rom[53784] = 12'h  0;
rom[53785] = 12'h  0;
rom[53786] = 12'h  0;
rom[53787] = 12'h  0;
rom[53788] = 12'h  0;
rom[53789] = 12'h  0;
rom[53790] = 12'h  0;
rom[53791] = 12'h  0;
rom[53792] = 12'h  0;
rom[53793] = 12'h  0;
rom[53794] = 12'h  0;
rom[53795] = 12'h  0;
rom[53796] = 12'h  0;
rom[53797] = 12'h  0;
rom[53798] = 12'h  0;
rom[53799] = 12'h  0;
rom[53800] = 12'h  0;
rom[53801] = 12'h  0;
rom[53802] = 12'h  0;
rom[53803] = 12'h  0;
rom[53804] = 12'h  0;
rom[53805] = 12'h  0;
rom[53806] = 12'h111;
rom[53807] = 12'h111;
rom[53808] = 12'h111;
rom[53809] = 12'h  0;
rom[53810] = 12'h  0;
rom[53811] = 12'h  0;
rom[53812] = 12'h111;
rom[53813] = 12'h111;
rom[53814] = 12'h111;
rom[53815] = 12'h  0;
rom[53816] = 12'h  0;
rom[53817] = 12'h  0;
rom[53818] = 12'h111;
rom[53819] = 12'h111;
rom[53820] = 12'h111;
rom[53821] = 12'h222;
rom[53822] = 12'h333;
rom[53823] = 12'h333;
rom[53824] = 12'h222;
rom[53825] = 12'h222;
rom[53826] = 12'h111;
rom[53827] = 12'h111;
rom[53828] = 12'h111;
rom[53829] = 12'h111;
rom[53830] = 12'h111;
rom[53831] = 12'h  0;
rom[53832] = 12'h  0;
rom[53833] = 12'h  0;
rom[53834] = 12'h  0;
rom[53835] = 12'h  0;
rom[53836] = 12'h  0;
rom[53837] = 12'h  0;
rom[53838] = 12'h  0;
rom[53839] = 12'h  0;
rom[53840] = 12'h  0;
rom[53841] = 12'h  0;
rom[53842] = 12'h  0;
rom[53843] = 12'h  0;
rom[53844] = 12'h  0;
rom[53845] = 12'h  0;
rom[53846] = 12'h  0;
rom[53847] = 12'h  0;
rom[53848] = 12'h  0;
rom[53849] = 12'h  0;
rom[53850] = 12'h  0;
rom[53851] = 12'h  0;
rom[53852] = 12'h  0;
rom[53853] = 12'h  0;
rom[53854] = 12'h  0;
rom[53855] = 12'h  0;
rom[53856] = 12'h  0;
rom[53857] = 12'h  0;
rom[53858] = 12'h  0;
rom[53859] = 12'h  0;
rom[53860] = 12'h  0;
rom[53861] = 12'h  0;
rom[53862] = 12'h  0;
rom[53863] = 12'h  0;
rom[53864] = 12'h  0;
rom[53865] = 12'h  0;
rom[53866] = 12'h  0;
rom[53867] = 12'h  0;
rom[53868] = 12'h  0;
rom[53869] = 12'h  0;
rom[53870] = 12'h  0;
rom[53871] = 12'h  0;
rom[53872] = 12'h111;
rom[53873] = 12'h111;
rom[53874] = 12'h222;
rom[53875] = 12'h222;
rom[53876] = 12'h333;
rom[53877] = 12'h333;
rom[53878] = 12'h222;
rom[53879] = 12'h333;
rom[53880] = 12'h333;
rom[53881] = 12'h333;
rom[53882] = 12'h333;
rom[53883] = 12'h333;
rom[53884] = 12'h444;
rom[53885] = 12'h555;
rom[53886] = 12'h555;
rom[53887] = 12'h555;
rom[53888] = 12'h444;
rom[53889] = 12'h444;
rom[53890] = 12'h444;
rom[53891] = 12'h444;
rom[53892] = 12'h555;
rom[53893] = 12'h555;
rom[53894] = 12'h666;
rom[53895] = 12'h666;
rom[53896] = 12'h777;
rom[53897] = 12'h777;
rom[53898] = 12'h666;
rom[53899] = 12'h666;
rom[53900] = 12'h666;
rom[53901] = 12'h666;
rom[53902] = 12'h666;
rom[53903] = 12'h666;
rom[53904] = 12'h666;
rom[53905] = 12'h666;
rom[53906] = 12'h666;
rom[53907] = 12'h666;
rom[53908] = 12'h666;
rom[53909] = 12'h666;
rom[53910] = 12'h666;
rom[53911] = 12'h666;
rom[53912] = 12'h666;
rom[53913] = 12'h666;
rom[53914] = 12'h555;
rom[53915] = 12'h555;
rom[53916] = 12'h555;
rom[53917] = 12'h555;
rom[53918] = 12'h666;
rom[53919] = 12'h666;
rom[53920] = 12'h555;
rom[53921] = 12'h555;
rom[53922] = 12'h555;
rom[53923] = 12'h555;
rom[53924] = 12'h555;
rom[53925] = 12'h555;
rom[53926] = 12'h555;
rom[53927] = 12'h555;
rom[53928] = 12'h555;
rom[53929] = 12'h555;
rom[53930] = 12'h555;
rom[53931] = 12'h555;
rom[53932] = 12'h555;
rom[53933] = 12'h555;
rom[53934] = 12'h555;
rom[53935] = 12'h555;
rom[53936] = 12'h555;
rom[53937] = 12'h555;
rom[53938] = 12'h555;
rom[53939] = 12'h666;
rom[53940] = 12'h666;
rom[53941] = 12'h666;
rom[53942] = 12'h666;
rom[53943] = 12'h666;
rom[53944] = 12'h666;
rom[53945] = 12'h666;
rom[53946] = 12'h666;
rom[53947] = 12'h777;
rom[53948] = 12'h777;
rom[53949] = 12'h777;
rom[53950] = 12'h777;
rom[53951] = 12'h777;
rom[53952] = 12'h888;
rom[53953] = 12'h888;
rom[53954] = 12'h888;
rom[53955] = 12'h999;
rom[53956] = 12'h999;
rom[53957] = 12'h999;
rom[53958] = 12'haaa;
rom[53959] = 12'haaa;
rom[53960] = 12'haaa;
rom[53961] = 12'haaa;
rom[53962] = 12'hbbb;
rom[53963] = 12'hbbb;
rom[53964] = 12'hbbb;
rom[53965] = 12'hccc;
rom[53966] = 12'hddd;
rom[53967] = 12'hddd;
rom[53968] = 12'hddd;
rom[53969] = 12'hddd;
rom[53970] = 12'hddd;
rom[53971] = 12'hddd;
rom[53972] = 12'hddd;
rom[53973] = 12'hccc;
rom[53974] = 12'hccc;
rom[53975] = 12'hccc;
rom[53976] = 12'hccc;
rom[53977] = 12'hccc;
rom[53978] = 12'hccc;
rom[53979] = 12'hccc;
rom[53980] = 12'hccc;
rom[53981] = 12'hccc;
rom[53982] = 12'hccc;
rom[53983] = 12'hccc;
rom[53984] = 12'hccc;
rom[53985] = 12'hccc;
rom[53986] = 12'hccc;
rom[53987] = 12'hccc;
rom[53988] = 12'hccc;
rom[53989] = 12'hccc;
rom[53990] = 12'hccc;
rom[53991] = 12'hccc;
rom[53992] = 12'hccc;
rom[53993] = 12'hccc;
rom[53994] = 12'hccc;
rom[53995] = 12'hddd;
rom[53996] = 12'hddd;
rom[53997] = 12'hddd;
rom[53998] = 12'hddd;
rom[53999] = 12'hddd;
rom[54000] = 12'hfff;
rom[54001] = 12'hfff;
rom[54002] = 12'hfff;
rom[54003] = 12'hfff;
rom[54004] = 12'hfff;
rom[54005] = 12'hfff;
rom[54006] = 12'hfff;
rom[54007] = 12'hfff;
rom[54008] = 12'hfff;
rom[54009] = 12'heee;
rom[54010] = 12'heee;
rom[54011] = 12'hddd;
rom[54012] = 12'hddd;
rom[54013] = 12'hccc;
rom[54014] = 12'hccc;
rom[54015] = 12'hccc;
rom[54016] = 12'hccc;
rom[54017] = 12'hccc;
rom[54018] = 12'hccc;
rom[54019] = 12'hbbb;
rom[54020] = 12'hbbb;
rom[54021] = 12'hbbb;
rom[54022] = 12'hbbb;
rom[54023] = 12'hbbb;
rom[54024] = 12'hccc;
rom[54025] = 12'hccc;
rom[54026] = 12'hbbb;
rom[54027] = 12'hbbb;
rom[54028] = 12'hbbb;
rom[54029] = 12'hbbb;
rom[54030] = 12'hccc;
rom[54031] = 12'hccc;
rom[54032] = 12'hbbb;
rom[54033] = 12'hbbb;
rom[54034] = 12'hbbb;
rom[54035] = 12'hccc;
rom[54036] = 12'hccc;
rom[54037] = 12'hccc;
rom[54038] = 12'hccc;
rom[54039] = 12'hccc;
rom[54040] = 12'hbbb;
rom[54041] = 12'hbbb;
rom[54042] = 12'hbbb;
rom[54043] = 12'hbbb;
rom[54044] = 12'hbbb;
rom[54045] = 12'hbbb;
rom[54046] = 12'hbbb;
rom[54047] = 12'hbbb;
rom[54048] = 12'hbbb;
rom[54049] = 12'hbbb;
rom[54050] = 12'hbbb;
rom[54051] = 12'hbbb;
rom[54052] = 12'hbbb;
rom[54053] = 12'hbbb;
rom[54054] = 12'hbbb;
rom[54055] = 12'hbbb;
rom[54056] = 12'hbbb;
rom[54057] = 12'hccc;
rom[54058] = 12'hccc;
rom[54059] = 12'hccc;
rom[54060] = 12'hccc;
rom[54061] = 12'hccc;
rom[54062] = 12'hccc;
rom[54063] = 12'hccc;
rom[54064] = 12'hddd;
rom[54065] = 12'hddd;
rom[54066] = 12'hddd;
rom[54067] = 12'hddd;
rom[54068] = 12'hddd;
rom[54069] = 12'hddd;
rom[54070] = 12'hddd;
rom[54071] = 12'hddd;
rom[54072] = 12'hddd;
rom[54073] = 12'hddd;
rom[54074] = 12'hddd;
rom[54075] = 12'hccc;
rom[54076] = 12'hccc;
rom[54077] = 12'hccc;
rom[54078] = 12'hccc;
rom[54079] = 12'hbbb;
rom[54080] = 12'haaa;
rom[54081] = 12'haaa;
rom[54082] = 12'haaa;
rom[54083] = 12'haaa;
rom[54084] = 12'haaa;
rom[54085] = 12'haaa;
rom[54086] = 12'haaa;
rom[54087] = 12'h999;
rom[54088] = 12'h999;
rom[54089] = 12'h999;
rom[54090] = 12'h999;
rom[54091] = 12'h999;
rom[54092] = 12'h999;
rom[54093] = 12'h999;
rom[54094] = 12'h999;
rom[54095] = 12'h999;
rom[54096] = 12'h999;
rom[54097] = 12'h999;
rom[54098] = 12'h999;
rom[54099] = 12'h888;
rom[54100] = 12'h888;
rom[54101] = 12'h777;
rom[54102] = 12'h777;
rom[54103] = 12'h777;
rom[54104] = 12'h777;
rom[54105] = 12'h888;
rom[54106] = 12'h888;
rom[54107] = 12'h888;
rom[54108] = 12'h777;
rom[54109] = 12'h777;
rom[54110] = 12'h888;
rom[54111] = 12'h888;
rom[54112] = 12'haaa;
rom[54113] = 12'haaa;
rom[54114] = 12'hbbb;
rom[54115] = 12'haaa;
rom[54116] = 12'haaa;
rom[54117] = 12'h999;
rom[54118] = 12'h888;
rom[54119] = 12'h888;
rom[54120] = 12'h555;
rom[54121] = 12'h555;
rom[54122] = 12'h555;
rom[54123] = 12'h555;
rom[54124] = 12'h555;
rom[54125] = 12'h555;
rom[54126] = 12'h444;
rom[54127] = 12'h444;
rom[54128] = 12'h555;
rom[54129] = 12'h555;
rom[54130] = 12'h444;
rom[54131] = 12'h444;
rom[54132] = 12'h333;
rom[54133] = 12'h333;
rom[54134] = 12'h333;
rom[54135] = 12'h222;
rom[54136] = 12'h222;
rom[54137] = 12'h222;
rom[54138] = 12'h222;
rom[54139] = 12'h222;
rom[54140] = 12'h222;
rom[54141] = 12'h222;
rom[54142] = 12'h222;
rom[54143] = 12'h222;
rom[54144] = 12'h222;
rom[54145] = 12'h111;
rom[54146] = 12'h111;
rom[54147] = 12'h111;
rom[54148] = 12'h111;
rom[54149] = 12'h111;
rom[54150] = 12'h111;
rom[54151] = 12'h111;
rom[54152] = 12'h111;
rom[54153] = 12'h111;
rom[54154] = 12'h222;
rom[54155] = 12'h222;
rom[54156] = 12'h222;
rom[54157] = 12'h222;
rom[54158] = 12'h222;
rom[54159] = 12'h222;
rom[54160] = 12'h222;
rom[54161] = 12'h111;
rom[54162] = 12'h111;
rom[54163] = 12'h111;
rom[54164] = 12'h111;
rom[54165] = 12'h111;
rom[54166] = 12'h111;
rom[54167] = 12'h111;
rom[54168] = 12'h111;
rom[54169] = 12'h111;
rom[54170] = 12'h111;
rom[54171] = 12'h111;
rom[54172] = 12'h111;
rom[54173] = 12'h111;
rom[54174] = 12'h111;
rom[54175] = 12'h111;
rom[54176] = 12'h111;
rom[54177] = 12'h  0;
rom[54178] = 12'h  0;
rom[54179] = 12'h  0;
rom[54180] = 12'h  0;
rom[54181] = 12'h  0;
rom[54182] = 12'h  0;
rom[54183] = 12'h  0;
rom[54184] = 12'h  0;
rom[54185] = 12'h  0;
rom[54186] = 12'h  0;
rom[54187] = 12'h  0;
rom[54188] = 12'h  0;
rom[54189] = 12'h  0;
rom[54190] = 12'h  0;
rom[54191] = 12'h  0;
rom[54192] = 12'h  0;
rom[54193] = 12'h  0;
rom[54194] = 12'h  0;
rom[54195] = 12'h  0;
rom[54196] = 12'h  0;
rom[54197] = 12'h  0;
rom[54198] = 12'h  0;
rom[54199] = 12'h  0;
rom[54200] = 12'h  0;
rom[54201] = 12'h  0;
rom[54202] = 12'h  0;
rom[54203] = 12'h  0;
rom[54204] = 12'h  0;
rom[54205] = 12'h  0;
rom[54206] = 12'h111;
rom[54207] = 12'h111;
rom[54208] = 12'h111;
rom[54209] = 12'h  0;
rom[54210] = 12'h  0;
rom[54211] = 12'h  0;
rom[54212] = 12'h111;
rom[54213] = 12'h111;
rom[54214] = 12'h111;
rom[54215] = 12'h  0;
rom[54216] = 12'h  0;
rom[54217] = 12'h  0;
rom[54218] = 12'h111;
rom[54219] = 12'h111;
rom[54220] = 12'h111;
rom[54221] = 12'h222;
rom[54222] = 12'h333;
rom[54223] = 12'h333;
rom[54224] = 12'h222;
rom[54225] = 12'h222;
rom[54226] = 12'h111;
rom[54227] = 12'h111;
rom[54228] = 12'h111;
rom[54229] = 12'h111;
rom[54230] = 12'h111;
rom[54231] = 12'h  0;
rom[54232] = 12'h  0;
rom[54233] = 12'h  0;
rom[54234] = 12'h  0;
rom[54235] = 12'h  0;
rom[54236] = 12'h  0;
rom[54237] = 12'h  0;
rom[54238] = 12'h  0;
rom[54239] = 12'h  0;
rom[54240] = 12'h  0;
rom[54241] = 12'h  0;
rom[54242] = 12'h  0;
rom[54243] = 12'h  0;
rom[54244] = 12'h  0;
rom[54245] = 12'h  0;
rom[54246] = 12'h  0;
rom[54247] = 12'h  0;
rom[54248] = 12'h  0;
rom[54249] = 12'h  0;
rom[54250] = 12'h  0;
rom[54251] = 12'h  0;
rom[54252] = 12'h  0;
rom[54253] = 12'h  0;
rom[54254] = 12'h  0;
rom[54255] = 12'h  0;
rom[54256] = 12'h  0;
rom[54257] = 12'h  0;
rom[54258] = 12'h  0;
rom[54259] = 12'h  0;
rom[54260] = 12'h  0;
rom[54261] = 12'h  0;
rom[54262] = 12'h  0;
rom[54263] = 12'h  0;
rom[54264] = 12'h  0;
rom[54265] = 12'h  0;
rom[54266] = 12'h  0;
rom[54267] = 12'h  0;
rom[54268] = 12'h  0;
rom[54269] = 12'h  0;
rom[54270] = 12'h  0;
rom[54271] = 12'h  0;
rom[54272] = 12'h111;
rom[54273] = 12'h111;
rom[54274] = 12'h222;
rom[54275] = 12'h222;
rom[54276] = 12'h333;
rom[54277] = 12'h333;
rom[54278] = 12'h222;
rom[54279] = 12'h333;
rom[54280] = 12'h333;
rom[54281] = 12'h333;
rom[54282] = 12'h333;
rom[54283] = 12'h333;
rom[54284] = 12'h444;
rom[54285] = 12'h555;
rom[54286] = 12'h555;
rom[54287] = 12'h555;
rom[54288] = 12'h444;
rom[54289] = 12'h444;
rom[54290] = 12'h444;
rom[54291] = 12'h444;
rom[54292] = 12'h555;
rom[54293] = 12'h555;
rom[54294] = 12'h666;
rom[54295] = 12'h666;
rom[54296] = 12'h777;
rom[54297] = 12'h666;
rom[54298] = 12'h666;
rom[54299] = 12'h666;
rom[54300] = 12'h777;
rom[54301] = 12'h666;
rom[54302] = 12'h666;
rom[54303] = 12'h666;
rom[54304] = 12'h666;
rom[54305] = 12'h666;
rom[54306] = 12'h666;
rom[54307] = 12'h666;
rom[54308] = 12'h666;
rom[54309] = 12'h666;
rom[54310] = 12'h555;
rom[54311] = 12'h555;
rom[54312] = 12'h666;
rom[54313] = 12'h666;
rom[54314] = 12'h555;
rom[54315] = 12'h666;
rom[54316] = 12'h666;
rom[54317] = 12'h666;
rom[54318] = 12'h666;
rom[54319] = 12'h666;
rom[54320] = 12'h666;
rom[54321] = 12'h666;
rom[54322] = 12'h666;
rom[54323] = 12'h666;
rom[54324] = 12'h555;
rom[54325] = 12'h555;
rom[54326] = 12'h555;
rom[54327] = 12'h555;
rom[54328] = 12'h555;
rom[54329] = 12'h555;
rom[54330] = 12'h555;
rom[54331] = 12'h555;
rom[54332] = 12'h555;
rom[54333] = 12'h555;
rom[54334] = 12'h555;
rom[54335] = 12'h555;
rom[54336] = 12'h666;
rom[54337] = 12'h666;
rom[54338] = 12'h666;
rom[54339] = 12'h666;
rom[54340] = 12'h666;
rom[54341] = 12'h666;
rom[54342] = 12'h666;
rom[54343] = 12'h666;
rom[54344] = 12'h666;
rom[54345] = 12'h666;
rom[54346] = 12'h666;
rom[54347] = 12'h777;
rom[54348] = 12'h777;
rom[54349] = 12'h777;
rom[54350] = 12'h777;
rom[54351] = 12'h777;
rom[54352] = 12'h888;
rom[54353] = 12'h888;
rom[54354] = 12'h888;
rom[54355] = 12'h999;
rom[54356] = 12'h999;
rom[54357] = 12'h999;
rom[54358] = 12'haaa;
rom[54359] = 12'haaa;
rom[54360] = 12'haaa;
rom[54361] = 12'hbbb;
rom[54362] = 12'hbbb;
rom[54363] = 12'hbbb;
rom[54364] = 12'hccc;
rom[54365] = 12'hccc;
rom[54366] = 12'hddd;
rom[54367] = 12'hddd;
rom[54368] = 12'hddd;
rom[54369] = 12'hddd;
rom[54370] = 12'hddd;
rom[54371] = 12'hddd;
rom[54372] = 12'hddd;
rom[54373] = 12'hddd;
rom[54374] = 12'hccc;
rom[54375] = 12'hccc;
rom[54376] = 12'hccc;
rom[54377] = 12'hccc;
rom[54378] = 12'hccc;
rom[54379] = 12'hccc;
rom[54380] = 12'hccc;
rom[54381] = 12'hccc;
rom[54382] = 12'hccc;
rom[54383] = 12'hbbb;
rom[54384] = 12'hccc;
rom[54385] = 12'hccc;
rom[54386] = 12'hccc;
rom[54387] = 12'hbbb;
rom[54388] = 12'hbbb;
rom[54389] = 12'hbbb;
rom[54390] = 12'hbbb;
rom[54391] = 12'hbbb;
rom[54392] = 12'hbbb;
rom[54393] = 12'hbbb;
rom[54394] = 12'hccc;
rom[54395] = 12'hccc;
rom[54396] = 12'hccc;
rom[54397] = 12'hccc;
rom[54398] = 12'hccc;
rom[54399] = 12'hccc;
rom[54400] = 12'hfff;
rom[54401] = 12'hfff;
rom[54402] = 12'hfff;
rom[54403] = 12'hfff;
rom[54404] = 12'hfff;
rom[54405] = 12'hfff;
rom[54406] = 12'hfff;
rom[54407] = 12'hfff;
rom[54408] = 12'hfff;
rom[54409] = 12'hfff;
rom[54410] = 12'hfff;
rom[54411] = 12'hfff;
rom[54412] = 12'heee;
rom[54413] = 12'heee;
rom[54414] = 12'hddd;
rom[54415] = 12'hddd;
rom[54416] = 12'hccc;
rom[54417] = 12'hccc;
rom[54418] = 12'hccc;
rom[54419] = 12'hccc;
rom[54420] = 12'hccc;
rom[54421] = 12'hccc;
rom[54422] = 12'hccc;
rom[54423] = 12'hccc;
rom[54424] = 12'hccc;
rom[54425] = 12'hccc;
rom[54426] = 12'hccc;
rom[54427] = 12'hccc;
rom[54428] = 12'hccc;
rom[54429] = 12'hccc;
rom[54430] = 12'hccc;
rom[54431] = 12'hccc;
rom[54432] = 12'hccc;
rom[54433] = 12'hccc;
rom[54434] = 12'hccc;
rom[54435] = 12'hccc;
rom[54436] = 12'hccc;
rom[54437] = 12'hccc;
rom[54438] = 12'hccc;
rom[54439] = 12'hccc;
rom[54440] = 12'hbbb;
rom[54441] = 12'hbbb;
rom[54442] = 12'hbbb;
rom[54443] = 12'hbbb;
rom[54444] = 12'hbbb;
rom[54445] = 12'hbbb;
rom[54446] = 12'hbbb;
rom[54447] = 12'hbbb;
rom[54448] = 12'hccc;
rom[54449] = 12'hccc;
rom[54450] = 12'hccc;
rom[54451] = 12'hccc;
rom[54452] = 12'hccc;
rom[54453] = 12'hccc;
rom[54454] = 12'hccc;
rom[54455] = 12'hccc;
rom[54456] = 12'hccc;
rom[54457] = 12'hccc;
rom[54458] = 12'hccc;
rom[54459] = 12'hddd;
rom[54460] = 12'hddd;
rom[54461] = 12'hddd;
rom[54462] = 12'hddd;
rom[54463] = 12'hddd;
rom[54464] = 12'hddd;
rom[54465] = 12'hddd;
rom[54466] = 12'hddd;
rom[54467] = 12'hddd;
rom[54468] = 12'hddd;
rom[54469] = 12'hddd;
rom[54470] = 12'hddd;
rom[54471] = 12'hddd;
rom[54472] = 12'hddd;
rom[54473] = 12'hddd;
rom[54474] = 12'hddd;
rom[54475] = 12'hddd;
rom[54476] = 12'hddd;
rom[54477] = 12'hddd;
rom[54478] = 12'hccc;
rom[54479] = 12'hccc;
rom[54480] = 12'hccc;
rom[54481] = 12'hbbb;
rom[54482] = 12'hbbb;
rom[54483] = 12'haaa;
rom[54484] = 12'haaa;
rom[54485] = 12'haaa;
rom[54486] = 12'haaa;
rom[54487] = 12'haaa;
rom[54488] = 12'haaa;
rom[54489] = 12'haaa;
rom[54490] = 12'haaa;
rom[54491] = 12'haaa;
rom[54492] = 12'haaa;
rom[54493] = 12'haaa;
rom[54494] = 12'haaa;
rom[54495] = 12'h999;
rom[54496] = 12'haaa;
rom[54497] = 12'haaa;
rom[54498] = 12'h999;
rom[54499] = 12'h999;
rom[54500] = 12'h999;
rom[54501] = 12'h999;
rom[54502] = 12'h888;
rom[54503] = 12'h888;
rom[54504] = 12'h888;
rom[54505] = 12'h888;
rom[54506] = 12'h888;
rom[54507] = 12'h777;
rom[54508] = 12'h777;
rom[54509] = 12'h888;
rom[54510] = 12'h888;
rom[54511] = 12'h888;
rom[54512] = 12'h888;
rom[54513] = 12'h888;
rom[54514] = 12'h999;
rom[54515] = 12'haaa;
rom[54516] = 12'hbbb;
rom[54517] = 12'hbbb;
rom[54518] = 12'haaa;
rom[54519] = 12'haaa;
rom[54520] = 12'h888;
rom[54521] = 12'h777;
rom[54522] = 12'h666;
rom[54523] = 12'h666;
rom[54524] = 12'h555;
rom[54525] = 12'h555;
rom[54526] = 12'h555;
rom[54527] = 12'h555;
rom[54528] = 12'h555;
rom[54529] = 12'h555;
rom[54530] = 12'h555;
rom[54531] = 12'h444;
rom[54532] = 12'h444;
rom[54533] = 12'h444;
rom[54534] = 12'h333;
rom[54535] = 12'h333;
rom[54536] = 12'h333;
rom[54537] = 12'h333;
rom[54538] = 12'h333;
rom[54539] = 12'h222;
rom[54540] = 12'h222;
rom[54541] = 12'h222;
rom[54542] = 12'h222;
rom[54543] = 12'h222;
rom[54544] = 12'h111;
rom[54545] = 12'h111;
rom[54546] = 12'h111;
rom[54547] = 12'h111;
rom[54548] = 12'h111;
rom[54549] = 12'h111;
rom[54550] = 12'h111;
rom[54551] = 12'h222;
rom[54552] = 12'h222;
rom[54553] = 12'h222;
rom[54554] = 12'h222;
rom[54555] = 12'h222;
rom[54556] = 12'h222;
rom[54557] = 12'h222;
rom[54558] = 12'h111;
rom[54559] = 12'h111;
rom[54560] = 12'h111;
rom[54561] = 12'h111;
rom[54562] = 12'h111;
rom[54563] = 12'h111;
rom[54564] = 12'h111;
rom[54565] = 12'h111;
rom[54566] = 12'h111;
rom[54567] = 12'h111;
rom[54568] = 12'h111;
rom[54569] = 12'h111;
rom[54570] = 12'h111;
rom[54571] = 12'h111;
rom[54572] = 12'h111;
rom[54573] = 12'h111;
rom[54574] = 12'h111;
rom[54575] = 12'h111;
rom[54576] = 12'h111;
rom[54577] = 12'h111;
rom[54578] = 12'h  0;
rom[54579] = 12'h  0;
rom[54580] = 12'h  0;
rom[54581] = 12'h  0;
rom[54582] = 12'h  0;
rom[54583] = 12'h  0;
rom[54584] = 12'h  0;
rom[54585] = 12'h  0;
rom[54586] = 12'h  0;
rom[54587] = 12'h  0;
rom[54588] = 12'h  0;
rom[54589] = 12'h  0;
rom[54590] = 12'h  0;
rom[54591] = 12'h  0;
rom[54592] = 12'h  0;
rom[54593] = 12'h  0;
rom[54594] = 12'h  0;
rom[54595] = 12'h  0;
rom[54596] = 12'h  0;
rom[54597] = 12'h  0;
rom[54598] = 12'h  0;
rom[54599] = 12'h  0;
rom[54600] = 12'h  0;
rom[54601] = 12'h  0;
rom[54602] = 12'h  0;
rom[54603] = 12'h  0;
rom[54604] = 12'h  0;
rom[54605] = 12'h  0;
rom[54606] = 12'h111;
rom[54607] = 12'h111;
rom[54608] = 12'h111;
rom[54609] = 12'h  0;
rom[54610] = 12'h111;
rom[54611] = 12'h111;
rom[54612] = 12'h111;
rom[54613] = 12'h111;
rom[54614] = 12'h111;
rom[54615] = 12'h  0;
rom[54616] = 12'h111;
rom[54617] = 12'h111;
rom[54618] = 12'h111;
rom[54619] = 12'h111;
rom[54620] = 12'h222;
rom[54621] = 12'h333;
rom[54622] = 12'h333;
rom[54623] = 12'h222;
rom[54624] = 12'h222;
rom[54625] = 12'h222;
rom[54626] = 12'h111;
rom[54627] = 12'h111;
rom[54628] = 12'h111;
rom[54629] = 12'h111;
rom[54630] = 12'h111;
rom[54631] = 12'h  0;
rom[54632] = 12'h  0;
rom[54633] = 12'h  0;
rom[54634] = 12'h  0;
rom[54635] = 12'h  0;
rom[54636] = 12'h  0;
rom[54637] = 12'h  0;
rom[54638] = 12'h  0;
rom[54639] = 12'h  0;
rom[54640] = 12'h  0;
rom[54641] = 12'h  0;
rom[54642] = 12'h  0;
rom[54643] = 12'h  0;
rom[54644] = 12'h  0;
rom[54645] = 12'h  0;
rom[54646] = 12'h  0;
rom[54647] = 12'h  0;
rom[54648] = 12'h  0;
rom[54649] = 12'h  0;
rom[54650] = 12'h  0;
rom[54651] = 12'h  0;
rom[54652] = 12'h  0;
rom[54653] = 12'h  0;
rom[54654] = 12'h  0;
rom[54655] = 12'h  0;
rom[54656] = 12'h  0;
rom[54657] = 12'h  0;
rom[54658] = 12'h  0;
rom[54659] = 12'h  0;
rom[54660] = 12'h  0;
rom[54661] = 12'h  0;
rom[54662] = 12'h  0;
rom[54663] = 12'h  0;
rom[54664] = 12'h  0;
rom[54665] = 12'h  0;
rom[54666] = 12'h  0;
rom[54667] = 12'h  0;
rom[54668] = 12'h  0;
rom[54669] = 12'h  0;
rom[54670] = 12'h  0;
rom[54671] = 12'h  0;
rom[54672] = 12'h111;
rom[54673] = 12'h111;
rom[54674] = 12'h222;
rom[54675] = 12'h222;
rom[54676] = 12'h222;
rom[54677] = 12'h333;
rom[54678] = 12'h333;
rom[54679] = 12'h333;
rom[54680] = 12'h333;
rom[54681] = 12'h333;
rom[54682] = 12'h333;
rom[54683] = 12'h333;
rom[54684] = 12'h555;
rom[54685] = 12'h666;
rom[54686] = 12'h555;
rom[54687] = 12'h444;
rom[54688] = 12'h333;
rom[54689] = 12'h333;
rom[54690] = 12'h444;
rom[54691] = 12'h444;
rom[54692] = 12'h444;
rom[54693] = 12'h555;
rom[54694] = 12'h555;
rom[54695] = 12'h666;
rom[54696] = 12'h777;
rom[54697] = 12'h666;
rom[54698] = 12'h666;
rom[54699] = 12'h666;
rom[54700] = 12'h666;
rom[54701] = 12'h666;
rom[54702] = 12'h666;
rom[54703] = 12'h666;
rom[54704] = 12'h666;
rom[54705] = 12'h666;
rom[54706] = 12'h666;
rom[54707] = 12'h666;
rom[54708] = 12'h666;
rom[54709] = 12'h555;
rom[54710] = 12'h555;
rom[54711] = 12'h555;
rom[54712] = 12'h555;
rom[54713] = 12'h555;
rom[54714] = 12'h555;
rom[54715] = 12'h555;
rom[54716] = 12'h555;
rom[54717] = 12'h555;
rom[54718] = 12'h555;
rom[54719] = 12'h555;
rom[54720] = 12'h555;
rom[54721] = 12'h555;
rom[54722] = 12'h666;
rom[54723] = 12'h666;
rom[54724] = 12'h666;
rom[54725] = 12'h666;
rom[54726] = 12'h666;
rom[54727] = 12'h666;
rom[54728] = 12'h555;
rom[54729] = 12'h666;
rom[54730] = 12'h666;
rom[54731] = 12'h666;
rom[54732] = 12'h666;
rom[54733] = 12'h666;
rom[54734] = 12'h666;
rom[54735] = 12'h666;
rom[54736] = 12'h666;
rom[54737] = 12'h666;
rom[54738] = 12'h666;
rom[54739] = 12'h666;
rom[54740] = 12'h666;
rom[54741] = 12'h666;
rom[54742] = 12'h666;
rom[54743] = 12'h666;
rom[54744] = 12'h666;
rom[54745] = 12'h777;
rom[54746] = 12'h777;
rom[54747] = 12'h777;
rom[54748] = 12'h777;
rom[54749] = 12'h777;
rom[54750] = 12'h777;
rom[54751] = 12'h888;
rom[54752] = 12'h888;
rom[54753] = 12'h999;
rom[54754] = 12'h999;
rom[54755] = 12'h999;
rom[54756] = 12'haaa;
rom[54757] = 12'haaa;
rom[54758] = 12'haaa;
rom[54759] = 12'haaa;
rom[54760] = 12'haaa;
rom[54761] = 12'hbbb;
rom[54762] = 12'hbbb;
rom[54763] = 12'hbbb;
rom[54764] = 12'hccc;
rom[54765] = 12'hddd;
rom[54766] = 12'hddd;
rom[54767] = 12'heee;
rom[54768] = 12'heee;
rom[54769] = 12'hddd;
rom[54770] = 12'hddd;
rom[54771] = 12'hddd;
rom[54772] = 12'hddd;
rom[54773] = 12'hccc;
rom[54774] = 12'hccc;
rom[54775] = 12'hccc;
rom[54776] = 12'hccc;
rom[54777] = 12'hccc;
rom[54778] = 12'hccc;
rom[54779] = 12'hccc;
rom[54780] = 12'hccc;
rom[54781] = 12'hccc;
rom[54782] = 12'hbbb;
rom[54783] = 12'hbbb;
rom[54784] = 12'hbbb;
rom[54785] = 12'hbbb;
rom[54786] = 12'hbbb;
rom[54787] = 12'hbbb;
rom[54788] = 12'hbbb;
rom[54789] = 12'haaa;
rom[54790] = 12'haaa;
rom[54791] = 12'haaa;
rom[54792] = 12'hbbb;
rom[54793] = 12'hbbb;
rom[54794] = 12'hbbb;
rom[54795] = 12'hbbb;
rom[54796] = 12'hbbb;
rom[54797] = 12'hbbb;
rom[54798] = 12'hbbb;
rom[54799] = 12'hbbb;
rom[54800] = 12'hfff;
rom[54801] = 12'hfff;
rom[54802] = 12'hfff;
rom[54803] = 12'hfff;
rom[54804] = 12'hfff;
rom[54805] = 12'hfff;
rom[54806] = 12'hfff;
rom[54807] = 12'hfff;
rom[54808] = 12'hfff;
rom[54809] = 12'hfff;
rom[54810] = 12'hfff;
rom[54811] = 12'hfff;
rom[54812] = 12'hfff;
rom[54813] = 12'heee;
rom[54814] = 12'heee;
rom[54815] = 12'heee;
rom[54816] = 12'hddd;
rom[54817] = 12'hddd;
rom[54818] = 12'hddd;
rom[54819] = 12'hddd;
rom[54820] = 12'hddd;
rom[54821] = 12'hddd;
rom[54822] = 12'hddd;
rom[54823] = 12'hddd;
rom[54824] = 12'hddd;
rom[54825] = 12'hddd;
rom[54826] = 12'hccc;
rom[54827] = 12'hccc;
rom[54828] = 12'hccc;
rom[54829] = 12'hccc;
rom[54830] = 12'hccc;
rom[54831] = 12'hccc;
rom[54832] = 12'hccc;
rom[54833] = 12'hccc;
rom[54834] = 12'hccc;
rom[54835] = 12'hccc;
rom[54836] = 12'hccc;
rom[54837] = 12'hccc;
rom[54838] = 12'hccc;
rom[54839] = 12'hccc;
rom[54840] = 12'hbbb;
rom[54841] = 12'hbbb;
rom[54842] = 12'hbbb;
rom[54843] = 12'hbbb;
rom[54844] = 12'hbbb;
rom[54845] = 12'hccc;
rom[54846] = 12'hccc;
rom[54847] = 12'hccc;
rom[54848] = 12'hccc;
rom[54849] = 12'hccc;
rom[54850] = 12'hccc;
rom[54851] = 12'hccc;
rom[54852] = 12'hccc;
rom[54853] = 12'hccc;
rom[54854] = 12'hccc;
rom[54855] = 12'hccc;
rom[54856] = 12'hddd;
rom[54857] = 12'hddd;
rom[54858] = 12'hddd;
rom[54859] = 12'hddd;
rom[54860] = 12'hddd;
rom[54861] = 12'hddd;
rom[54862] = 12'hddd;
rom[54863] = 12'hddd;
rom[54864] = 12'hddd;
rom[54865] = 12'hddd;
rom[54866] = 12'hddd;
rom[54867] = 12'hddd;
rom[54868] = 12'hddd;
rom[54869] = 12'heee;
rom[54870] = 12'heee;
rom[54871] = 12'heee;
rom[54872] = 12'heee;
rom[54873] = 12'heee;
rom[54874] = 12'heee;
rom[54875] = 12'heee;
rom[54876] = 12'hddd;
rom[54877] = 12'hddd;
rom[54878] = 12'hddd;
rom[54879] = 12'hddd;
rom[54880] = 12'hccc;
rom[54881] = 12'hccc;
rom[54882] = 12'hccc;
rom[54883] = 12'hbbb;
rom[54884] = 12'hbbb;
rom[54885] = 12'hbbb;
rom[54886] = 12'hbbb;
rom[54887] = 12'hbbb;
rom[54888] = 12'hbbb;
rom[54889] = 12'haaa;
rom[54890] = 12'haaa;
rom[54891] = 12'haaa;
rom[54892] = 12'haaa;
rom[54893] = 12'haaa;
rom[54894] = 12'haaa;
rom[54895] = 12'haaa;
rom[54896] = 12'haaa;
rom[54897] = 12'haaa;
rom[54898] = 12'haaa;
rom[54899] = 12'haaa;
rom[54900] = 12'haaa;
rom[54901] = 12'haaa;
rom[54902] = 12'h999;
rom[54903] = 12'h999;
rom[54904] = 12'h999;
rom[54905] = 12'h888;
rom[54906] = 12'h888;
rom[54907] = 12'h888;
rom[54908] = 12'h888;
rom[54909] = 12'h888;
rom[54910] = 12'h888;
rom[54911] = 12'h888;
rom[54912] = 12'h888;
rom[54913] = 12'h888;
rom[54914] = 12'h888;
rom[54915] = 12'h999;
rom[54916] = 12'haaa;
rom[54917] = 12'haaa;
rom[54918] = 12'hbbb;
rom[54919] = 12'hbbb;
rom[54920] = 12'haaa;
rom[54921] = 12'h999;
rom[54922] = 12'h999;
rom[54923] = 12'h888;
rom[54924] = 12'h666;
rom[54925] = 12'h666;
rom[54926] = 12'h555;
rom[54927] = 12'h555;
rom[54928] = 12'h555;
rom[54929] = 12'h444;
rom[54930] = 12'h444;
rom[54931] = 12'h555;
rom[54932] = 12'h555;
rom[54933] = 12'h555;
rom[54934] = 12'h444;
rom[54935] = 12'h444;
rom[54936] = 12'h333;
rom[54937] = 12'h333;
rom[54938] = 12'h333;
rom[54939] = 12'h333;
rom[54940] = 12'h222;
rom[54941] = 12'h222;
rom[54942] = 12'h222;
rom[54943] = 12'h222;
rom[54944] = 12'h111;
rom[54945] = 12'h111;
rom[54946] = 12'h111;
rom[54947] = 12'h111;
rom[54948] = 12'h111;
rom[54949] = 12'h222;
rom[54950] = 12'h222;
rom[54951] = 12'h222;
rom[54952] = 12'h222;
rom[54953] = 12'h222;
rom[54954] = 12'h222;
rom[54955] = 12'h222;
rom[54956] = 12'h222;
rom[54957] = 12'h222;
rom[54958] = 12'h111;
rom[54959] = 12'h111;
rom[54960] = 12'h111;
rom[54961] = 12'h111;
rom[54962] = 12'h111;
rom[54963] = 12'h111;
rom[54964] = 12'h111;
rom[54965] = 12'h111;
rom[54966] = 12'h111;
rom[54967] = 12'h111;
rom[54968] = 12'h111;
rom[54969] = 12'h111;
rom[54970] = 12'h111;
rom[54971] = 12'h111;
rom[54972] = 12'h111;
rom[54973] = 12'h111;
rom[54974] = 12'h111;
rom[54975] = 12'h  0;
rom[54976] = 12'h111;
rom[54977] = 12'h  0;
rom[54978] = 12'h  0;
rom[54979] = 12'h  0;
rom[54980] = 12'h  0;
rom[54981] = 12'h  0;
rom[54982] = 12'h  0;
rom[54983] = 12'h  0;
rom[54984] = 12'h  0;
rom[54985] = 12'h  0;
rom[54986] = 12'h  0;
rom[54987] = 12'h  0;
rom[54988] = 12'h  0;
rom[54989] = 12'h  0;
rom[54990] = 12'h  0;
rom[54991] = 12'h  0;
rom[54992] = 12'h  0;
rom[54993] = 12'h  0;
rom[54994] = 12'h  0;
rom[54995] = 12'h  0;
rom[54996] = 12'h  0;
rom[54997] = 12'h  0;
rom[54998] = 12'h  0;
rom[54999] = 12'h  0;
rom[55000] = 12'h  0;
rom[55001] = 12'h  0;
rom[55002] = 12'h  0;
rom[55003] = 12'h  0;
rom[55004] = 12'h  0;
rom[55005] = 12'h  0;
rom[55006] = 12'h111;
rom[55007] = 12'h111;
rom[55008] = 12'h111;
rom[55009] = 12'h111;
rom[55010] = 12'h111;
rom[55011] = 12'h111;
rom[55012] = 12'h111;
rom[55013] = 12'h111;
rom[55014] = 12'h111;
rom[55015] = 12'h  0;
rom[55016] = 12'h111;
rom[55017] = 12'h111;
rom[55018] = 12'h111;
rom[55019] = 12'h111;
rom[55020] = 12'h222;
rom[55021] = 12'h333;
rom[55022] = 12'h333;
rom[55023] = 12'h222;
rom[55024] = 12'h222;
rom[55025] = 12'h222;
rom[55026] = 12'h111;
rom[55027] = 12'h111;
rom[55028] = 12'h111;
rom[55029] = 12'h111;
rom[55030] = 12'h111;
rom[55031] = 12'h  0;
rom[55032] = 12'h  0;
rom[55033] = 12'h  0;
rom[55034] = 12'h  0;
rom[55035] = 12'h  0;
rom[55036] = 12'h  0;
rom[55037] = 12'h  0;
rom[55038] = 12'h  0;
rom[55039] = 12'h  0;
rom[55040] = 12'h  0;
rom[55041] = 12'h  0;
rom[55042] = 12'h  0;
rom[55043] = 12'h  0;
rom[55044] = 12'h  0;
rom[55045] = 12'h  0;
rom[55046] = 12'h  0;
rom[55047] = 12'h  0;
rom[55048] = 12'h  0;
rom[55049] = 12'h  0;
rom[55050] = 12'h  0;
rom[55051] = 12'h  0;
rom[55052] = 12'h  0;
rom[55053] = 12'h  0;
rom[55054] = 12'h  0;
rom[55055] = 12'h  0;
rom[55056] = 12'h  0;
rom[55057] = 12'h  0;
rom[55058] = 12'h  0;
rom[55059] = 12'h  0;
rom[55060] = 12'h  0;
rom[55061] = 12'h  0;
rom[55062] = 12'h  0;
rom[55063] = 12'h  0;
rom[55064] = 12'h  0;
rom[55065] = 12'h  0;
rom[55066] = 12'h  0;
rom[55067] = 12'h  0;
rom[55068] = 12'h  0;
rom[55069] = 12'h  0;
rom[55070] = 12'h  0;
rom[55071] = 12'h  0;
rom[55072] = 12'h111;
rom[55073] = 12'h111;
rom[55074] = 12'h222;
rom[55075] = 12'h222;
rom[55076] = 12'h222;
rom[55077] = 12'h333;
rom[55078] = 12'h333;
rom[55079] = 12'h333;
rom[55080] = 12'h333;
rom[55081] = 12'h333;
rom[55082] = 12'h333;
rom[55083] = 12'h444;
rom[55084] = 12'h555;
rom[55085] = 12'h666;
rom[55086] = 12'h555;
rom[55087] = 12'h444;
rom[55088] = 12'h333;
rom[55089] = 12'h333;
rom[55090] = 12'h333;
rom[55091] = 12'h444;
rom[55092] = 12'h444;
rom[55093] = 12'h555;
rom[55094] = 12'h555;
rom[55095] = 12'h666;
rom[55096] = 12'h777;
rom[55097] = 12'h666;
rom[55098] = 12'h666;
rom[55099] = 12'h666;
rom[55100] = 12'h666;
rom[55101] = 12'h666;
rom[55102] = 12'h666;
rom[55103] = 12'h666;
rom[55104] = 12'h666;
rom[55105] = 12'h666;
rom[55106] = 12'h555;
rom[55107] = 12'h666;
rom[55108] = 12'h666;
rom[55109] = 12'h555;
rom[55110] = 12'h555;
rom[55111] = 12'h555;
rom[55112] = 12'h555;
rom[55113] = 12'h555;
rom[55114] = 12'h555;
rom[55115] = 12'h555;
rom[55116] = 12'h555;
rom[55117] = 12'h555;
rom[55118] = 12'h555;
rom[55119] = 12'h555;
rom[55120] = 12'h555;
rom[55121] = 12'h555;
rom[55122] = 12'h555;
rom[55123] = 12'h555;
rom[55124] = 12'h666;
rom[55125] = 12'h666;
rom[55126] = 12'h666;
rom[55127] = 12'h666;
rom[55128] = 12'h666;
rom[55129] = 12'h666;
rom[55130] = 12'h666;
rom[55131] = 12'h666;
rom[55132] = 12'h666;
rom[55133] = 12'h666;
rom[55134] = 12'h666;
rom[55135] = 12'h666;
rom[55136] = 12'h666;
rom[55137] = 12'h666;
rom[55138] = 12'h666;
rom[55139] = 12'h666;
rom[55140] = 12'h666;
rom[55141] = 12'h777;
rom[55142] = 12'h777;
rom[55143] = 12'h777;
rom[55144] = 12'h777;
rom[55145] = 12'h777;
rom[55146] = 12'h777;
rom[55147] = 12'h777;
rom[55148] = 12'h888;
rom[55149] = 12'h888;
rom[55150] = 12'h888;
rom[55151] = 12'h888;
rom[55152] = 12'h999;
rom[55153] = 12'h999;
rom[55154] = 12'h999;
rom[55155] = 12'h999;
rom[55156] = 12'haaa;
rom[55157] = 12'haaa;
rom[55158] = 12'haaa;
rom[55159] = 12'haaa;
rom[55160] = 12'hbbb;
rom[55161] = 12'hbbb;
rom[55162] = 12'hbbb;
rom[55163] = 12'hccc;
rom[55164] = 12'hccc;
rom[55165] = 12'hddd;
rom[55166] = 12'hddd;
rom[55167] = 12'heee;
rom[55168] = 12'hddd;
rom[55169] = 12'hddd;
rom[55170] = 12'hddd;
rom[55171] = 12'hddd;
rom[55172] = 12'hccc;
rom[55173] = 12'hccc;
rom[55174] = 12'hccc;
rom[55175] = 12'hccc;
rom[55176] = 12'hccc;
rom[55177] = 12'hccc;
rom[55178] = 12'hccc;
rom[55179] = 12'hbbb;
rom[55180] = 12'hbbb;
rom[55181] = 12'hbbb;
rom[55182] = 12'hbbb;
rom[55183] = 12'hbbb;
rom[55184] = 12'hbbb;
rom[55185] = 12'hbbb;
rom[55186] = 12'hbbb;
rom[55187] = 12'haaa;
rom[55188] = 12'haaa;
rom[55189] = 12'haaa;
rom[55190] = 12'haaa;
rom[55191] = 12'haaa;
rom[55192] = 12'haaa;
rom[55193] = 12'haaa;
rom[55194] = 12'haaa;
rom[55195] = 12'haaa;
rom[55196] = 12'haaa;
rom[55197] = 12'haaa;
rom[55198] = 12'haaa;
rom[55199] = 12'haaa;
rom[55200] = 12'hfff;
rom[55201] = 12'hfff;
rom[55202] = 12'hfff;
rom[55203] = 12'hfff;
rom[55204] = 12'hfff;
rom[55205] = 12'hfff;
rom[55206] = 12'hfff;
rom[55207] = 12'hfff;
rom[55208] = 12'hfff;
rom[55209] = 12'hfff;
rom[55210] = 12'hfff;
rom[55211] = 12'hfff;
rom[55212] = 12'hfff;
rom[55213] = 12'hfff;
rom[55214] = 12'hfff;
rom[55215] = 12'hfff;
rom[55216] = 12'hfff;
rom[55217] = 12'heee;
rom[55218] = 12'heee;
rom[55219] = 12'heee;
rom[55220] = 12'heee;
rom[55221] = 12'heee;
rom[55222] = 12'heee;
rom[55223] = 12'heee;
rom[55224] = 12'hddd;
rom[55225] = 12'hddd;
rom[55226] = 12'hddd;
rom[55227] = 12'hddd;
rom[55228] = 12'hccc;
rom[55229] = 12'hccc;
rom[55230] = 12'hddd;
rom[55231] = 12'hddd;
rom[55232] = 12'hddd;
rom[55233] = 12'hddd;
rom[55234] = 12'hddd;
rom[55235] = 12'hccc;
rom[55236] = 12'hccc;
rom[55237] = 12'hccc;
rom[55238] = 12'hccc;
rom[55239] = 12'hccc;
rom[55240] = 12'hccc;
rom[55241] = 12'hccc;
rom[55242] = 12'hccc;
rom[55243] = 12'hccc;
rom[55244] = 12'hccc;
rom[55245] = 12'hccc;
rom[55246] = 12'hccc;
rom[55247] = 12'hccc;
rom[55248] = 12'hccc;
rom[55249] = 12'hccc;
rom[55250] = 12'hccc;
rom[55251] = 12'hddd;
rom[55252] = 12'hddd;
rom[55253] = 12'hddd;
rom[55254] = 12'hddd;
rom[55255] = 12'hddd;
rom[55256] = 12'hddd;
rom[55257] = 12'hddd;
rom[55258] = 12'hddd;
rom[55259] = 12'hddd;
rom[55260] = 12'heee;
rom[55261] = 12'heee;
rom[55262] = 12'heee;
rom[55263] = 12'heee;
rom[55264] = 12'heee;
rom[55265] = 12'heee;
rom[55266] = 12'heee;
rom[55267] = 12'heee;
rom[55268] = 12'heee;
rom[55269] = 12'heee;
rom[55270] = 12'heee;
rom[55271] = 12'heee;
rom[55272] = 12'heee;
rom[55273] = 12'heee;
rom[55274] = 12'heee;
rom[55275] = 12'heee;
rom[55276] = 12'heee;
rom[55277] = 12'heee;
rom[55278] = 12'hddd;
rom[55279] = 12'hddd;
rom[55280] = 12'hddd;
rom[55281] = 12'hddd;
rom[55282] = 12'hddd;
rom[55283] = 12'hddd;
rom[55284] = 12'hddd;
rom[55285] = 12'hccc;
rom[55286] = 12'hccc;
rom[55287] = 12'hccc;
rom[55288] = 12'hbbb;
rom[55289] = 12'hbbb;
rom[55290] = 12'hbbb;
rom[55291] = 12'hbbb;
rom[55292] = 12'hbbb;
rom[55293] = 12'hbbb;
rom[55294] = 12'haaa;
rom[55295] = 12'haaa;
rom[55296] = 12'h999;
rom[55297] = 12'h999;
rom[55298] = 12'h999;
rom[55299] = 12'haaa;
rom[55300] = 12'haaa;
rom[55301] = 12'haaa;
rom[55302] = 12'haaa;
rom[55303] = 12'haaa;
rom[55304] = 12'h999;
rom[55305] = 12'h999;
rom[55306] = 12'h999;
rom[55307] = 12'h999;
rom[55308] = 12'h999;
rom[55309] = 12'h888;
rom[55310] = 12'h888;
rom[55311] = 12'h777;
rom[55312] = 12'h888;
rom[55313] = 12'h888;
rom[55314] = 12'h888;
rom[55315] = 12'h888;
rom[55316] = 12'h888;
rom[55317] = 12'h999;
rom[55318] = 12'haaa;
rom[55319] = 12'haaa;
rom[55320] = 12'hbbb;
rom[55321] = 12'hbbb;
rom[55322] = 12'hbbb;
rom[55323] = 12'haaa;
rom[55324] = 12'h999;
rom[55325] = 12'h777;
rom[55326] = 12'h666;
rom[55327] = 12'h666;
rom[55328] = 12'h555;
rom[55329] = 12'h555;
rom[55330] = 12'h555;
rom[55331] = 12'h555;
rom[55332] = 12'h555;
rom[55333] = 12'h555;
rom[55334] = 12'h555;
rom[55335] = 12'h444;
rom[55336] = 12'h444;
rom[55337] = 12'h444;
rom[55338] = 12'h333;
rom[55339] = 12'h333;
rom[55340] = 12'h333;
rom[55341] = 12'h222;
rom[55342] = 12'h222;
rom[55343] = 12'h222;
rom[55344] = 12'h222;
rom[55345] = 12'h222;
rom[55346] = 12'h222;
rom[55347] = 12'h222;
rom[55348] = 12'h222;
rom[55349] = 12'h222;
rom[55350] = 12'h222;
rom[55351] = 12'h222;
rom[55352] = 12'h222;
rom[55353] = 12'h222;
rom[55354] = 12'h222;
rom[55355] = 12'h222;
rom[55356] = 12'h111;
rom[55357] = 12'h111;
rom[55358] = 12'h111;
rom[55359] = 12'h111;
rom[55360] = 12'h111;
rom[55361] = 12'h111;
rom[55362] = 12'h111;
rom[55363] = 12'h111;
rom[55364] = 12'h111;
rom[55365] = 12'h111;
rom[55366] = 12'h111;
rom[55367] = 12'h111;
rom[55368] = 12'h111;
rom[55369] = 12'h111;
rom[55370] = 12'h111;
rom[55371] = 12'h111;
rom[55372] = 12'h111;
rom[55373] = 12'h111;
rom[55374] = 12'h  0;
rom[55375] = 12'h  0;
rom[55376] = 12'h  0;
rom[55377] = 12'h  0;
rom[55378] = 12'h  0;
rom[55379] = 12'h  0;
rom[55380] = 12'h  0;
rom[55381] = 12'h  0;
rom[55382] = 12'h  0;
rom[55383] = 12'h  0;
rom[55384] = 12'h  0;
rom[55385] = 12'h  0;
rom[55386] = 12'h  0;
rom[55387] = 12'h  0;
rom[55388] = 12'h  0;
rom[55389] = 12'h  0;
rom[55390] = 12'h  0;
rom[55391] = 12'h  0;
rom[55392] = 12'h  0;
rom[55393] = 12'h  0;
rom[55394] = 12'h  0;
rom[55395] = 12'h  0;
rom[55396] = 12'h  0;
rom[55397] = 12'h  0;
rom[55398] = 12'h  0;
rom[55399] = 12'h  0;
rom[55400] = 12'h  0;
rom[55401] = 12'h  0;
rom[55402] = 12'h  0;
rom[55403] = 12'h  0;
rom[55404] = 12'h  0;
rom[55405] = 12'h  0;
rom[55406] = 12'h111;
rom[55407] = 12'h111;
rom[55408] = 12'h111;
rom[55409] = 12'h111;
rom[55410] = 12'h111;
rom[55411] = 12'h111;
rom[55412] = 12'h111;
rom[55413] = 12'h111;
rom[55414] = 12'h111;
rom[55415] = 12'h  0;
rom[55416] = 12'h  0;
rom[55417] = 12'h111;
rom[55418] = 12'h111;
rom[55419] = 12'h111;
rom[55420] = 12'h222;
rom[55421] = 12'h333;
rom[55422] = 12'h333;
rom[55423] = 12'h222;
rom[55424] = 12'h222;
rom[55425] = 12'h111;
rom[55426] = 12'h111;
rom[55427] = 12'h111;
rom[55428] = 12'h111;
rom[55429] = 12'h111;
rom[55430] = 12'h  0;
rom[55431] = 12'h  0;
rom[55432] = 12'h  0;
rom[55433] = 12'h  0;
rom[55434] = 12'h  0;
rom[55435] = 12'h  0;
rom[55436] = 12'h  0;
rom[55437] = 12'h  0;
rom[55438] = 12'h  0;
rom[55439] = 12'h  0;
rom[55440] = 12'h  0;
rom[55441] = 12'h  0;
rom[55442] = 12'h  0;
rom[55443] = 12'h  0;
rom[55444] = 12'h  0;
rom[55445] = 12'h  0;
rom[55446] = 12'h  0;
rom[55447] = 12'h  0;
rom[55448] = 12'h  0;
rom[55449] = 12'h  0;
rom[55450] = 12'h  0;
rom[55451] = 12'h  0;
rom[55452] = 12'h  0;
rom[55453] = 12'h  0;
rom[55454] = 12'h  0;
rom[55455] = 12'h  0;
rom[55456] = 12'h  0;
rom[55457] = 12'h  0;
rom[55458] = 12'h  0;
rom[55459] = 12'h  0;
rom[55460] = 12'h  0;
rom[55461] = 12'h  0;
rom[55462] = 12'h  0;
rom[55463] = 12'h  0;
rom[55464] = 12'h  0;
rom[55465] = 12'h  0;
rom[55466] = 12'h  0;
rom[55467] = 12'h  0;
rom[55468] = 12'h  0;
rom[55469] = 12'h  0;
rom[55470] = 12'h  0;
rom[55471] = 12'h  0;
rom[55472] = 12'h111;
rom[55473] = 12'h111;
rom[55474] = 12'h222;
rom[55475] = 12'h222;
rom[55476] = 12'h222;
rom[55477] = 12'h333;
rom[55478] = 12'h333;
rom[55479] = 12'h333;
rom[55480] = 12'h333;
rom[55481] = 12'h333;
rom[55482] = 12'h333;
rom[55483] = 12'h444;
rom[55484] = 12'h555;
rom[55485] = 12'h555;
rom[55486] = 12'h555;
rom[55487] = 12'h333;
rom[55488] = 12'h333;
rom[55489] = 12'h333;
rom[55490] = 12'h333;
rom[55491] = 12'h444;
rom[55492] = 12'h444;
rom[55493] = 12'h444;
rom[55494] = 12'h555;
rom[55495] = 12'h666;
rom[55496] = 12'h666;
rom[55497] = 12'h666;
rom[55498] = 12'h666;
rom[55499] = 12'h666;
rom[55500] = 12'h666;
rom[55501] = 12'h666;
rom[55502] = 12'h666;
rom[55503] = 12'h666;
rom[55504] = 12'h666;
rom[55505] = 12'h555;
rom[55506] = 12'h555;
rom[55507] = 12'h555;
rom[55508] = 12'h666;
rom[55509] = 12'h666;
rom[55510] = 12'h555;
rom[55511] = 12'h555;
rom[55512] = 12'h555;
rom[55513] = 12'h555;
rom[55514] = 12'h555;
rom[55515] = 12'h555;
rom[55516] = 12'h555;
rom[55517] = 12'h555;
rom[55518] = 12'h555;
rom[55519] = 12'h555;
rom[55520] = 12'h555;
rom[55521] = 12'h555;
rom[55522] = 12'h555;
rom[55523] = 12'h555;
rom[55524] = 12'h555;
rom[55525] = 12'h555;
rom[55526] = 12'h555;
rom[55527] = 12'h555;
rom[55528] = 12'h666;
rom[55529] = 12'h666;
rom[55530] = 12'h666;
rom[55531] = 12'h666;
rom[55532] = 12'h666;
rom[55533] = 12'h666;
rom[55534] = 12'h666;
rom[55535] = 12'h666;
rom[55536] = 12'h666;
rom[55537] = 12'h666;
rom[55538] = 12'h777;
rom[55539] = 12'h777;
rom[55540] = 12'h777;
rom[55541] = 12'h777;
rom[55542] = 12'h777;
rom[55543] = 12'h777;
rom[55544] = 12'h777;
rom[55545] = 12'h888;
rom[55546] = 12'h888;
rom[55547] = 12'h888;
rom[55548] = 12'h888;
rom[55549] = 12'h888;
rom[55550] = 12'h888;
rom[55551] = 12'h999;
rom[55552] = 12'h999;
rom[55553] = 12'h999;
rom[55554] = 12'h999;
rom[55555] = 12'haaa;
rom[55556] = 12'haaa;
rom[55557] = 12'haaa;
rom[55558] = 12'hbbb;
rom[55559] = 12'hbbb;
rom[55560] = 12'hbbb;
rom[55561] = 12'hccc;
rom[55562] = 12'hccc;
rom[55563] = 12'hddd;
rom[55564] = 12'hddd;
rom[55565] = 12'hddd;
rom[55566] = 12'hddd;
rom[55567] = 12'heee;
rom[55568] = 12'hddd;
rom[55569] = 12'hddd;
rom[55570] = 12'hddd;
rom[55571] = 12'hccc;
rom[55572] = 12'hccc;
rom[55573] = 12'hccc;
rom[55574] = 12'hccc;
rom[55575] = 12'hccc;
rom[55576] = 12'hbbb;
rom[55577] = 12'hbbb;
rom[55578] = 12'hbbb;
rom[55579] = 12'hbbb;
rom[55580] = 12'hbbb;
rom[55581] = 12'hbbb;
rom[55582] = 12'hbbb;
rom[55583] = 12'haaa;
rom[55584] = 12'haaa;
rom[55585] = 12'haaa;
rom[55586] = 12'haaa;
rom[55587] = 12'haaa;
rom[55588] = 12'haaa;
rom[55589] = 12'haaa;
rom[55590] = 12'haaa;
rom[55591] = 12'haaa;
rom[55592] = 12'haaa;
rom[55593] = 12'h999;
rom[55594] = 12'h999;
rom[55595] = 12'h999;
rom[55596] = 12'h999;
rom[55597] = 12'haaa;
rom[55598] = 12'haaa;
rom[55599] = 12'haaa;
rom[55600] = 12'hfff;
rom[55601] = 12'hfff;
rom[55602] = 12'hfff;
rom[55603] = 12'hfff;
rom[55604] = 12'hfff;
rom[55605] = 12'hfff;
rom[55606] = 12'hfff;
rom[55607] = 12'hfff;
rom[55608] = 12'hfff;
rom[55609] = 12'hfff;
rom[55610] = 12'hfff;
rom[55611] = 12'hfff;
rom[55612] = 12'hfff;
rom[55613] = 12'hfff;
rom[55614] = 12'hfff;
rom[55615] = 12'hfff;
rom[55616] = 12'hfff;
rom[55617] = 12'hfff;
rom[55618] = 12'hfff;
rom[55619] = 12'hfff;
rom[55620] = 12'heee;
rom[55621] = 12'heee;
rom[55622] = 12'heee;
rom[55623] = 12'heee;
rom[55624] = 12'heee;
rom[55625] = 12'hddd;
rom[55626] = 12'hddd;
rom[55627] = 12'hddd;
rom[55628] = 12'hddd;
rom[55629] = 12'hddd;
rom[55630] = 12'hddd;
rom[55631] = 12'hddd;
rom[55632] = 12'hddd;
rom[55633] = 12'hddd;
rom[55634] = 12'hddd;
rom[55635] = 12'hddd;
rom[55636] = 12'hddd;
rom[55637] = 12'hddd;
rom[55638] = 12'hccc;
rom[55639] = 12'hccc;
rom[55640] = 12'hccc;
rom[55641] = 12'hccc;
rom[55642] = 12'hccc;
rom[55643] = 12'hccc;
rom[55644] = 12'hccc;
rom[55645] = 12'hddd;
rom[55646] = 12'hddd;
rom[55647] = 12'hddd;
rom[55648] = 12'hddd;
rom[55649] = 12'hddd;
rom[55650] = 12'hddd;
rom[55651] = 12'hddd;
rom[55652] = 12'hddd;
rom[55653] = 12'hddd;
rom[55654] = 12'hddd;
rom[55655] = 12'heee;
rom[55656] = 12'heee;
rom[55657] = 12'heee;
rom[55658] = 12'heee;
rom[55659] = 12'heee;
rom[55660] = 12'heee;
rom[55661] = 12'heee;
rom[55662] = 12'heee;
rom[55663] = 12'heee;
rom[55664] = 12'heee;
rom[55665] = 12'heee;
rom[55666] = 12'heee;
rom[55667] = 12'heee;
rom[55668] = 12'heee;
rom[55669] = 12'heee;
rom[55670] = 12'heee;
rom[55671] = 12'hfff;
rom[55672] = 12'hfff;
rom[55673] = 12'heee;
rom[55674] = 12'heee;
rom[55675] = 12'heee;
rom[55676] = 12'heee;
rom[55677] = 12'heee;
rom[55678] = 12'heee;
rom[55679] = 12'heee;
rom[55680] = 12'heee;
rom[55681] = 12'hddd;
rom[55682] = 12'hddd;
rom[55683] = 12'hddd;
rom[55684] = 12'hddd;
rom[55685] = 12'hddd;
rom[55686] = 12'hddd;
rom[55687] = 12'hccc;
rom[55688] = 12'hccc;
rom[55689] = 12'hccc;
rom[55690] = 12'hbbb;
rom[55691] = 12'hbbb;
rom[55692] = 12'hbbb;
rom[55693] = 12'hbbb;
rom[55694] = 12'hbbb;
rom[55695] = 12'hbbb;
rom[55696] = 12'haaa;
rom[55697] = 12'haaa;
rom[55698] = 12'h999;
rom[55699] = 12'h999;
rom[55700] = 12'h999;
rom[55701] = 12'h999;
rom[55702] = 12'h999;
rom[55703] = 12'h999;
rom[55704] = 12'haaa;
rom[55705] = 12'haaa;
rom[55706] = 12'h999;
rom[55707] = 12'h999;
rom[55708] = 12'h999;
rom[55709] = 12'h999;
rom[55710] = 12'h888;
rom[55711] = 12'h888;
rom[55712] = 12'h888;
rom[55713] = 12'h888;
rom[55714] = 12'h888;
rom[55715] = 12'h888;
rom[55716] = 12'h777;
rom[55717] = 12'h888;
rom[55718] = 12'h888;
rom[55719] = 12'h888;
rom[55720] = 12'h999;
rom[55721] = 12'haaa;
rom[55722] = 12'hbbb;
rom[55723] = 12'hbbb;
rom[55724] = 12'hbbb;
rom[55725] = 12'haaa;
rom[55726] = 12'h888;
rom[55727] = 12'h888;
rom[55728] = 12'h777;
rom[55729] = 12'h666;
rom[55730] = 12'h666;
rom[55731] = 12'h666;
rom[55732] = 12'h555;
rom[55733] = 12'h555;
rom[55734] = 12'h555;
rom[55735] = 12'h555;
rom[55736] = 12'h555;
rom[55737] = 12'h444;
rom[55738] = 12'h444;
rom[55739] = 12'h444;
rom[55740] = 12'h333;
rom[55741] = 12'h333;
rom[55742] = 12'h333;
rom[55743] = 12'h333;
rom[55744] = 12'h333;
rom[55745] = 12'h333;
rom[55746] = 12'h333;
rom[55747] = 12'h333;
rom[55748] = 12'h333;
rom[55749] = 12'h333;
rom[55750] = 12'h333;
rom[55751] = 12'h333;
rom[55752] = 12'h222;
rom[55753] = 12'h222;
rom[55754] = 12'h222;
rom[55755] = 12'h111;
rom[55756] = 12'h111;
rom[55757] = 12'h111;
rom[55758] = 12'h111;
rom[55759] = 12'h111;
rom[55760] = 12'h111;
rom[55761] = 12'h111;
rom[55762] = 12'h111;
rom[55763] = 12'h111;
rom[55764] = 12'h111;
rom[55765] = 12'h111;
rom[55766] = 12'h111;
rom[55767] = 12'h111;
rom[55768] = 12'h111;
rom[55769] = 12'h111;
rom[55770] = 12'h111;
rom[55771] = 12'h111;
rom[55772] = 12'h111;
rom[55773] = 12'h111;
rom[55774] = 12'h111;
rom[55775] = 12'h  0;
rom[55776] = 12'h  0;
rom[55777] = 12'h  0;
rom[55778] = 12'h  0;
rom[55779] = 12'h  0;
rom[55780] = 12'h  0;
rom[55781] = 12'h  0;
rom[55782] = 12'h  0;
rom[55783] = 12'h  0;
rom[55784] = 12'h  0;
rom[55785] = 12'h  0;
rom[55786] = 12'h  0;
rom[55787] = 12'h  0;
rom[55788] = 12'h  0;
rom[55789] = 12'h  0;
rom[55790] = 12'h  0;
rom[55791] = 12'h  0;
rom[55792] = 12'h  0;
rom[55793] = 12'h  0;
rom[55794] = 12'h  0;
rom[55795] = 12'h  0;
rom[55796] = 12'h  0;
rom[55797] = 12'h  0;
rom[55798] = 12'h  0;
rom[55799] = 12'h  0;
rom[55800] = 12'h  0;
rom[55801] = 12'h  0;
rom[55802] = 12'h  0;
rom[55803] = 12'h  0;
rom[55804] = 12'h  0;
rom[55805] = 12'h  0;
rom[55806] = 12'h111;
rom[55807] = 12'h111;
rom[55808] = 12'h111;
rom[55809] = 12'h111;
rom[55810] = 12'h111;
rom[55811] = 12'h111;
rom[55812] = 12'h111;
rom[55813] = 12'h111;
rom[55814] = 12'h111;
rom[55815] = 12'h  0;
rom[55816] = 12'h  0;
rom[55817] = 12'h111;
rom[55818] = 12'h222;
rom[55819] = 12'h222;
rom[55820] = 12'h333;
rom[55821] = 12'h333;
rom[55822] = 12'h222;
rom[55823] = 12'h222;
rom[55824] = 12'h111;
rom[55825] = 12'h111;
rom[55826] = 12'h111;
rom[55827] = 12'h111;
rom[55828] = 12'h111;
rom[55829] = 12'h111;
rom[55830] = 12'h  0;
rom[55831] = 12'h  0;
rom[55832] = 12'h  0;
rom[55833] = 12'h  0;
rom[55834] = 12'h  0;
rom[55835] = 12'h  0;
rom[55836] = 12'h  0;
rom[55837] = 12'h  0;
rom[55838] = 12'h  0;
rom[55839] = 12'h  0;
rom[55840] = 12'h  0;
rom[55841] = 12'h  0;
rom[55842] = 12'h  0;
rom[55843] = 12'h  0;
rom[55844] = 12'h  0;
rom[55845] = 12'h  0;
rom[55846] = 12'h  0;
rom[55847] = 12'h  0;
rom[55848] = 12'h  0;
rom[55849] = 12'h  0;
rom[55850] = 12'h  0;
rom[55851] = 12'h  0;
rom[55852] = 12'h  0;
rom[55853] = 12'h  0;
rom[55854] = 12'h  0;
rom[55855] = 12'h  0;
rom[55856] = 12'h  0;
rom[55857] = 12'h  0;
rom[55858] = 12'h  0;
rom[55859] = 12'h  0;
rom[55860] = 12'h  0;
rom[55861] = 12'h  0;
rom[55862] = 12'h  0;
rom[55863] = 12'h  0;
rom[55864] = 12'h  0;
rom[55865] = 12'h  0;
rom[55866] = 12'h  0;
rom[55867] = 12'h  0;
rom[55868] = 12'h  0;
rom[55869] = 12'h  0;
rom[55870] = 12'h  0;
rom[55871] = 12'h  0;
rom[55872] = 12'h111;
rom[55873] = 12'h111;
rom[55874] = 12'h222;
rom[55875] = 12'h222;
rom[55876] = 12'h222;
rom[55877] = 12'h222;
rom[55878] = 12'h333;
rom[55879] = 12'h333;
rom[55880] = 12'h333;
rom[55881] = 12'h333;
rom[55882] = 12'h333;
rom[55883] = 12'h444;
rom[55884] = 12'h555;
rom[55885] = 12'h555;
rom[55886] = 12'h444;
rom[55887] = 12'h333;
rom[55888] = 12'h333;
rom[55889] = 12'h333;
rom[55890] = 12'h333;
rom[55891] = 12'h333;
rom[55892] = 12'h444;
rom[55893] = 12'h444;
rom[55894] = 12'h555;
rom[55895] = 12'h555;
rom[55896] = 12'h666;
rom[55897] = 12'h666;
rom[55898] = 12'h666;
rom[55899] = 12'h666;
rom[55900] = 12'h555;
rom[55901] = 12'h555;
rom[55902] = 12'h666;
rom[55903] = 12'h666;
rom[55904] = 12'h666;
rom[55905] = 12'h555;
rom[55906] = 12'h555;
rom[55907] = 12'h555;
rom[55908] = 12'h555;
rom[55909] = 12'h666;
rom[55910] = 12'h666;
rom[55911] = 12'h555;
rom[55912] = 12'h666;
rom[55913] = 12'h555;
rom[55914] = 12'h555;
rom[55915] = 12'h555;
rom[55916] = 12'h555;
rom[55917] = 12'h555;
rom[55918] = 12'h555;
rom[55919] = 12'h555;
rom[55920] = 12'h555;
rom[55921] = 12'h555;
rom[55922] = 12'h555;
rom[55923] = 12'h555;
rom[55924] = 12'h555;
rom[55925] = 12'h555;
rom[55926] = 12'h555;
rom[55927] = 12'h555;
rom[55928] = 12'h666;
rom[55929] = 12'h666;
rom[55930] = 12'h666;
rom[55931] = 12'h666;
rom[55932] = 12'h666;
rom[55933] = 12'h666;
rom[55934] = 12'h666;
rom[55935] = 12'h666;
rom[55936] = 12'h777;
rom[55937] = 12'h777;
rom[55938] = 12'h777;
rom[55939] = 12'h777;
rom[55940] = 12'h777;
rom[55941] = 12'h777;
rom[55942] = 12'h777;
rom[55943] = 12'h777;
rom[55944] = 12'h888;
rom[55945] = 12'h888;
rom[55946] = 12'h888;
rom[55947] = 12'h888;
rom[55948] = 12'h888;
rom[55949] = 12'h999;
rom[55950] = 12'h999;
rom[55951] = 12'h999;
rom[55952] = 12'h999;
rom[55953] = 12'h999;
rom[55954] = 12'h999;
rom[55955] = 12'haaa;
rom[55956] = 12'haaa;
rom[55957] = 12'haaa;
rom[55958] = 12'hbbb;
rom[55959] = 12'hbbb;
rom[55960] = 12'hbbb;
rom[55961] = 12'hccc;
rom[55962] = 12'hccc;
rom[55963] = 12'hddd;
rom[55964] = 12'heee;
rom[55965] = 12'heee;
rom[55966] = 12'heee;
rom[55967] = 12'hddd;
rom[55968] = 12'hddd;
rom[55969] = 12'hddd;
rom[55970] = 12'hccc;
rom[55971] = 12'hccc;
rom[55972] = 12'hccc;
rom[55973] = 12'hccc;
rom[55974] = 12'hccc;
rom[55975] = 12'hbbb;
rom[55976] = 12'hbbb;
rom[55977] = 12'hbbb;
rom[55978] = 12'hbbb;
rom[55979] = 12'hbbb;
rom[55980] = 12'hbbb;
rom[55981] = 12'hbbb;
rom[55982] = 12'haaa;
rom[55983] = 12'haaa;
rom[55984] = 12'haaa;
rom[55985] = 12'haaa;
rom[55986] = 12'haaa;
rom[55987] = 12'haaa;
rom[55988] = 12'h999;
rom[55989] = 12'h999;
rom[55990] = 12'h999;
rom[55991] = 12'h999;
rom[55992] = 12'h999;
rom[55993] = 12'h999;
rom[55994] = 12'h999;
rom[55995] = 12'h999;
rom[55996] = 12'h999;
rom[55997] = 12'h999;
rom[55998] = 12'haaa;
rom[55999] = 12'haaa;
rom[56000] = 12'hfff;
rom[56001] = 12'hfff;
rom[56002] = 12'hfff;
rom[56003] = 12'hfff;
rom[56004] = 12'hfff;
rom[56005] = 12'hfff;
rom[56006] = 12'hfff;
rom[56007] = 12'hfff;
rom[56008] = 12'hfff;
rom[56009] = 12'hfff;
rom[56010] = 12'hfff;
rom[56011] = 12'hfff;
rom[56012] = 12'hfff;
rom[56013] = 12'hfff;
rom[56014] = 12'hfff;
rom[56015] = 12'hfff;
rom[56016] = 12'hfff;
rom[56017] = 12'hfff;
rom[56018] = 12'hfff;
rom[56019] = 12'hfff;
rom[56020] = 12'hfff;
rom[56021] = 12'hfff;
rom[56022] = 12'hfff;
rom[56023] = 12'hfff;
rom[56024] = 12'heee;
rom[56025] = 12'heee;
rom[56026] = 12'heee;
rom[56027] = 12'heee;
rom[56028] = 12'heee;
rom[56029] = 12'heee;
rom[56030] = 12'heee;
rom[56031] = 12'heee;
rom[56032] = 12'hddd;
rom[56033] = 12'hddd;
rom[56034] = 12'hddd;
rom[56035] = 12'hddd;
rom[56036] = 12'hddd;
rom[56037] = 12'hddd;
rom[56038] = 12'hddd;
rom[56039] = 12'hddd;
rom[56040] = 12'hddd;
rom[56041] = 12'hddd;
rom[56042] = 12'hddd;
rom[56043] = 12'hddd;
rom[56044] = 12'hddd;
rom[56045] = 12'hddd;
rom[56046] = 12'hddd;
rom[56047] = 12'hddd;
rom[56048] = 12'hddd;
rom[56049] = 12'hddd;
rom[56050] = 12'heee;
rom[56051] = 12'heee;
rom[56052] = 12'heee;
rom[56053] = 12'heee;
rom[56054] = 12'heee;
rom[56055] = 12'heee;
rom[56056] = 12'heee;
rom[56057] = 12'heee;
rom[56058] = 12'heee;
rom[56059] = 12'heee;
rom[56060] = 12'heee;
rom[56061] = 12'hfff;
rom[56062] = 12'heee;
rom[56063] = 12'heee;
rom[56064] = 12'hfff;
rom[56065] = 12'hfff;
rom[56066] = 12'hfff;
rom[56067] = 12'hfff;
rom[56068] = 12'hfff;
rom[56069] = 12'hfff;
rom[56070] = 12'hfff;
rom[56071] = 12'hfff;
rom[56072] = 12'hfff;
rom[56073] = 12'hfff;
rom[56074] = 12'hfff;
rom[56075] = 12'hfff;
rom[56076] = 12'hfff;
rom[56077] = 12'hfff;
rom[56078] = 12'heee;
rom[56079] = 12'heee;
rom[56080] = 12'heee;
rom[56081] = 12'heee;
rom[56082] = 12'hddd;
rom[56083] = 12'hddd;
rom[56084] = 12'hddd;
rom[56085] = 12'hddd;
rom[56086] = 12'hddd;
rom[56087] = 12'hddd;
rom[56088] = 12'hccc;
rom[56089] = 12'hccc;
rom[56090] = 12'hccc;
rom[56091] = 12'hccc;
rom[56092] = 12'hccc;
rom[56093] = 12'hccc;
rom[56094] = 12'hccc;
rom[56095] = 12'hccc;
rom[56096] = 12'hbbb;
rom[56097] = 12'hbbb;
rom[56098] = 12'haaa;
rom[56099] = 12'haaa;
rom[56100] = 12'h999;
rom[56101] = 12'h999;
rom[56102] = 12'h999;
rom[56103] = 12'h999;
rom[56104] = 12'h999;
rom[56105] = 12'h999;
rom[56106] = 12'h999;
rom[56107] = 12'h999;
rom[56108] = 12'h999;
rom[56109] = 12'h999;
rom[56110] = 12'h999;
rom[56111] = 12'h888;
rom[56112] = 12'h888;
rom[56113] = 12'h888;
rom[56114] = 12'h888;
rom[56115] = 12'h888;
rom[56116] = 12'h888;
rom[56117] = 12'h888;
rom[56118] = 12'h888;
rom[56119] = 12'h777;
rom[56120] = 12'h888;
rom[56121] = 12'h888;
rom[56122] = 12'h999;
rom[56123] = 12'haaa;
rom[56124] = 12'hbbb;
rom[56125] = 12'hbbb;
rom[56126] = 12'haaa;
rom[56127] = 12'haaa;
rom[56128] = 12'h888;
rom[56129] = 12'h888;
rom[56130] = 12'h777;
rom[56131] = 12'h666;
rom[56132] = 12'h666;
rom[56133] = 12'h666;
rom[56134] = 12'h666;
rom[56135] = 12'h666;
rom[56136] = 12'h555;
rom[56137] = 12'h555;
rom[56138] = 12'h555;
rom[56139] = 12'h555;
rom[56140] = 12'h444;
rom[56141] = 12'h444;
rom[56142] = 12'h444;
rom[56143] = 12'h444;
rom[56144] = 12'h444;
rom[56145] = 12'h444;
rom[56146] = 12'h333;
rom[56147] = 12'h333;
rom[56148] = 12'h333;
rom[56149] = 12'h333;
rom[56150] = 12'h333;
rom[56151] = 12'h333;
rom[56152] = 12'h222;
rom[56153] = 12'h222;
rom[56154] = 12'h222;
rom[56155] = 12'h222;
rom[56156] = 12'h222;
rom[56157] = 12'h222;
rom[56158] = 12'h222;
rom[56159] = 12'h222;
rom[56160] = 12'h111;
rom[56161] = 12'h111;
rom[56162] = 12'h111;
rom[56163] = 12'h111;
rom[56164] = 12'h111;
rom[56165] = 12'h111;
rom[56166] = 12'h111;
rom[56167] = 12'h111;
rom[56168] = 12'h111;
rom[56169] = 12'h111;
rom[56170] = 12'h111;
rom[56171] = 12'h111;
rom[56172] = 12'h111;
rom[56173] = 12'h111;
rom[56174] = 12'h111;
rom[56175] = 12'h  0;
rom[56176] = 12'h  0;
rom[56177] = 12'h  0;
rom[56178] = 12'h  0;
rom[56179] = 12'h  0;
rom[56180] = 12'h  0;
rom[56181] = 12'h  0;
rom[56182] = 12'h  0;
rom[56183] = 12'h  0;
rom[56184] = 12'h  0;
rom[56185] = 12'h  0;
rom[56186] = 12'h  0;
rom[56187] = 12'h  0;
rom[56188] = 12'h  0;
rom[56189] = 12'h  0;
rom[56190] = 12'h  0;
rom[56191] = 12'h  0;
rom[56192] = 12'h  0;
rom[56193] = 12'h  0;
rom[56194] = 12'h  0;
rom[56195] = 12'h  0;
rom[56196] = 12'h  0;
rom[56197] = 12'h  0;
rom[56198] = 12'h  0;
rom[56199] = 12'h  0;
rom[56200] = 12'h  0;
rom[56201] = 12'h  0;
rom[56202] = 12'h  0;
rom[56203] = 12'h  0;
rom[56204] = 12'h  0;
rom[56205] = 12'h111;
rom[56206] = 12'h111;
rom[56207] = 12'h111;
rom[56208] = 12'h111;
rom[56209] = 12'h111;
rom[56210] = 12'h111;
rom[56211] = 12'h111;
rom[56212] = 12'h111;
rom[56213] = 12'h111;
rom[56214] = 12'h111;
rom[56215] = 12'h  0;
rom[56216] = 12'h111;
rom[56217] = 12'h111;
rom[56218] = 12'h222;
rom[56219] = 12'h333;
rom[56220] = 12'h333;
rom[56221] = 12'h333;
rom[56222] = 12'h222;
rom[56223] = 12'h111;
rom[56224] = 12'h111;
rom[56225] = 12'h111;
rom[56226] = 12'h111;
rom[56227] = 12'h111;
rom[56228] = 12'h111;
rom[56229] = 12'h  0;
rom[56230] = 12'h  0;
rom[56231] = 12'h  0;
rom[56232] = 12'h  0;
rom[56233] = 12'h  0;
rom[56234] = 12'h  0;
rom[56235] = 12'h  0;
rom[56236] = 12'h  0;
rom[56237] = 12'h  0;
rom[56238] = 12'h  0;
rom[56239] = 12'h  0;
rom[56240] = 12'h  0;
rom[56241] = 12'h  0;
rom[56242] = 12'h  0;
rom[56243] = 12'h  0;
rom[56244] = 12'h  0;
rom[56245] = 12'h  0;
rom[56246] = 12'h  0;
rom[56247] = 12'h  0;
rom[56248] = 12'h  0;
rom[56249] = 12'h  0;
rom[56250] = 12'h  0;
rom[56251] = 12'h  0;
rom[56252] = 12'h  0;
rom[56253] = 12'h  0;
rom[56254] = 12'h  0;
rom[56255] = 12'h  0;
rom[56256] = 12'h  0;
rom[56257] = 12'h  0;
rom[56258] = 12'h  0;
rom[56259] = 12'h  0;
rom[56260] = 12'h  0;
rom[56261] = 12'h  0;
rom[56262] = 12'h  0;
rom[56263] = 12'h  0;
rom[56264] = 12'h  0;
rom[56265] = 12'h  0;
rom[56266] = 12'h  0;
rom[56267] = 12'h  0;
rom[56268] = 12'h  0;
rom[56269] = 12'h  0;
rom[56270] = 12'h  0;
rom[56271] = 12'h  0;
rom[56272] = 12'h111;
rom[56273] = 12'h111;
rom[56274] = 12'h222;
rom[56275] = 12'h222;
rom[56276] = 12'h222;
rom[56277] = 12'h222;
rom[56278] = 12'h333;
rom[56279] = 12'h333;
rom[56280] = 12'h333;
rom[56281] = 12'h333;
rom[56282] = 12'h444;
rom[56283] = 12'h555;
rom[56284] = 12'h555;
rom[56285] = 12'h555;
rom[56286] = 12'h444;
rom[56287] = 12'h333;
rom[56288] = 12'h333;
rom[56289] = 12'h333;
rom[56290] = 12'h333;
rom[56291] = 12'h333;
rom[56292] = 12'h333;
rom[56293] = 12'h444;
rom[56294] = 12'h444;
rom[56295] = 12'h555;
rom[56296] = 12'h666;
rom[56297] = 12'h666;
rom[56298] = 12'h666;
rom[56299] = 12'h666;
rom[56300] = 12'h555;
rom[56301] = 12'h555;
rom[56302] = 12'h666;
rom[56303] = 12'h666;
rom[56304] = 12'h666;
rom[56305] = 12'h666;
rom[56306] = 12'h555;
rom[56307] = 12'h555;
rom[56308] = 12'h555;
rom[56309] = 12'h666;
rom[56310] = 12'h666;
rom[56311] = 12'h555;
rom[56312] = 12'h666;
rom[56313] = 12'h555;
rom[56314] = 12'h555;
rom[56315] = 12'h555;
rom[56316] = 12'h555;
rom[56317] = 12'h555;
rom[56318] = 12'h555;
rom[56319] = 12'h555;
rom[56320] = 12'h555;
rom[56321] = 12'h555;
rom[56322] = 12'h555;
rom[56323] = 12'h555;
rom[56324] = 12'h555;
rom[56325] = 12'h555;
rom[56326] = 12'h555;
rom[56327] = 12'h555;
rom[56328] = 12'h555;
rom[56329] = 12'h555;
rom[56330] = 12'h666;
rom[56331] = 12'h666;
rom[56332] = 12'h666;
rom[56333] = 12'h666;
rom[56334] = 12'h666;
rom[56335] = 12'h666;
rom[56336] = 12'h777;
rom[56337] = 12'h777;
rom[56338] = 12'h777;
rom[56339] = 12'h777;
rom[56340] = 12'h777;
rom[56341] = 12'h777;
rom[56342] = 12'h777;
rom[56343] = 12'h888;
rom[56344] = 12'h888;
rom[56345] = 12'h888;
rom[56346] = 12'h888;
rom[56347] = 12'h888;
rom[56348] = 12'h999;
rom[56349] = 12'h999;
rom[56350] = 12'h999;
rom[56351] = 12'h999;
rom[56352] = 12'haaa;
rom[56353] = 12'haaa;
rom[56354] = 12'haaa;
rom[56355] = 12'haaa;
rom[56356] = 12'haaa;
rom[56357] = 12'hbbb;
rom[56358] = 12'hbbb;
rom[56359] = 12'hbbb;
rom[56360] = 12'hccc;
rom[56361] = 12'hccc;
rom[56362] = 12'hddd;
rom[56363] = 12'hddd;
rom[56364] = 12'heee;
rom[56365] = 12'heee;
rom[56366] = 12'hddd;
rom[56367] = 12'hddd;
rom[56368] = 12'hddd;
rom[56369] = 12'hccc;
rom[56370] = 12'hccc;
rom[56371] = 12'hccc;
rom[56372] = 12'hccc;
rom[56373] = 12'hbbb;
rom[56374] = 12'hbbb;
rom[56375] = 12'hbbb;
rom[56376] = 12'hbbb;
rom[56377] = 12'hbbb;
rom[56378] = 12'haaa;
rom[56379] = 12'haaa;
rom[56380] = 12'haaa;
rom[56381] = 12'haaa;
rom[56382] = 12'haaa;
rom[56383] = 12'haaa;
rom[56384] = 12'haaa;
rom[56385] = 12'haaa;
rom[56386] = 12'h999;
rom[56387] = 12'h999;
rom[56388] = 12'h999;
rom[56389] = 12'h999;
rom[56390] = 12'h999;
rom[56391] = 12'h999;
rom[56392] = 12'h999;
rom[56393] = 12'h999;
rom[56394] = 12'h999;
rom[56395] = 12'h999;
rom[56396] = 12'h999;
rom[56397] = 12'h999;
rom[56398] = 12'haaa;
rom[56399] = 12'haaa;
rom[56400] = 12'hfff;
rom[56401] = 12'hfff;
rom[56402] = 12'hfff;
rom[56403] = 12'hfff;
rom[56404] = 12'hfff;
rom[56405] = 12'hfff;
rom[56406] = 12'hfff;
rom[56407] = 12'hfff;
rom[56408] = 12'hfff;
rom[56409] = 12'hfff;
rom[56410] = 12'hfff;
rom[56411] = 12'hfff;
rom[56412] = 12'hfff;
rom[56413] = 12'hfff;
rom[56414] = 12'hfff;
rom[56415] = 12'hfff;
rom[56416] = 12'hfff;
rom[56417] = 12'hfff;
rom[56418] = 12'hfff;
rom[56419] = 12'hfff;
rom[56420] = 12'hfff;
rom[56421] = 12'hfff;
rom[56422] = 12'hfff;
rom[56423] = 12'hfff;
rom[56424] = 12'hfff;
rom[56425] = 12'hfff;
rom[56426] = 12'hfff;
rom[56427] = 12'hfff;
rom[56428] = 12'heee;
rom[56429] = 12'heee;
rom[56430] = 12'heee;
rom[56431] = 12'heee;
rom[56432] = 12'heee;
rom[56433] = 12'heee;
rom[56434] = 12'heee;
rom[56435] = 12'heee;
rom[56436] = 12'heee;
rom[56437] = 12'heee;
rom[56438] = 12'heee;
rom[56439] = 12'heee;
rom[56440] = 12'heee;
rom[56441] = 12'heee;
rom[56442] = 12'heee;
rom[56443] = 12'heee;
rom[56444] = 12'heee;
rom[56445] = 12'heee;
rom[56446] = 12'heee;
rom[56447] = 12'heee;
rom[56448] = 12'heee;
rom[56449] = 12'heee;
rom[56450] = 12'heee;
rom[56451] = 12'heee;
rom[56452] = 12'heee;
rom[56453] = 12'hfff;
rom[56454] = 12'hfff;
rom[56455] = 12'hfff;
rom[56456] = 12'hfff;
rom[56457] = 12'hfff;
rom[56458] = 12'hfff;
rom[56459] = 12'hfff;
rom[56460] = 12'hfff;
rom[56461] = 12'hfff;
rom[56462] = 12'hfff;
rom[56463] = 12'hfff;
rom[56464] = 12'hfff;
rom[56465] = 12'hfff;
rom[56466] = 12'hfff;
rom[56467] = 12'hfff;
rom[56468] = 12'hfff;
rom[56469] = 12'hfff;
rom[56470] = 12'hfff;
rom[56471] = 12'hfff;
rom[56472] = 12'hfff;
rom[56473] = 12'hfff;
rom[56474] = 12'hfff;
rom[56475] = 12'hfff;
rom[56476] = 12'hfff;
rom[56477] = 12'hfff;
rom[56478] = 12'hfff;
rom[56479] = 12'hfff;
rom[56480] = 12'heee;
rom[56481] = 12'heee;
rom[56482] = 12'heee;
rom[56483] = 12'hddd;
rom[56484] = 12'hddd;
rom[56485] = 12'hddd;
rom[56486] = 12'hddd;
rom[56487] = 12'hddd;
rom[56488] = 12'hddd;
rom[56489] = 12'hccc;
rom[56490] = 12'hccc;
rom[56491] = 12'hccc;
rom[56492] = 12'hccc;
rom[56493] = 12'hddd;
rom[56494] = 12'hccc;
rom[56495] = 12'hccc;
rom[56496] = 12'hddd;
rom[56497] = 12'hccc;
rom[56498] = 12'hccc;
rom[56499] = 12'hbbb;
rom[56500] = 12'hbbb;
rom[56501] = 12'haaa;
rom[56502] = 12'haaa;
rom[56503] = 12'haaa;
rom[56504] = 12'h999;
rom[56505] = 12'h999;
rom[56506] = 12'h999;
rom[56507] = 12'h999;
rom[56508] = 12'haaa;
rom[56509] = 12'haaa;
rom[56510] = 12'haaa;
rom[56511] = 12'h999;
rom[56512] = 12'h999;
rom[56513] = 12'h888;
rom[56514] = 12'h888;
rom[56515] = 12'h888;
rom[56516] = 12'h888;
rom[56517] = 12'h888;
rom[56518] = 12'h777;
rom[56519] = 12'h777;
rom[56520] = 12'h777;
rom[56521] = 12'h777;
rom[56522] = 12'h777;
rom[56523] = 12'h888;
rom[56524] = 12'h999;
rom[56525] = 12'haaa;
rom[56526] = 12'hbbb;
rom[56527] = 12'hbbb;
rom[56528] = 12'h999;
rom[56529] = 12'h999;
rom[56530] = 12'h888;
rom[56531] = 12'h777;
rom[56532] = 12'h777;
rom[56533] = 12'h666;
rom[56534] = 12'h666;
rom[56535] = 12'h666;
rom[56536] = 12'h666;
rom[56537] = 12'h555;
rom[56538] = 12'h555;
rom[56539] = 12'h555;
rom[56540] = 12'h555;
rom[56541] = 12'h555;
rom[56542] = 12'h444;
rom[56543] = 12'h444;
rom[56544] = 12'h444;
rom[56545] = 12'h444;
rom[56546] = 12'h444;
rom[56547] = 12'h333;
rom[56548] = 12'h333;
rom[56549] = 12'h333;
rom[56550] = 12'h333;
rom[56551] = 12'h333;
rom[56552] = 12'h333;
rom[56553] = 12'h222;
rom[56554] = 12'h222;
rom[56555] = 12'h222;
rom[56556] = 12'h222;
rom[56557] = 12'h222;
rom[56558] = 12'h222;
rom[56559] = 12'h222;
rom[56560] = 12'h111;
rom[56561] = 12'h111;
rom[56562] = 12'h111;
rom[56563] = 12'h111;
rom[56564] = 12'h111;
rom[56565] = 12'h111;
rom[56566] = 12'h111;
rom[56567] = 12'h111;
rom[56568] = 12'h111;
rom[56569] = 12'h111;
rom[56570] = 12'h111;
rom[56571] = 12'h111;
rom[56572] = 12'h111;
rom[56573] = 12'h111;
rom[56574] = 12'h111;
rom[56575] = 12'h  0;
rom[56576] = 12'h  0;
rom[56577] = 12'h  0;
rom[56578] = 12'h  0;
rom[56579] = 12'h  0;
rom[56580] = 12'h  0;
rom[56581] = 12'h  0;
rom[56582] = 12'h  0;
rom[56583] = 12'h  0;
rom[56584] = 12'h  0;
rom[56585] = 12'h  0;
rom[56586] = 12'h  0;
rom[56587] = 12'h  0;
rom[56588] = 12'h  0;
rom[56589] = 12'h  0;
rom[56590] = 12'h  0;
rom[56591] = 12'h  0;
rom[56592] = 12'h  0;
rom[56593] = 12'h  0;
rom[56594] = 12'h  0;
rom[56595] = 12'h  0;
rom[56596] = 12'h  0;
rom[56597] = 12'h  0;
rom[56598] = 12'h  0;
rom[56599] = 12'h  0;
rom[56600] = 12'h  0;
rom[56601] = 12'h  0;
rom[56602] = 12'h  0;
rom[56603] = 12'h  0;
rom[56604] = 12'h  0;
rom[56605] = 12'h111;
rom[56606] = 12'h111;
rom[56607] = 12'h111;
rom[56608] = 12'h111;
rom[56609] = 12'h111;
rom[56610] = 12'h  0;
rom[56611] = 12'h  0;
rom[56612] = 12'h111;
rom[56613] = 12'h111;
rom[56614] = 12'h111;
rom[56615] = 12'h111;
rom[56616] = 12'h111;
rom[56617] = 12'h222;
rom[56618] = 12'h333;
rom[56619] = 12'h333;
rom[56620] = 12'h333;
rom[56621] = 12'h222;
rom[56622] = 12'h222;
rom[56623] = 12'h111;
rom[56624] = 12'h111;
rom[56625] = 12'h111;
rom[56626] = 12'h111;
rom[56627] = 12'h111;
rom[56628] = 12'h  0;
rom[56629] = 12'h  0;
rom[56630] = 12'h  0;
rom[56631] = 12'h  0;
rom[56632] = 12'h  0;
rom[56633] = 12'h  0;
rom[56634] = 12'h  0;
rom[56635] = 12'h  0;
rom[56636] = 12'h  0;
rom[56637] = 12'h  0;
rom[56638] = 12'h  0;
rom[56639] = 12'h  0;
rom[56640] = 12'h  0;
rom[56641] = 12'h  0;
rom[56642] = 12'h  0;
rom[56643] = 12'h  0;
rom[56644] = 12'h  0;
rom[56645] = 12'h  0;
rom[56646] = 12'h  0;
rom[56647] = 12'h  0;
rom[56648] = 12'h  0;
rom[56649] = 12'h  0;
rom[56650] = 12'h  0;
rom[56651] = 12'h  0;
rom[56652] = 12'h  0;
rom[56653] = 12'h  0;
rom[56654] = 12'h  0;
rom[56655] = 12'h  0;
rom[56656] = 12'h  0;
rom[56657] = 12'h  0;
rom[56658] = 12'h  0;
rom[56659] = 12'h  0;
rom[56660] = 12'h  0;
rom[56661] = 12'h  0;
rom[56662] = 12'h  0;
rom[56663] = 12'h  0;
rom[56664] = 12'h  0;
rom[56665] = 12'h  0;
rom[56666] = 12'h  0;
rom[56667] = 12'h  0;
rom[56668] = 12'h  0;
rom[56669] = 12'h  0;
rom[56670] = 12'h  0;
rom[56671] = 12'h  0;
rom[56672] = 12'h  0;
rom[56673] = 12'h111;
rom[56674] = 12'h111;
rom[56675] = 12'h222;
rom[56676] = 12'h222;
rom[56677] = 12'h222;
rom[56678] = 12'h333;
rom[56679] = 12'h333;
rom[56680] = 12'h333;
rom[56681] = 12'h333;
rom[56682] = 12'h444;
rom[56683] = 12'h555;
rom[56684] = 12'h555;
rom[56685] = 12'h444;
rom[56686] = 12'h333;
rom[56687] = 12'h333;
rom[56688] = 12'h333;
rom[56689] = 12'h333;
rom[56690] = 12'h333;
rom[56691] = 12'h333;
rom[56692] = 12'h333;
rom[56693] = 12'h333;
rom[56694] = 12'h444;
rom[56695] = 12'h555;
rom[56696] = 12'h666;
rom[56697] = 12'h666;
rom[56698] = 12'h666;
rom[56699] = 12'h666;
rom[56700] = 12'h555;
rom[56701] = 12'h555;
rom[56702] = 12'h555;
rom[56703] = 12'h666;
rom[56704] = 12'h666;
rom[56705] = 12'h666;
rom[56706] = 12'h555;
rom[56707] = 12'h555;
rom[56708] = 12'h555;
rom[56709] = 12'h555;
rom[56710] = 12'h555;
rom[56711] = 12'h555;
rom[56712] = 12'h555;
rom[56713] = 12'h555;
rom[56714] = 12'h555;
rom[56715] = 12'h555;
rom[56716] = 12'h555;
rom[56717] = 12'h555;
rom[56718] = 12'h555;
rom[56719] = 12'h555;
rom[56720] = 12'h555;
rom[56721] = 12'h555;
rom[56722] = 12'h555;
rom[56723] = 12'h555;
rom[56724] = 12'h555;
rom[56725] = 12'h555;
rom[56726] = 12'h555;
rom[56727] = 12'h555;
rom[56728] = 12'h555;
rom[56729] = 12'h555;
rom[56730] = 12'h555;
rom[56731] = 12'h666;
rom[56732] = 12'h666;
rom[56733] = 12'h666;
rom[56734] = 12'h666;
rom[56735] = 12'h666;
rom[56736] = 12'h666;
rom[56737] = 12'h777;
rom[56738] = 12'h777;
rom[56739] = 12'h777;
rom[56740] = 12'h777;
rom[56741] = 12'h777;
rom[56742] = 12'h888;
rom[56743] = 12'h888;
rom[56744] = 12'h888;
rom[56745] = 12'h888;
rom[56746] = 12'h888;
rom[56747] = 12'h999;
rom[56748] = 12'h999;
rom[56749] = 12'h999;
rom[56750] = 12'h999;
rom[56751] = 12'h999;
rom[56752] = 12'haaa;
rom[56753] = 12'haaa;
rom[56754] = 12'haaa;
rom[56755] = 12'haaa;
rom[56756] = 12'hbbb;
rom[56757] = 12'hbbb;
rom[56758] = 12'hbbb;
rom[56759] = 12'hccc;
rom[56760] = 12'hccc;
rom[56761] = 12'hccc;
rom[56762] = 12'hddd;
rom[56763] = 12'heee;
rom[56764] = 12'heee;
rom[56765] = 12'heee;
rom[56766] = 12'hddd;
rom[56767] = 12'hddd;
rom[56768] = 12'hccc;
rom[56769] = 12'hccc;
rom[56770] = 12'hccc;
rom[56771] = 12'hbbb;
rom[56772] = 12'hbbb;
rom[56773] = 12'hbbb;
rom[56774] = 12'hbbb;
rom[56775] = 12'hbbb;
rom[56776] = 12'hbbb;
rom[56777] = 12'haaa;
rom[56778] = 12'haaa;
rom[56779] = 12'haaa;
rom[56780] = 12'haaa;
rom[56781] = 12'haaa;
rom[56782] = 12'haaa;
rom[56783] = 12'haaa;
rom[56784] = 12'h999;
rom[56785] = 12'h999;
rom[56786] = 12'h999;
rom[56787] = 12'h999;
rom[56788] = 12'h999;
rom[56789] = 12'h999;
rom[56790] = 12'h999;
rom[56791] = 12'h999;
rom[56792] = 12'h999;
rom[56793] = 12'h999;
rom[56794] = 12'h999;
rom[56795] = 12'h999;
rom[56796] = 12'h999;
rom[56797] = 12'h999;
rom[56798] = 12'h999;
rom[56799] = 12'h999;
rom[56800] = 12'hfff;
rom[56801] = 12'hfff;
rom[56802] = 12'hfff;
rom[56803] = 12'hfff;
rom[56804] = 12'hfff;
rom[56805] = 12'hfff;
rom[56806] = 12'hfff;
rom[56807] = 12'hfff;
rom[56808] = 12'hfff;
rom[56809] = 12'hfff;
rom[56810] = 12'hfff;
rom[56811] = 12'hfff;
rom[56812] = 12'hfff;
rom[56813] = 12'hfff;
rom[56814] = 12'hfff;
rom[56815] = 12'hfff;
rom[56816] = 12'hfff;
rom[56817] = 12'hfff;
rom[56818] = 12'hfff;
rom[56819] = 12'hfff;
rom[56820] = 12'hfff;
rom[56821] = 12'hfff;
rom[56822] = 12'hfff;
rom[56823] = 12'hfff;
rom[56824] = 12'hfff;
rom[56825] = 12'hfff;
rom[56826] = 12'hfff;
rom[56827] = 12'hfff;
rom[56828] = 12'hfff;
rom[56829] = 12'hfff;
rom[56830] = 12'hfff;
rom[56831] = 12'hfff;
rom[56832] = 12'hfff;
rom[56833] = 12'hfff;
rom[56834] = 12'hfff;
rom[56835] = 12'hfff;
rom[56836] = 12'hfff;
rom[56837] = 12'hfff;
rom[56838] = 12'hfff;
rom[56839] = 12'hfff;
rom[56840] = 12'hfff;
rom[56841] = 12'hfff;
rom[56842] = 12'hfff;
rom[56843] = 12'hfff;
rom[56844] = 12'hfff;
rom[56845] = 12'hfff;
rom[56846] = 12'hfff;
rom[56847] = 12'hfff;
rom[56848] = 12'hfff;
rom[56849] = 12'hfff;
rom[56850] = 12'hfff;
rom[56851] = 12'hfff;
rom[56852] = 12'hfff;
rom[56853] = 12'hfff;
rom[56854] = 12'hfff;
rom[56855] = 12'hfff;
rom[56856] = 12'hfff;
rom[56857] = 12'hfff;
rom[56858] = 12'hfff;
rom[56859] = 12'hfff;
rom[56860] = 12'hfff;
rom[56861] = 12'hfff;
rom[56862] = 12'hfff;
rom[56863] = 12'hfff;
rom[56864] = 12'hfff;
rom[56865] = 12'hfff;
rom[56866] = 12'hfff;
rom[56867] = 12'hfff;
rom[56868] = 12'hfff;
rom[56869] = 12'hfff;
rom[56870] = 12'hfff;
rom[56871] = 12'hfff;
rom[56872] = 12'hfff;
rom[56873] = 12'hfff;
rom[56874] = 12'hfff;
rom[56875] = 12'hfff;
rom[56876] = 12'hfff;
rom[56877] = 12'hfff;
rom[56878] = 12'hfff;
rom[56879] = 12'hfff;
rom[56880] = 12'hfff;
rom[56881] = 12'hfff;
rom[56882] = 12'heee;
rom[56883] = 12'heee;
rom[56884] = 12'heee;
rom[56885] = 12'hddd;
rom[56886] = 12'hddd;
rom[56887] = 12'hddd;
rom[56888] = 12'hccc;
rom[56889] = 12'hccc;
rom[56890] = 12'hccc;
rom[56891] = 12'hccc;
rom[56892] = 12'hccc;
rom[56893] = 12'hddd;
rom[56894] = 12'hccc;
rom[56895] = 12'hccc;
rom[56896] = 12'hddd;
rom[56897] = 12'hddd;
rom[56898] = 12'hddd;
rom[56899] = 12'hddd;
rom[56900] = 12'hddd;
rom[56901] = 12'hccc;
rom[56902] = 12'hccc;
rom[56903] = 12'hbbb;
rom[56904] = 12'haaa;
rom[56905] = 12'haaa;
rom[56906] = 12'haaa;
rom[56907] = 12'haaa;
rom[56908] = 12'haaa;
rom[56909] = 12'haaa;
rom[56910] = 12'haaa;
rom[56911] = 12'haaa;
rom[56912] = 12'haaa;
rom[56913] = 12'h999;
rom[56914] = 12'h999;
rom[56915] = 12'h888;
rom[56916] = 12'h888;
rom[56917] = 12'h777;
rom[56918] = 12'h777;
rom[56919] = 12'h777;
rom[56920] = 12'h777;
rom[56921] = 12'h777;
rom[56922] = 12'h777;
rom[56923] = 12'h777;
rom[56924] = 12'h888;
rom[56925] = 12'h999;
rom[56926] = 12'h999;
rom[56927] = 12'haaa;
rom[56928] = 12'haaa;
rom[56929] = 12'haaa;
rom[56930] = 12'h999;
rom[56931] = 12'h888;
rom[56932] = 12'h777;
rom[56933] = 12'h666;
rom[56934] = 12'h666;
rom[56935] = 12'h555;
rom[56936] = 12'h555;
rom[56937] = 12'h555;
rom[56938] = 12'h555;
rom[56939] = 12'h555;
rom[56940] = 12'h555;
rom[56941] = 12'h555;
rom[56942] = 12'h444;
rom[56943] = 12'h444;
rom[56944] = 12'h444;
rom[56945] = 12'h444;
rom[56946] = 12'h333;
rom[56947] = 12'h333;
rom[56948] = 12'h333;
rom[56949] = 12'h222;
rom[56950] = 12'h222;
rom[56951] = 12'h222;
rom[56952] = 12'h222;
rom[56953] = 12'h222;
rom[56954] = 12'h222;
rom[56955] = 12'h222;
rom[56956] = 12'h222;
rom[56957] = 12'h222;
rom[56958] = 12'h111;
rom[56959] = 12'h111;
rom[56960] = 12'h111;
rom[56961] = 12'h111;
rom[56962] = 12'h111;
rom[56963] = 12'h111;
rom[56964] = 12'h111;
rom[56965] = 12'h111;
rom[56966] = 12'h111;
rom[56967] = 12'h111;
rom[56968] = 12'h111;
rom[56969] = 12'h111;
rom[56970] = 12'h111;
rom[56971] = 12'h111;
rom[56972] = 12'h111;
rom[56973] = 12'h  0;
rom[56974] = 12'h  0;
rom[56975] = 12'h  0;
rom[56976] = 12'h  0;
rom[56977] = 12'h  0;
rom[56978] = 12'h  0;
rom[56979] = 12'h  0;
rom[56980] = 12'h  0;
rom[56981] = 12'h  0;
rom[56982] = 12'h  0;
rom[56983] = 12'h  0;
rom[56984] = 12'h  0;
rom[56985] = 12'h  0;
rom[56986] = 12'h  0;
rom[56987] = 12'h  0;
rom[56988] = 12'h  0;
rom[56989] = 12'h  0;
rom[56990] = 12'h  0;
rom[56991] = 12'h  0;
rom[56992] = 12'h  0;
rom[56993] = 12'h  0;
rom[56994] = 12'h  0;
rom[56995] = 12'h  0;
rom[56996] = 12'h  0;
rom[56997] = 12'h  0;
rom[56998] = 12'h  0;
rom[56999] = 12'h  0;
rom[57000] = 12'h  0;
rom[57001] = 12'h  0;
rom[57002] = 12'h  0;
rom[57003] = 12'h  0;
rom[57004] = 12'h111;
rom[57005] = 12'h111;
rom[57006] = 12'h111;
rom[57007] = 12'h111;
rom[57008] = 12'h111;
rom[57009] = 12'h111;
rom[57010] = 12'h  0;
rom[57011] = 12'h  0;
rom[57012] = 12'h111;
rom[57013] = 12'h111;
rom[57014] = 12'h111;
rom[57015] = 12'h111;
rom[57016] = 12'h222;
rom[57017] = 12'h222;
rom[57018] = 12'h333;
rom[57019] = 12'h333;
rom[57020] = 12'h333;
rom[57021] = 12'h222;
rom[57022] = 12'h111;
rom[57023] = 12'h111;
rom[57024] = 12'h111;
rom[57025] = 12'h111;
rom[57026] = 12'h111;
rom[57027] = 12'h  0;
rom[57028] = 12'h  0;
rom[57029] = 12'h  0;
rom[57030] = 12'h  0;
rom[57031] = 12'h  0;
rom[57032] = 12'h  0;
rom[57033] = 12'h  0;
rom[57034] = 12'h  0;
rom[57035] = 12'h  0;
rom[57036] = 12'h  0;
rom[57037] = 12'h  0;
rom[57038] = 12'h  0;
rom[57039] = 12'h  0;
rom[57040] = 12'h  0;
rom[57041] = 12'h  0;
rom[57042] = 12'h  0;
rom[57043] = 12'h  0;
rom[57044] = 12'h  0;
rom[57045] = 12'h  0;
rom[57046] = 12'h  0;
rom[57047] = 12'h  0;
rom[57048] = 12'h  0;
rom[57049] = 12'h  0;
rom[57050] = 12'h  0;
rom[57051] = 12'h  0;
rom[57052] = 12'h  0;
rom[57053] = 12'h  0;
rom[57054] = 12'h  0;
rom[57055] = 12'h  0;
rom[57056] = 12'h  0;
rom[57057] = 12'h  0;
rom[57058] = 12'h  0;
rom[57059] = 12'h  0;
rom[57060] = 12'h  0;
rom[57061] = 12'h  0;
rom[57062] = 12'h  0;
rom[57063] = 12'h  0;
rom[57064] = 12'h  0;
rom[57065] = 12'h  0;
rom[57066] = 12'h  0;
rom[57067] = 12'h  0;
rom[57068] = 12'h  0;
rom[57069] = 12'h  0;
rom[57070] = 12'h  0;
rom[57071] = 12'h  0;
rom[57072] = 12'h  0;
rom[57073] = 12'h111;
rom[57074] = 12'h111;
rom[57075] = 12'h222;
rom[57076] = 12'h222;
rom[57077] = 12'h222;
rom[57078] = 12'h222;
rom[57079] = 12'h333;
rom[57080] = 12'h333;
rom[57081] = 12'h333;
rom[57082] = 12'h444;
rom[57083] = 12'h555;
rom[57084] = 12'h555;
rom[57085] = 12'h444;
rom[57086] = 12'h333;
rom[57087] = 12'h222;
rom[57088] = 12'h333;
rom[57089] = 12'h333;
rom[57090] = 12'h333;
rom[57091] = 12'h333;
rom[57092] = 12'h333;
rom[57093] = 12'h333;
rom[57094] = 12'h444;
rom[57095] = 12'h555;
rom[57096] = 12'h666;
rom[57097] = 12'h666;
rom[57098] = 12'h666;
rom[57099] = 12'h666;
rom[57100] = 12'h555;
rom[57101] = 12'h555;
rom[57102] = 12'h555;
rom[57103] = 12'h555;
rom[57104] = 12'h666;
rom[57105] = 12'h666;
rom[57106] = 12'h666;
rom[57107] = 12'h555;
rom[57108] = 12'h555;
rom[57109] = 12'h555;
rom[57110] = 12'h555;
rom[57111] = 12'h555;
rom[57112] = 12'h555;
rom[57113] = 12'h555;
rom[57114] = 12'h555;
rom[57115] = 12'h555;
rom[57116] = 12'h555;
rom[57117] = 12'h555;
rom[57118] = 12'h555;
rom[57119] = 12'h555;
rom[57120] = 12'h555;
rom[57121] = 12'h555;
rom[57122] = 12'h555;
rom[57123] = 12'h555;
rom[57124] = 12'h555;
rom[57125] = 12'h555;
rom[57126] = 12'h555;
rom[57127] = 12'h666;
rom[57128] = 12'h555;
rom[57129] = 12'h666;
rom[57130] = 12'h666;
rom[57131] = 12'h666;
rom[57132] = 12'h666;
rom[57133] = 12'h666;
rom[57134] = 12'h666;
rom[57135] = 12'h666;
rom[57136] = 12'h666;
rom[57137] = 12'h777;
rom[57138] = 12'h777;
rom[57139] = 12'h777;
rom[57140] = 12'h777;
rom[57141] = 12'h777;
rom[57142] = 12'h888;
rom[57143] = 12'h888;
rom[57144] = 12'h888;
rom[57145] = 12'h888;
rom[57146] = 12'h999;
rom[57147] = 12'h999;
rom[57148] = 12'h999;
rom[57149] = 12'h999;
rom[57150] = 12'h999;
rom[57151] = 12'h999;
rom[57152] = 12'haaa;
rom[57153] = 12'haaa;
rom[57154] = 12'haaa;
rom[57155] = 12'hbbb;
rom[57156] = 12'hbbb;
rom[57157] = 12'hbbb;
rom[57158] = 12'hccc;
rom[57159] = 12'hccc;
rom[57160] = 12'hddd;
rom[57161] = 12'hddd;
rom[57162] = 12'heee;
rom[57163] = 12'heee;
rom[57164] = 12'heee;
rom[57165] = 12'hddd;
rom[57166] = 12'hddd;
rom[57167] = 12'hccc;
rom[57168] = 12'hccc;
rom[57169] = 12'hccc;
rom[57170] = 12'hbbb;
rom[57171] = 12'hbbb;
rom[57172] = 12'hbbb;
rom[57173] = 12'hbbb;
rom[57174] = 12'hbbb;
rom[57175] = 12'hbbb;
rom[57176] = 12'haaa;
rom[57177] = 12'haaa;
rom[57178] = 12'haaa;
rom[57179] = 12'haaa;
rom[57180] = 12'haaa;
rom[57181] = 12'haaa;
rom[57182] = 12'haaa;
rom[57183] = 12'h999;
rom[57184] = 12'h999;
rom[57185] = 12'h999;
rom[57186] = 12'h999;
rom[57187] = 12'h999;
rom[57188] = 12'h999;
rom[57189] = 12'h999;
rom[57190] = 12'h999;
rom[57191] = 12'h999;
rom[57192] = 12'h999;
rom[57193] = 12'h999;
rom[57194] = 12'h999;
rom[57195] = 12'h999;
rom[57196] = 12'h999;
rom[57197] = 12'h999;
rom[57198] = 12'h999;
rom[57199] = 12'h999;
rom[57200] = 12'hfff;
rom[57201] = 12'hfff;
rom[57202] = 12'hfff;
rom[57203] = 12'hfff;
rom[57204] = 12'hfff;
rom[57205] = 12'hfff;
rom[57206] = 12'hfff;
rom[57207] = 12'hfff;
rom[57208] = 12'hfff;
rom[57209] = 12'hfff;
rom[57210] = 12'hfff;
rom[57211] = 12'hfff;
rom[57212] = 12'hfff;
rom[57213] = 12'hfff;
rom[57214] = 12'hfff;
rom[57215] = 12'hfff;
rom[57216] = 12'hfff;
rom[57217] = 12'hfff;
rom[57218] = 12'hfff;
rom[57219] = 12'hfff;
rom[57220] = 12'hfff;
rom[57221] = 12'hfff;
rom[57222] = 12'hfff;
rom[57223] = 12'hfff;
rom[57224] = 12'hfff;
rom[57225] = 12'hfff;
rom[57226] = 12'hfff;
rom[57227] = 12'hfff;
rom[57228] = 12'hfff;
rom[57229] = 12'hfff;
rom[57230] = 12'hfff;
rom[57231] = 12'hfff;
rom[57232] = 12'hfff;
rom[57233] = 12'hfff;
rom[57234] = 12'hfff;
rom[57235] = 12'hfff;
rom[57236] = 12'hfff;
rom[57237] = 12'hfff;
rom[57238] = 12'hfff;
rom[57239] = 12'hfff;
rom[57240] = 12'hfff;
rom[57241] = 12'hfff;
rom[57242] = 12'hfff;
rom[57243] = 12'hfff;
rom[57244] = 12'hfff;
rom[57245] = 12'hfff;
rom[57246] = 12'hfff;
rom[57247] = 12'hfff;
rom[57248] = 12'hfff;
rom[57249] = 12'hfff;
rom[57250] = 12'hfff;
rom[57251] = 12'hfff;
rom[57252] = 12'hfff;
rom[57253] = 12'hfff;
rom[57254] = 12'hfff;
rom[57255] = 12'hfff;
rom[57256] = 12'hfff;
rom[57257] = 12'hfff;
rom[57258] = 12'hfff;
rom[57259] = 12'hfff;
rom[57260] = 12'hfff;
rom[57261] = 12'hfff;
rom[57262] = 12'hfff;
rom[57263] = 12'hfff;
rom[57264] = 12'hfff;
rom[57265] = 12'hfff;
rom[57266] = 12'hfff;
rom[57267] = 12'hfff;
rom[57268] = 12'hfff;
rom[57269] = 12'hfff;
rom[57270] = 12'hfff;
rom[57271] = 12'hfff;
rom[57272] = 12'hfff;
rom[57273] = 12'hfff;
rom[57274] = 12'hfff;
rom[57275] = 12'hfff;
rom[57276] = 12'hfff;
rom[57277] = 12'hfff;
rom[57278] = 12'hfff;
rom[57279] = 12'hfff;
rom[57280] = 12'hfff;
rom[57281] = 12'hfff;
rom[57282] = 12'hfff;
rom[57283] = 12'hfff;
rom[57284] = 12'heee;
rom[57285] = 12'heee;
rom[57286] = 12'hddd;
rom[57287] = 12'hccc;
rom[57288] = 12'hccc;
rom[57289] = 12'hccc;
rom[57290] = 12'hccc;
rom[57291] = 12'hccc;
rom[57292] = 12'hccc;
rom[57293] = 12'hccc;
rom[57294] = 12'hccc;
rom[57295] = 12'hccc;
rom[57296] = 12'hccc;
rom[57297] = 12'hccc;
rom[57298] = 12'hddd;
rom[57299] = 12'heee;
rom[57300] = 12'heee;
rom[57301] = 12'heee;
rom[57302] = 12'hddd;
rom[57303] = 12'hccc;
rom[57304] = 12'hbbb;
rom[57305] = 12'hbbb;
rom[57306] = 12'hbbb;
rom[57307] = 12'haaa;
rom[57308] = 12'haaa;
rom[57309] = 12'haaa;
rom[57310] = 12'haaa;
rom[57311] = 12'haaa;
rom[57312] = 12'haaa;
rom[57313] = 12'haaa;
rom[57314] = 12'haaa;
rom[57315] = 12'h999;
rom[57316] = 12'h999;
rom[57317] = 12'h888;
rom[57318] = 12'h888;
rom[57319] = 12'h888;
rom[57320] = 12'h777;
rom[57321] = 12'h777;
rom[57322] = 12'h777;
rom[57323] = 12'h777;
rom[57324] = 12'h777;
rom[57325] = 12'h777;
rom[57326] = 12'h888;
rom[57327] = 12'h888;
rom[57328] = 12'h999;
rom[57329] = 12'h999;
rom[57330] = 12'h999;
rom[57331] = 12'h888;
rom[57332] = 12'h888;
rom[57333] = 12'h777;
rom[57334] = 12'h666;
rom[57335] = 12'h555;
rom[57336] = 12'h555;
rom[57337] = 12'h555;
rom[57338] = 12'h555;
rom[57339] = 12'h555;
rom[57340] = 12'h555;
rom[57341] = 12'h444;
rom[57342] = 12'h444;
rom[57343] = 12'h444;
rom[57344] = 12'h444;
rom[57345] = 12'h333;
rom[57346] = 12'h333;
rom[57347] = 12'h333;
rom[57348] = 12'h222;
rom[57349] = 12'h222;
rom[57350] = 12'h222;
rom[57351] = 12'h222;
rom[57352] = 12'h222;
rom[57353] = 12'h222;
rom[57354] = 12'h222;
rom[57355] = 12'h222;
rom[57356] = 12'h222;
rom[57357] = 12'h111;
rom[57358] = 12'h111;
rom[57359] = 12'h111;
rom[57360] = 12'h111;
rom[57361] = 12'h111;
rom[57362] = 12'h111;
rom[57363] = 12'h111;
rom[57364] = 12'h111;
rom[57365] = 12'h111;
rom[57366] = 12'h111;
rom[57367] = 12'h111;
rom[57368] = 12'h111;
rom[57369] = 12'h111;
rom[57370] = 12'h111;
rom[57371] = 12'h111;
rom[57372] = 12'h  0;
rom[57373] = 12'h  0;
rom[57374] = 12'h  0;
rom[57375] = 12'h  0;
rom[57376] = 12'h  0;
rom[57377] = 12'h  0;
rom[57378] = 12'h111;
rom[57379] = 12'h111;
rom[57380] = 12'h111;
rom[57381] = 12'h111;
rom[57382] = 12'h  0;
rom[57383] = 12'h  0;
rom[57384] = 12'h  0;
rom[57385] = 12'h  0;
rom[57386] = 12'h  0;
rom[57387] = 12'h  0;
rom[57388] = 12'h  0;
rom[57389] = 12'h  0;
rom[57390] = 12'h  0;
rom[57391] = 12'h  0;
rom[57392] = 12'h  0;
rom[57393] = 12'h  0;
rom[57394] = 12'h  0;
rom[57395] = 12'h  0;
rom[57396] = 12'h  0;
rom[57397] = 12'h  0;
rom[57398] = 12'h  0;
rom[57399] = 12'h  0;
rom[57400] = 12'h  0;
rom[57401] = 12'h  0;
rom[57402] = 12'h  0;
rom[57403] = 12'h  0;
rom[57404] = 12'h111;
rom[57405] = 12'h111;
rom[57406] = 12'h111;
rom[57407] = 12'h111;
rom[57408] = 12'h111;
rom[57409] = 12'h111;
rom[57410] = 12'h  0;
rom[57411] = 12'h111;
rom[57412] = 12'h111;
rom[57413] = 12'h111;
rom[57414] = 12'h111;
rom[57415] = 12'h111;
rom[57416] = 12'h222;
rom[57417] = 12'h222;
rom[57418] = 12'h333;
rom[57419] = 12'h333;
rom[57420] = 12'h333;
rom[57421] = 12'h222;
rom[57422] = 12'h111;
rom[57423] = 12'h222;
rom[57424] = 12'h111;
rom[57425] = 12'h111;
rom[57426] = 12'h111;
rom[57427] = 12'h  0;
rom[57428] = 12'h  0;
rom[57429] = 12'h  0;
rom[57430] = 12'h  0;
rom[57431] = 12'h  0;
rom[57432] = 12'h  0;
rom[57433] = 12'h  0;
rom[57434] = 12'h  0;
rom[57435] = 12'h  0;
rom[57436] = 12'h  0;
rom[57437] = 12'h  0;
rom[57438] = 12'h  0;
rom[57439] = 12'h  0;
rom[57440] = 12'h  0;
rom[57441] = 12'h  0;
rom[57442] = 12'h  0;
rom[57443] = 12'h  0;
rom[57444] = 12'h  0;
rom[57445] = 12'h  0;
rom[57446] = 12'h  0;
rom[57447] = 12'h  0;
rom[57448] = 12'h  0;
rom[57449] = 12'h  0;
rom[57450] = 12'h  0;
rom[57451] = 12'h  0;
rom[57452] = 12'h  0;
rom[57453] = 12'h  0;
rom[57454] = 12'h  0;
rom[57455] = 12'h  0;
rom[57456] = 12'h  0;
rom[57457] = 12'h  0;
rom[57458] = 12'h  0;
rom[57459] = 12'h  0;
rom[57460] = 12'h  0;
rom[57461] = 12'h  0;
rom[57462] = 12'h  0;
rom[57463] = 12'h  0;
rom[57464] = 12'h  0;
rom[57465] = 12'h  0;
rom[57466] = 12'h  0;
rom[57467] = 12'h  0;
rom[57468] = 12'h  0;
rom[57469] = 12'h  0;
rom[57470] = 12'h  0;
rom[57471] = 12'h  0;
rom[57472] = 12'h  0;
rom[57473] = 12'h111;
rom[57474] = 12'h111;
rom[57475] = 12'h222;
rom[57476] = 12'h222;
rom[57477] = 12'h222;
rom[57478] = 12'h222;
rom[57479] = 12'h333;
rom[57480] = 12'h333;
rom[57481] = 12'h333;
rom[57482] = 12'h444;
rom[57483] = 12'h555;
rom[57484] = 12'h555;
rom[57485] = 12'h444;
rom[57486] = 12'h333;
rom[57487] = 12'h222;
rom[57488] = 12'h222;
rom[57489] = 12'h222;
rom[57490] = 12'h333;
rom[57491] = 12'h333;
rom[57492] = 12'h333;
rom[57493] = 12'h333;
rom[57494] = 12'h444;
rom[57495] = 12'h555;
rom[57496] = 12'h666;
rom[57497] = 12'h666;
rom[57498] = 12'h666;
rom[57499] = 12'h666;
rom[57500] = 12'h666;
rom[57501] = 12'h555;
rom[57502] = 12'h555;
rom[57503] = 12'h555;
rom[57504] = 12'h666;
rom[57505] = 12'h666;
rom[57506] = 12'h666;
rom[57507] = 12'h555;
rom[57508] = 12'h555;
rom[57509] = 12'h555;
rom[57510] = 12'h555;
rom[57511] = 12'h555;
rom[57512] = 12'h555;
rom[57513] = 12'h555;
rom[57514] = 12'h555;
rom[57515] = 12'h666;
rom[57516] = 12'h666;
rom[57517] = 12'h555;
rom[57518] = 12'h555;
rom[57519] = 12'h555;
rom[57520] = 12'h555;
rom[57521] = 12'h555;
rom[57522] = 12'h555;
rom[57523] = 12'h555;
rom[57524] = 12'h555;
rom[57525] = 12'h666;
rom[57526] = 12'h666;
rom[57527] = 12'h666;
rom[57528] = 12'h666;
rom[57529] = 12'h666;
rom[57530] = 12'h666;
rom[57531] = 12'h666;
rom[57532] = 12'h666;
rom[57533] = 12'h666;
rom[57534] = 12'h666;
rom[57535] = 12'h777;
rom[57536] = 12'h777;
rom[57537] = 12'h777;
rom[57538] = 12'h777;
rom[57539] = 12'h777;
rom[57540] = 12'h777;
rom[57541] = 12'h888;
rom[57542] = 12'h888;
rom[57543] = 12'h888;
rom[57544] = 12'h888;
rom[57545] = 12'h999;
rom[57546] = 12'h999;
rom[57547] = 12'h999;
rom[57548] = 12'h999;
rom[57549] = 12'h999;
rom[57550] = 12'h999;
rom[57551] = 12'haaa;
rom[57552] = 12'haaa;
rom[57553] = 12'haaa;
rom[57554] = 12'hbbb;
rom[57555] = 12'hbbb;
rom[57556] = 12'hbbb;
rom[57557] = 12'hccc;
rom[57558] = 12'hccc;
rom[57559] = 12'hccc;
rom[57560] = 12'hddd;
rom[57561] = 12'heee;
rom[57562] = 12'heee;
rom[57563] = 12'heee;
rom[57564] = 12'heee;
rom[57565] = 12'hddd;
rom[57566] = 12'hccc;
rom[57567] = 12'hccc;
rom[57568] = 12'hccc;
rom[57569] = 12'hccc;
rom[57570] = 12'hbbb;
rom[57571] = 12'hbbb;
rom[57572] = 12'hbbb;
rom[57573] = 12'hbbb;
rom[57574] = 12'haaa;
rom[57575] = 12'haaa;
rom[57576] = 12'haaa;
rom[57577] = 12'haaa;
rom[57578] = 12'haaa;
rom[57579] = 12'haaa;
rom[57580] = 12'haaa;
rom[57581] = 12'haaa;
rom[57582] = 12'h999;
rom[57583] = 12'h999;
rom[57584] = 12'h999;
rom[57585] = 12'h999;
rom[57586] = 12'h999;
rom[57587] = 12'h999;
rom[57588] = 12'h999;
rom[57589] = 12'h999;
rom[57590] = 12'h999;
rom[57591] = 12'h999;
rom[57592] = 12'h999;
rom[57593] = 12'h999;
rom[57594] = 12'h999;
rom[57595] = 12'h999;
rom[57596] = 12'h999;
rom[57597] = 12'h999;
rom[57598] = 12'h999;
rom[57599] = 12'h999;
rom[57600] = 12'hfff;
rom[57601] = 12'hfff;
rom[57602] = 12'hfff;
rom[57603] = 12'hfff;
rom[57604] = 12'hfff;
rom[57605] = 12'hfff;
rom[57606] = 12'hfff;
rom[57607] = 12'hfff;
rom[57608] = 12'hfff;
rom[57609] = 12'hfff;
rom[57610] = 12'hfff;
rom[57611] = 12'hfff;
rom[57612] = 12'hfff;
rom[57613] = 12'hfff;
rom[57614] = 12'hfff;
rom[57615] = 12'hfff;
rom[57616] = 12'hfff;
rom[57617] = 12'hfff;
rom[57618] = 12'hfff;
rom[57619] = 12'hfff;
rom[57620] = 12'hfff;
rom[57621] = 12'hfff;
rom[57622] = 12'hfff;
rom[57623] = 12'hfff;
rom[57624] = 12'hfff;
rom[57625] = 12'hfff;
rom[57626] = 12'hfff;
rom[57627] = 12'hfff;
rom[57628] = 12'hfff;
rom[57629] = 12'hfff;
rom[57630] = 12'hfff;
rom[57631] = 12'hfff;
rom[57632] = 12'hfff;
rom[57633] = 12'hfff;
rom[57634] = 12'hfff;
rom[57635] = 12'hfff;
rom[57636] = 12'hfff;
rom[57637] = 12'hfff;
rom[57638] = 12'hfff;
rom[57639] = 12'hfff;
rom[57640] = 12'hfff;
rom[57641] = 12'hfff;
rom[57642] = 12'hfff;
rom[57643] = 12'hfff;
rom[57644] = 12'hfff;
rom[57645] = 12'hfff;
rom[57646] = 12'hfff;
rom[57647] = 12'hfff;
rom[57648] = 12'hfff;
rom[57649] = 12'hfff;
rom[57650] = 12'hfff;
rom[57651] = 12'hfff;
rom[57652] = 12'hfff;
rom[57653] = 12'hfff;
rom[57654] = 12'hfff;
rom[57655] = 12'hfff;
rom[57656] = 12'hfff;
rom[57657] = 12'hfff;
rom[57658] = 12'hfff;
rom[57659] = 12'hfff;
rom[57660] = 12'hfff;
rom[57661] = 12'hfff;
rom[57662] = 12'hfff;
rom[57663] = 12'hfff;
rom[57664] = 12'hfff;
rom[57665] = 12'hfff;
rom[57666] = 12'hfff;
rom[57667] = 12'hfff;
rom[57668] = 12'hfff;
rom[57669] = 12'hfff;
rom[57670] = 12'hfff;
rom[57671] = 12'hfff;
rom[57672] = 12'hfff;
rom[57673] = 12'hfff;
rom[57674] = 12'hfff;
rom[57675] = 12'hfff;
rom[57676] = 12'hfff;
rom[57677] = 12'hfff;
rom[57678] = 12'hfff;
rom[57679] = 12'hfff;
rom[57680] = 12'hfff;
rom[57681] = 12'hfff;
rom[57682] = 12'hfff;
rom[57683] = 12'hfff;
rom[57684] = 12'hfff;
rom[57685] = 12'heee;
rom[57686] = 12'heee;
rom[57687] = 12'hddd;
rom[57688] = 12'hddd;
rom[57689] = 12'hddd;
rom[57690] = 12'hddd;
rom[57691] = 12'hccc;
rom[57692] = 12'hccc;
rom[57693] = 12'hccc;
rom[57694] = 12'hccc;
rom[57695] = 12'hccc;
rom[57696] = 12'hbbb;
rom[57697] = 12'hbbb;
rom[57698] = 12'hccc;
rom[57699] = 12'hccc;
rom[57700] = 12'hccc;
rom[57701] = 12'hddd;
rom[57702] = 12'hddd;
rom[57703] = 12'hddd;
rom[57704] = 12'heee;
rom[57705] = 12'hddd;
rom[57706] = 12'hddd;
rom[57707] = 12'hddd;
rom[57708] = 12'hccc;
rom[57709] = 12'hbbb;
rom[57710] = 12'haaa;
rom[57711] = 12'haaa;
rom[57712] = 12'haaa;
rom[57713] = 12'haaa;
rom[57714] = 12'haaa;
rom[57715] = 12'haaa;
rom[57716] = 12'h999;
rom[57717] = 12'h999;
rom[57718] = 12'h888;
rom[57719] = 12'h888;
rom[57720] = 12'h888;
rom[57721] = 12'h888;
rom[57722] = 12'h888;
rom[57723] = 12'h888;
rom[57724] = 12'h888;
rom[57725] = 12'h888;
rom[57726] = 12'h888;
rom[57727] = 12'h777;
rom[57728] = 12'h999;
rom[57729] = 12'h888;
rom[57730] = 12'h888;
rom[57731] = 12'h888;
rom[57732] = 12'h888;
rom[57733] = 12'h777;
rom[57734] = 12'h777;
rom[57735] = 12'h666;
rom[57736] = 12'h666;
rom[57737] = 12'h666;
rom[57738] = 12'h555;
rom[57739] = 12'h555;
rom[57740] = 12'h555;
rom[57741] = 12'h444;
rom[57742] = 12'h444;
rom[57743] = 12'h333;
rom[57744] = 12'h333;
rom[57745] = 12'h333;
rom[57746] = 12'h333;
rom[57747] = 12'h222;
rom[57748] = 12'h222;
rom[57749] = 12'h222;
rom[57750] = 12'h222;
rom[57751] = 12'h222;
rom[57752] = 12'h222;
rom[57753] = 12'h222;
rom[57754] = 12'h222;
rom[57755] = 12'h222;
rom[57756] = 12'h222;
rom[57757] = 12'h222;
rom[57758] = 12'h222;
rom[57759] = 12'h111;
rom[57760] = 12'h111;
rom[57761] = 12'h111;
rom[57762] = 12'h111;
rom[57763] = 12'h111;
rom[57764] = 12'h111;
rom[57765] = 12'h111;
rom[57766] = 12'h111;
rom[57767] = 12'h111;
rom[57768] = 12'h111;
rom[57769] = 12'h111;
rom[57770] = 12'h111;
rom[57771] = 12'h111;
rom[57772] = 12'h111;
rom[57773] = 12'h111;
rom[57774] = 12'h111;
rom[57775] = 12'h111;
rom[57776] = 12'h111;
rom[57777] = 12'h111;
rom[57778] = 12'h111;
rom[57779] = 12'h111;
rom[57780] = 12'h111;
rom[57781] = 12'h111;
rom[57782] = 12'h  0;
rom[57783] = 12'h  0;
rom[57784] = 12'h  0;
rom[57785] = 12'h  0;
rom[57786] = 12'h  0;
rom[57787] = 12'h  0;
rom[57788] = 12'h  0;
rom[57789] = 12'h  0;
rom[57790] = 12'h  0;
rom[57791] = 12'h  0;
rom[57792] = 12'h  0;
rom[57793] = 12'h  0;
rom[57794] = 12'h  0;
rom[57795] = 12'h  0;
rom[57796] = 12'h  0;
rom[57797] = 12'h  0;
rom[57798] = 12'h  0;
rom[57799] = 12'h  0;
rom[57800] = 12'h  0;
rom[57801] = 12'h  0;
rom[57802] = 12'h  0;
rom[57803] = 12'h111;
rom[57804] = 12'h111;
rom[57805] = 12'h111;
rom[57806] = 12'h111;
rom[57807] = 12'h111;
rom[57808] = 12'h111;
rom[57809] = 12'h  0;
rom[57810] = 12'h  0;
rom[57811] = 12'h111;
rom[57812] = 12'h111;
rom[57813] = 12'h111;
rom[57814] = 12'h111;
rom[57815] = 12'h222;
rom[57816] = 12'h222;
rom[57817] = 12'h333;
rom[57818] = 12'h333;
rom[57819] = 12'h333;
rom[57820] = 12'h222;
rom[57821] = 12'h111;
rom[57822] = 12'h111;
rom[57823] = 12'h111;
rom[57824] = 12'h111;
rom[57825] = 12'h111;
rom[57826] = 12'h  0;
rom[57827] = 12'h  0;
rom[57828] = 12'h  0;
rom[57829] = 12'h  0;
rom[57830] = 12'h  0;
rom[57831] = 12'h  0;
rom[57832] = 12'h  0;
rom[57833] = 12'h  0;
rom[57834] = 12'h  0;
rom[57835] = 12'h  0;
rom[57836] = 12'h  0;
rom[57837] = 12'h  0;
rom[57838] = 12'h  0;
rom[57839] = 12'h  0;
rom[57840] = 12'h  0;
rom[57841] = 12'h  0;
rom[57842] = 12'h  0;
rom[57843] = 12'h  0;
rom[57844] = 12'h  0;
rom[57845] = 12'h  0;
rom[57846] = 12'h  0;
rom[57847] = 12'h  0;
rom[57848] = 12'h  0;
rom[57849] = 12'h  0;
rom[57850] = 12'h  0;
rom[57851] = 12'h  0;
rom[57852] = 12'h  0;
rom[57853] = 12'h  0;
rom[57854] = 12'h  0;
rom[57855] = 12'h  0;
rom[57856] = 12'h  0;
rom[57857] = 12'h  0;
rom[57858] = 12'h  0;
rom[57859] = 12'h  0;
rom[57860] = 12'h  0;
rom[57861] = 12'h  0;
rom[57862] = 12'h  0;
rom[57863] = 12'h  0;
rom[57864] = 12'h  0;
rom[57865] = 12'h  0;
rom[57866] = 12'h  0;
rom[57867] = 12'h  0;
rom[57868] = 12'h  0;
rom[57869] = 12'h  0;
rom[57870] = 12'h  0;
rom[57871] = 12'h  0;
rom[57872] = 12'h  0;
rom[57873] = 12'h111;
rom[57874] = 12'h111;
rom[57875] = 12'h222;
rom[57876] = 12'h222;
rom[57877] = 12'h222;
rom[57878] = 12'h333;
rom[57879] = 12'h333;
rom[57880] = 12'h333;
rom[57881] = 12'h444;
rom[57882] = 12'h444;
rom[57883] = 12'h555;
rom[57884] = 12'h444;
rom[57885] = 12'h333;
rom[57886] = 12'h222;
rom[57887] = 12'h222;
rom[57888] = 12'h222;
rom[57889] = 12'h222;
rom[57890] = 12'h333;
rom[57891] = 12'h333;
rom[57892] = 12'h333;
rom[57893] = 12'h333;
rom[57894] = 12'h444;
rom[57895] = 12'h444;
rom[57896] = 12'h555;
rom[57897] = 12'h666;
rom[57898] = 12'h666;
rom[57899] = 12'h666;
rom[57900] = 12'h666;
rom[57901] = 12'h555;
rom[57902] = 12'h555;
rom[57903] = 12'h555;
rom[57904] = 12'h666;
rom[57905] = 12'h666;
rom[57906] = 12'h666;
rom[57907] = 12'h666;
rom[57908] = 12'h555;
rom[57909] = 12'h555;
rom[57910] = 12'h555;
rom[57911] = 12'h555;
rom[57912] = 12'h555;
rom[57913] = 12'h555;
rom[57914] = 12'h555;
rom[57915] = 12'h555;
rom[57916] = 12'h666;
rom[57917] = 12'h666;
rom[57918] = 12'h666;
rom[57919] = 12'h666;
rom[57920] = 12'h555;
rom[57921] = 12'h555;
rom[57922] = 12'h555;
rom[57923] = 12'h666;
rom[57924] = 12'h666;
rom[57925] = 12'h666;
rom[57926] = 12'h666;
rom[57927] = 12'h666;
rom[57928] = 12'h666;
rom[57929] = 12'h666;
rom[57930] = 12'h666;
rom[57931] = 12'h666;
rom[57932] = 12'h666;
rom[57933] = 12'h666;
rom[57934] = 12'h666;
rom[57935] = 12'h777;
rom[57936] = 12'h777;
rom[57937] = 12'h777;
rom[57938] = 12'h777;
rom[57939] = 12'h777;
rom[57940] = 12'h888;
rom[57941] = 12'h888;
rom[57942] = 12'h888;
rom[57943] = 12'h888;
rom[57944] = 12'h888;
rom[57945] = 12'h999;
rom[57946] = 12'h999;
rom[57947] = 12'h999;
rom[57948] = 12'h999;
rom[57949] = 12'h999;
rom[57950] = 12'haaa;
rom[57951] = 12'haaa;
rom[57952] = 12'haaa;
rom[57953] = 12'haaa;
rom[57954] = 12'hbbb;
rom[57955] = 12'hbbb;
rom[57956] = 12'hbbb;
rom[57957] = 12'hccc;
rom[57958] = 12'hddd;
rom[57959] = 12'hddd;
rom[57960] = 12'hddd;
rom[57961] = 12'heee;
rom[57962] = 12'heee;
rom[57963] = 12'heee;
rom[57964] = 12'hddd;
rom[57965] = 12'hddd;
rom[57966] = 12'hccc;
rom[57967] = 12'hccc;
rom[57968] = 12'hccc;
rom[57969] = 12'hbbb;
rom[57970] = 12'hbbb;
rom[57971] = 12'hbbb;
rom[57972] = 12'hbbb;
rom[57973] = 12'hbbb;
rom[57974] = 12'haaa;
rom[57975] = 12'haaa;
rom[57976] = 12'haaa;
rom[57977] = 12'haaa;
rom[57978] = 12'haaa;
rom[57979] = 12'haaa;
rom[57980] = 12'h999;
rom[57981] = 12'h999;
rom[57982] = 12'h999;
rom[57983] = 12'h999;
rom[57984] = 12'h999;
rom[57985] = 12'h999;
rom[57986] = 12'h999;
rom[57987] = 12'h999;
rom[57988] = 12'h999;
rom[57989] = 12'h999;
rom[57990] = 12'h999;
rom[57991] = 12'h999;
rom[57992] = 12'h999;
rom[57993] = 12'h999;
rom[57994] = 12'h999;
rom[57995] = 12'h999;
rom[57996] = 12'h999;
rom[57997] = 12'h999;
rom[57998] = 12'h999;
rom[57999] = 12'h999;
rom[58000] = 12'hfff;
rom[58001] = 12'hfff;
rom[58002] = 12'hfff;
rom[58003] = 12'hfff;
rom[58004] = 12'hfff;
rom[58005] = 12'hfff;
rom[58006] = 12'hfff;
rom[58007] = 12'hfff;
rom[58008] = 12'hfff;
rom[58009] = 12'hfff;
rom[58010] = 12'hfff;
rom[58011] = 12'hfff;
rom[58012] = 12'hfff;
rom[58013] = 12'hfff;
rom[58014] = 12'hfff;
rom[58015] = 12'hfff;
rom[58016] = 12'hfff;
rom[58017] = 12'hfff;
rom[58018] = 12'hfff;
rom[58019] = 12'hfff;
rom[58020] = 12'hfff;
rom[58021] = 12'hfff;
rom[58022] = 12'hfff;
rom[58023] = 12'hfff;
rom[58024] = 12'hfff;
rom[58025] = 12'hfff;
rom[58026] = 12'hfff;
rom[58027] = 12'hfff;
rom[58028] = 12'hfff;
rom[58029] = 12'hfff;
rom[58030] = 12'hfff;
rom[58031] = 12'hfff;
rom[58032] = 12'hfff;
rom[58033] = 12'hfff;
rom[58034] = 12'hfff;
rom[58035] = 12'hfff;
rom[58036] = 12'hfff;
rom[58037] = 12'hfff;
rom[58038] = 12'hfff;
rom[58039] = 12'hfff;
rom[58040] = 12'hfff;
rom[58041] = 12'hfff;
rom[58042] = 12'hfff;
rom[58043] = 12'hfff;
rom[58044] = 12'hfff;
rom[58045] = 12'hfff;
rom[58046] = 12'hfff;
rom[58047] = 12'hfff;
rom[58048] = 12'hfff;
rom[58049] = 12'hfff;
rom[58050] = 12'hfff;
rom[58051] = 12'hfff;
rom[58052] = 12'hfff;
rom[58053] = 12'hfff;
rom[58054] = 12'hfff;
rom[58055] = 12'hfff;
rom[58056] = 12'hfff;
rom[58057] = 12'hfff;
rom[58058] = 12'hfff;
rom[58059] = 12'hfff;
rom[58060] = 12'hfff;
rom[58061] = 12'hfff;
rom[58062] = 12'hfff;
rom[58063] = 12'hfff;
rom[58064] = 12'hfff;
rom[58065] = 12'hfff;
rom[58066] = 12'hfff;
rom[58067] = 12'hfff;
rom[58068] = 12'hfff;
rom[58069] = 12'hfff;
rom[58070] = 12'hfff;
rom[58071] = 12'hfff;
rom[58072] = 12'hfff;
rom[58073] = 12'hfff;
rom[58074] = 12'hfff;
rom[58075] = 12'hfff;
rom[58076] = 12'hfff;
rom[58077] = 12'hfff;
rom[58078] = 12'hfff;
rom[58079] = 12'hfff;
rom[58080] = 12'hfff;
rom[58081] = 12'hfff;
rom[58082] = 12'hfff;
rom[58083] = 12'hfff;
rom[58084] = 12'hfff;
rom[58085] = 12'hfff;
rom[58086] = 12'heee;
rom[58087] = 12'heee;
rom[58088] = 12'heee;
rom[58089] = 12'hddd;
rom[58090] = 12'hddd;
rom[58091] = 12'hddd;
rom[58092] = 12'hccc;
rom[58093] = 12'hccc;
rom[58094] = 12'hccc;
rom[58095] = 12'hccc;
rom[58096] = 12'hccc;
rom[58097] = 12'hbbb;
rom[58098] = 12'hbbb;
rom[58099] = 12'hbbb;
rom[58100] = 12'hccc;
rom[58101] = 12'hccc;
rom[58102] = 12'hccc;
rom[58103] = 12'hccc;
rom[58104] = 12'hddd;
rom[58105] = 12'heee;
rom[58106] = 12'heee;
rom[58107] = 12'heee;
rom[58108] = 12'hddd;
rom[58109] = 12'hddd;
rom[58110] = 12'hccc;
rom[58111] = 12'hccc;
rom[58112] = 12'hbbb;
rom[58113] = 12'hbbb;
rom[58114] = 12'haaa;
rom[58115] = 12'haaa;
rom[58116] = 12'haaa;
rom[58117] = 12'h999;
rom[58118] = 12'h999;
rom[58119] = 12'h999;
rom[58120] = 12'h888;
rom[58121] = 12'h888;
rom[58122] = 12'h888;
rom[58123] = 12'h888;
rom[58124] = 12'h888;
rom[58125] = 12'h888;
rom[58126] = 12'h888;
rom[58127] = 12'h888;
rom[58128] = 12'h777;
rom[58129] = 12'h888;
rom[58130] = 12'h888;
rom[58131] = 12'h888;
rom[58132] = 12'h888;
rom[58133] = 12'h888;
rom[58134] = 12'h777;
rom[58135] = 12'h777;
rom[58136] = 12'h666;
rom[58137] = 12'h666;
rom[58138] = 12'h555;
rom[58139] = 12'h555;
rom[58140] = 12'h444;
rom[58141] = 12'h444;
rom[58142] = 12'h444;
rom[58143] = 12'h333;
rom[58144] = 12'h333;
rom[58145] = 12'h333;
rom[58146] = 12'h333;
rom[58147] = 12'h222;
rom[58148] = 12'h222;
rom[58149] = 12'h222;
rom[58150] = 12'h222;
rom[58151] = 12'h222;
rom[58152] = 12'h222;
rom[58153] = 12'h222;
rom[58154] = 12'h111;
rom[58155] = 12'h111;
rom[58156] = 12'h222;
rom[58157] = 12'h222;
rom[58158] = 12'h111;
rom[58159] = 12'h111;
rom[58160] = 12'h111;
rom[58161] = 12'h111;
rom[58162] = 12'h111;
rom[58163] = 12'h111;
rom[58164] = 12'h111;
rom[58165] = 12'h111;
rom[58166] = 12'h111;
rom[58167] = 12'h111;
rom[58168] = 12'h111;
rom[58169] = 12'h111;
rom[58170] = 12'h111;
rom[58171] = 12'h111;
rom[58172] = 12'h111;
rom[58173] = 12'h111;
rom[58174] = 12'h111;
rom[58175] = 12'h111;
rom[58176] = 12'h111;
rom[58177] = 12'h111;
rom[58178] = 12'h111;
rom[58179] = 12'h111;
rom[58180] = 12'h  0;
rom[58181] = 12'h  0;
rom[58182] = 12'h  0;
rom[58183] = 12'h  0;
rom[58184] = 12'h  0;
rom[58185] = 12'h  0;
rom[58186] = 12'h  0;
rom[58187] = 12'h  0;
rom[58188] = 12'h  0;
rom[58189] = 12'h  0;
rom[58190] = 12'h  0;
rom[58191] = 12'h  0;
rom[58192] = 12'h  0;
rom[58193] = 12'h  0;
rom[58194] = 12'h  0;
rom[58195] = 12'h  0;
rom[58196] = 12'h  0;
rom[58197] = 12'h  0;
rom[58198] = 12'h  0;
rom[58199] = 12'h  0;
rom[58200] = 12'h  0;
rom[58201] = 12'h  0;
rom[58202] = 12'h  0;
rom[58203] = 12'h  0;
rom[58204] = 12'h111;
rom[58205] = 12'h111;
rom[58206] = 12'h111;
rom[58207] = 12'h111;
rom[58208] = 12'h111;
rom[58209] = 12'h  0;
rom[58210] = 12'h  0;
rom[58211] = 12'h111;
rom[58212] = 12'h111;
rom[58213] = 12'h111;
rom[58214] = 12'h111;
rom[58215] = 12'h222;
rom[58216] = 12'h333;
rom[58217] = 12'h333;
rom[58218] = 12'h333;
rom[58219] = 12'h222;
rom[58220] = 12'h222;
rom[58221] = 12'h111;
rom[58222] = 12'h111;
rom[58223] = 12'h111;
rom[58224] = 12'h111;
rom[58225] = 12'h111;
rom[58226] = 12'h  0;
rom[58227] = 12'h  0;
rom[58228] = 12'h  0;
rom[58229] = 12'h  0;
rom[58230] = 12'h  0;
rom[58231] = 12'h  0;
rom[58232] = 12'h  0;
rom[58233] = 12'h  0;
rom[58234] = 12'h  0;
rom[58235] = 12'h  0;
rom[58236] = 12'h  0;
rom[58237] = 12'h  0;
rom[58238] = 12'h  0;
rom[58239] = 12'h  0;
rom[58240] = 12'h  0;
rom[58241] = 12'h  0;
rom[58242] = 12'h  0;
rom[58243] = 12'h  0;
rom[58244] = 12'h  0;
rom[58245] = 12'h  0;
rom[58246] = 12'h  0;
rom[58247] = 12'h  0;
rom[58248] = 12'h  0;
rom[58249] = 12'h  0;
rom[58250] = 12'h  0;
rom[58251] = 12'h  0;
rom[58252] = 12'h  0;
rom[58253] = 12'h  0;
rom[58254] = 12'h  0;
rom[58255] = 12'h  0;
rom[58256] = 12'h  0;
rom[58257] = 12'h  0;
rom[58258] = 12'h  0;
rom[58259] = 12'h  0;
rom[58260] = 12'h  0;
rom[58261] = 12'h  0;
rom[58262] = 12'h  0;
rom[58263] = 12'h  0;
rom[58264] = 12'h  0;
rom[58265] = 12'h  0;
rom[58266] = 12'h  0;
rom[58267] = 12'h  0;
rom[58268] = 12'h  0;
rom[58269] = 12'h  0;
rom[58270] = 12'h  0;
rom[58271] = 12'h  0;
rom[58272] = 12'h  0;
rom[58273] = 12'h111;
rom[58274] = 12'h111;
rom[58275] = 12'h222;
rom[58276] = 12'h222;
rom[58277] = 12'h222;
rom[58278] = 12'h333;
rom[58279] = 12'h333;
rom[58280] = 12'h333;
rom[58281] = 12'h444;
rom[58282] = 12'h555;
rom[58283] = 12'h555;
rom[58284] = 12'h444;
rom[58285] = 12'h333;
rom[58286] = 12'h222;
rom[58287] = 12'h222;
rom[58288] = 12'h222;
rom[58289] = 12'h222;
rom[58290] = 12'h333;
rom[58291] = 12'h333;
rom[58292] = 12'h333;
rom[58293] = 12'h333;
rom[58294] = 12'h333;
rom[58295] = 12'h444;
rom[58296] = 12'h555;
rom[58297] = 12'h666;
rom[58298] = 12'h666;
rom[58299] = 12'h666;
rom[58300] = 12'h555;
rom[58301] = 12'h555;
rom[58302] = 12'h555;
rom[58303] = 12'h555;
rom[58304] = 12'h666;
rom[58305] = 12'h666;
rom[58306] = 12'h666;
rom[58307] = 12'h666;
rom[58308] = 12'h555;
rom[58309] = 12'h555;
rom[58310] = 12'h555;
rom[58311] = 12'h555;
rom[58312] = 12'h555;
rom[58313] = 12'h555;
rom[58314] = 12'h555;
rom[58315] = 12'h555;
rom[58316] = 12'h555;
rom[58317] = 12'h666;
rom[58318] = 12'h666;
rom[58319] = 12'h666;
rom[58320] = 12'h666;
rom[58321] = 12'h666;
rom[58322] = 12'h666;
rom[58323] = 12'h666;
rom[58324] = 12'h666;
rom[58325] = 12'h666;
rom[58326] = 12'h666;
rom[58327] = 12'h666;
rom[58328] = 12'h666;
rom[58329] = 12'h666;
rom[58330] = 12'h666;
rom[58331] = 12'h666;
rom[58332] = 12'h666;
rom[58333] = 12'h666;
rom[58334] = 12'h666;
rom[58335] = 12'h777;
rom[58336] = 12'h777;
rom[58337] = 12'h777;
rom[58338] = 12'h777;
rom[58339] = 12'h777;
rom[58340] = 12'h888;
rom[58341] = 12'h888;
rom[58342] = 12'h888;
rom[58343] = 12'h888;
rom[58344] = 12'h999;
rom[58345] = 12'h999;
rom[58346] = 12'h999;
rom[58347] = 12'h999;
rom[58348] = 12'h999;
rom[58349] = 12'haaa;
rom[58350] = 12'haaa;
rom[58351] = 12'haaa;
rom[58352] = 12'hbbb;
rom[58353] = 12'hbbb;
rom[58354] = 12'hbbb;
rom[58355] = 12'hccc;
rom[58356] = 12'hccc;
rom[58357] = 12'hccc;
rom[58358] = 12'hddd;
rom[58359] = 12'hddd;
rom[58360] = 12'heee;
rom[58361] = 12'heee;
rom[58362] = 12'heee;
rom[58363] = 12'hddd;
rom[58364] = 12'hddd;
rom[58365] = 12'hccc;
rom[58366] = 12'hccc;
rom[58367] = 12'hccc;
rom[58368] = 12'hbbb;
rom[58369] = 12'hbbb;
rom[58370] = 12'hbbb;
rom[58371] = 12'hbbb;
rom[58372] = 12'hbbb;
rom[58373] = 12'haaa;
rom[58374] = 12'haaa;
rom[58375] = 12'haaa;
rom[58376] = 12'haaa;
rom[58377] = 12'haaa;
rom[58378] = 12'haaa;
rom[58379] = 12'h999;
rom[58380] = 12'h999;
rom[58381] = 12'h999;
rom[58382] = 12'h999;
rom[58383] = 12'h999;
rom[58384] = 12'h999;
rom[58385] = 12'h999;
rom[58386] = 12'h999;
rom[58387] = 12'h999;
rom[58388] = 12'h999;
rom[58389] = 12'h999;
rom[58390] = 12'h999;
rom[58391] = 12'h999;
rom[58392] = 12'h999;
rom[58393] = 12'h999;
rom[58394] = 12'h888;
rom[58395] = 12'h999;
rom[58396] = 12'h999;
rom[58397] = 12'h999;
rom[58398] = 12'h999;
rom[58399] = 12'h999;
rom[58400] = 12'hfff;
rom[58401] = 12'hfff;
rom[58402] = 12'hfff;
rom[58403] = 12'hfff;
rom[58404] = 12'hfff;
rom[58405] = 12'hfff;
rom[58406] = 12'hfff;
rom[58407] = 12'hfff;
rom[58408] = 12'hfff;
rom[58409] = 12'hfff;
rom[58410] = 12'hfff;
rom[58411] = 12'hfff;
rom[58412] = 12'hfff;
rom[58413] = 12'hfff;
rom[58414] = 12'hfff;
rom[58415] = 12'hfff;
rom[58416] = 12'hfff;
rom[58417] = 12'hfff;
rom[58418] = 12'hfff;
rom[58419] = 12'hfff;
rom[58420] = 12'hfff;
rom[58421] = 12'hfff;
rom[58422] = 12'hfff;
rom[58423] = 12'hfff;
rom[58424] = 12'hfff;
rom[58425] = 12'hfff;
rom[58426] = 12'hfff;
rom[58427] = 12'hfff;
rom[58428] = 12'hfff;
rom[58429] = 12'hfff;
rom[58430] = 12'hfff;
rom[58431] = 12'hfff;
rom[58432] = 12'hfff;
rom[58433] = 12'hfff;
rom[58434] = 12'hfff;
rom[58435] = 12'hfff;
rom[58436] = 12'hfff;
rom[58437] = 12'hfff;
rom[58438] = 12'hfff;
rom[58439] = 12'hfff;
rom[58440] = 12'hfff;
rom[58441] = 12'hfff;
rom[58442] = 12'hfff;
rom[58443] = 12'hfff;
rom[58444] = 12'hfff;
rom[58445] = 12'hfff;
rom[58446] = 12'hfff;
rom[58447] = 12'hfff;
rom[58448] = 12'hfff;
rom[58449] = 12'hfff;
rom[58450] = 12'hfff;
rom[58451] = 12'hfff;
rom[58452] = 12'hfff;
rom[58453] = 12'hfff;
rom[58454] = 12'hfff;
rom[58455] = 12'hfff;
rom[58456] = 12'hfff;
rom[58457] = 12'hfff;
rom[58458] = 12'hfff;
rom[58459] = 12'hfff;
rom[58460] = 12'hfff;
rom[58461] = 12'hfff;
rom[58462] = 12'hfff;
rom[58463] = 12'hfff;
rom[58464] = 12'hfff;
rom[58465] = 12'hfff;
rom[58466] = 12'hfff;
rom[58467] = 12'hfff;
rom[58468] = 12'hfff;
rom[58469] = 12'hfff;
rom[58470] = 12'hfff;
rom[58471] = 12'hfff;
rom[58472] = 12'hfff;
rom[58473] = 12'hfff;
rom[58474] = 12'hfff;
rom[58475] = 12'hfff;
rom[58476] = 12'hfff;
rom[58477] = 12'hfff;
rom[58478] = 12'hfff;
rom[58479] = 12'hfff;
rom[58480] = 12'hfff;
rom[58481] = 12'hfff;
rom[58482] = 12'hfff;
rom[58483] = 12'hfff;
rom[58484] = 12'hfff;
rom[58485] = 12'hfff;
rom[58486] = 12'hfff;
rom[58487] = 12'hfff;
rom[58488] = 12'heee;
rom[58489] = 12'heee;
rom[58490] = 12'heee;
rom[58491] = 12'hddd;
rom[58492] = 12'hddd;
rom[58493] = 12'hddd;
rom[58494] = 12'hccc;
rom[58495] = 12'hccc;
rom[58496] = 12'hccc;
rom[58497] = 12'hccc;
rom[58498] = 12'hccc;
rom[58499] = 12'hccc;
rom[58500] = 12'hbbb;
rom[58501] = 12'hbbb;
rom[58502] = 12'hbbb;
rom[58503] = 12'hbbb;
rom[58504] = 12'hccc;
rom[58505] = 12'hccc;
rom[58506] = 12'hddd;
rom[58507] = 12'hddd;
rom[58508] = 12'heee;
rom[58509] = 12'heee;
rom[58510] = 12'heee;
rom[58511] = 12'heee;
rom[58512] = 12'hddd;
rom[58513] = 12'hccc;
rom[58514] = 12'hbbb;
rom[58515] = 12'hbbb;
rom[58516] = 12'hbbb;
rom[58517] = 12'hbbb;
rom[58518] = 12'haaa;
rom[58519] = 12'haaa;
rom[58520] = 12'h999;
rom[58521] = 12'h888;
rom[58522] = 12'h888;
rom[58523] = 12'h888;
rom[58524] = 12'h888;
rom[58525] = 12'h888;
rom[58526] = 12'h888;
rom[58527] = 12'h888;
rom[58528] = 12'h777;
rom[58529] = 12'h777;
rom[58530] = 12'h888;
rom[58531] = 12'h888;
rom[58532] = 12'h888;
rom[58533] = 12'h888;
rom[58534] = 12'h777;
rom[58535] = 12'h777;
rom[58536] = 12'h666;
rom[58537] = 12'h666;
rom[58538] = 12'h555;
rom[58539] = 12'h555;
rom[58540] = 12'h444;
rom[58541] = 12'h444;
rom[58542] = 12'h444;
rom[58543] = 12'h333;
rom[58544] = 12'h333;
rom[58545] = 12'h333;
rom[58546] = 12'h333;
rom[58547] = 12'h222;
rom[58548] = 12'h222;
rom[58549] = 12'h222;
rom[58550] = 12'h222;
rom[58551] = 12'h222;
rom[58552] = 12'h222;
rom[58553] = 12'h111;
rom[58554] = 12'h111;
rom[58555] = 12'h111;
rom[58556] = 12'h222;
rom[58557] = 12'h222;
rom[58558] = 12'h111;
rom[58559] = 12'h111;
rom[58560] = 12'h111;
rom[58561] = 12'h111;
rom[58562] = 12'h111;
rom[58563] = 12'h111;
rom[58564] = 12'h111;
rom[58565] = 12'h111;
rom[58566] = 12'h111;
rom[58567] = 12'h111;
rom[58568] = 12'h111;
rom[58569] = 12'h111;
rom[58570] = 12'h111;
rom[58571] = 12'h111;
rom[58572] = 12'h111;
rom[58573] = 12'h111;
rom[58574] = 12'h111;
rom[58575] = 12'h111;
rom[58576] = 12'h111;
rom[58577] = 12'h111;
rom[58578] = 12'h  0;
rom[58579] = 12'h  0;
rom[58580] = 12'h  0;
rom[58581] = 12'h  0;
rom[58582] = 12'h  0;
rom[58583] = 12'h  0;
rom[58584] = 12'h  0;
rom[58585] = 12'h  0;
rom[58586] = 12'h  0;
rom[58587] = 12'h  0;
rom[58588] = 12'h  0;
rom[58589] = 12'h  0;
rom[58590] = 12'h  0;
rom[58591] = 12'h  0;
rom[58592] = 12'h  0;
rom[58593] = 12'h  0;
rom[58594] = 12'h  0;
rom[58595] = 12'h  0;
rom[58596] = 12'h  0;
rom[58597] = 12'h  0;
rom[58598] = 12'h  0;
rom[58599] = 12'h  0;
rom[58600] = 12'h  0;
rom[58601] = 12'h  0;
rom[58602] = 12'h  0;
rom[58603] = 12'h  0;
rom[58604] = 12'h111;
rom[58605] = 12'h111;
rom[58606] = 12'h111;
rom[58607] = 12'h111;
rom[58608] = 12'h111;
rom[58609] = 12'h  0;
rom[58610] = 12'h111;
rom[58611] = 12'h111;
rom[58612] = 12'h111;
rom[58613] = 12'h111;
rom[58614] = 12'h111;
rom[58615] = 12'h222;
rom[58616] = 12'h333;
rom[58617] = 12'h333;
rom[58618] = 12'h222;
rom[58619] = 12'h222;
rom[58620] = 12'h111;
rom[58621] = 12'h111;
rom[58622] = 12'h111;
rom[58623] = 12'h111;
rom[58624] = 12'h111;
rom[58625] = 12'h111;
rom[58626] = 12'h  0;
rom[58627] = 12'h  0;
rom[58628] = 12'h  0;
rom[58629] = 12'h  0;
rom[58630] = 12'h  0;
rom[58631] = 12'h  0;
rom[58632] = 12'h  0;
rom[58633] = 12'h  0;
rom[58634] = 12'h  0;
rom[58635] = 12'h  0;
rom[58636] = 12'h  0;
rom[58637] = 12'h  0;
rom[58638] = 12'h  0;
rom[58639] = 12'h  0;
rom[58640] = 12'h  0;
rom[58641] = 12'h  0;
rom[58642] = 12'h  0;
rom[58643] = 12'h  0;
rom[58644] = 12'h  0;
rom[58645] = 12'h  0;
rom[58646] = 12'h  0;
rom[58647] = 12'h  0;
rom[58648] = 12'h  0;
rom[58649] = 12'h  0;
rom[58650] = 12'h  0;
rom[58651] = 12'h  0;
rom[58652] = 12'h  0;
rom[58653] = 12'h  0;
rom[58654] = 12'h  0;
rom[58655] = 12'h  0;
rom[58656] = 12'h  0;
rom[58657] = 12'h  0;
rom[58658] = 12'h  0;
rom[58659] = 12'h  0;
rom[58660] = 12'h  0;
rom[58661] = 12'h  0;
rom[58662] = 12'h  0;
rom[58663] = 12'h  0;
rom[58664] = 12'h  0;
rom[58665] = 12'h  0;
rom[58666] = 12'h  0;
rom[58667] = 12'h  0;
rom[58668] = 12'h  0;
rom[58669] = 12'h  0;
rom[58670] = 12'h  0;
rom[58671] = 12'h  0;
rom[58672] = 12'h111;
rom[58673] = 12'h111;
rom[58674] = 12'h111;
rom[58675] = 12'h222;
rom[58676] = 12'h222;
rom[58677] = 12'h222;
rom[58678] = 12'h333;
rom[58679] = 12'h333;
rom[58680] = 12'h333;
rom[58681] = 12'h444;
rom[58682] = 12'h555;
rom[58683] = 12'h555;
rom[58684] = 12'h444;
rom[58685] = 12'h333;
rom[58686] = 12'h222;
rom[58687] = 12'h222;
rom[58688] = 12'h222;
rom[58689] = 12'h222;
rom[58690] = 12'h333;
rom[58691] = 12'h333;
rom[58692] = 12'h333;
rom[58693] = 12'h333;
rom[58694] = 12'h333;
rom[58695] = 12'h444;
rom[58696] = 12'h555;
rom[58697] = 12'h555;
rom[58698] = 12'h666;
rom[58699] = 12'h666;
rom[58700] = 12'h555;
rom[58701] = 12'h555;
rom[58702] = 12'h555;
rom[58703] = 12'h555;
rom[58704] = 12'h555;
rom[58705] = 12'h666;
rom[58706] = 12'h666;
rom[58707] = 12'h666;
rom[58708] = 12'h666;
rom[58709] = 12'h555;
rom[58710] = 12'h555;
rom[58711] = 12'h555;
rom[58712] = 12'h444;
rom[58713] = 12'h555;
rom[58714] = 12'h555;
rom[58715] = 12'h555;
rom[58716] = 12'h555;
rom[58717] = 12'h666;
rom[58718] = 12'h666;
rom[58719] = 12'h666;
rom[58720] = 12'h666;
rom[58721] = 12'h666;
rom[58722] = 12'h666;
rom[58723] = 12'h666;
rom[58724] = 12'h666;
rom[58725] = 12'h666;
rom[58726] = 12'h666;
rom[58727] = 12'h666;
rom[58728] = 12'h666;
rom[58729] = 12'h666;
rom[58730] = 12'h666;
rom[58731] = 12'h666;
rom[58732] = 12'h666;
rom[58733] = 12'h666;
rom[58734] = 12'h777;
rom[58735] = 12'h777;
rom[58736] = 12'h777;
rom[58737] = 12'h777;
rom[58738] = 12'h777;
rom[58739] = 12'h888;
rom[58740] = 12'h888;
rom[58741] = 12'h888;
rom[58742] = 12'h888;
rom[58743] = 12'h888;
rom[58744] = 12'h999;
rom[58745] = 12'h999;
rom[58746] = 12'h999;
rom[58747] = 12'haaa;
rom[58748] = 12'haaa;
rom[58749] = 12'haaa;
rom[58750] = 12'haaa;
rom[58751] = 12'hbbb;
rom[58752] = 12'hbbb;
rom[58753] = 12'hbbb;
rom[58754] = 12'hccc;
rom[58755] = 12'hccc;
rom[58756] = 12'hccc;
rom[58757] = 12'hddd;
rom[58758] = 12'heee;
rom[58759] = 12'heee;
rom[58760] = 12'heee;
rom[58761] = 12'heee;
rom[58762] = 12'heee;
rom[58763] = 12'hddd;
rom[58764] = 12'hddd;
rom[58765] = 12'hccc;
rom[58766] = 12'hccc;
rom[58767] = 12'hbbb;
rom[58768] = 12'hbbb;
rom[58769] = 12'hbbb;
rom[58770] = 12'hbbb;
rom[58771] = 12'hbbb;
rom[58772] = 12'haaa;
rom[58773] = 12'haaa;
rom[58774] = 12'haaa;
rom[58775] = 12'haaa;
rom[58776] = 12'haaa;
rom[58777] = 12'haaa;
rom[58778] = 12'h999;
rom[58779] = 12'h999;
rom[58780] = 12'h999;
rom[58781] = 12'h999;
rom[58782] = 12'h999;
rom[58783] = 12'h999;
rom[58784] = 12'h999;
rom[58785] = 12'h999;
rom[58786] = 12'h999;
rom[58787] = 12'h999;
rom[58788] = 12'h999;
rom[58789] = 12'h999;
rom[58790] = 12'h999;
rom[58791] = 12'h999;
rom[58792] = 12'h888;
rom[58793] = 12'h888;
rom[58794] = 12'h888;
rom[58795] = 12'h888;
rom[58796] = 12'h888;
rom[58797] = 12'h888;
rom[58798] = 12'h888;
rom[58799] = 12'h888;
rom[58800] = 12'hfff;
rom[58801] = 12'hfff;
rom[58802] = 12'hfff;
rom[58803] = 12'hfff;
rom[58804] = 12'hfff;
rom[58805] = 12'hfff;
rom[58806] = 12'hfff;
rom[58807] = 12'hfff;
rom[58808] = 12'hfff;
rom[58809] = 12'hfff;
rom[58810] = 12'hfff;
rom[58811] = 12'hfff;
rom[58812] = 12'hfff;
rom[58813] = 12'hfff;
rom[58814] = 12'hfff;
rom[58815] = 12'hfff;
rom[58816] = 12'hfff;
rom[58817] = 12'hfff;
rom[58818] = 12'hfff;
rom[58819] = 12'hfff;
rom[58820] = 12'hfff;
rom[58821] = 12'hfff;
rom[58822] = 12'hfff;
rom[58823] = 12'hfff;
rom[58824] = 12'hfff;
rom[58825] = 12'hfff;
rom[58826] = 12'hfff;
rom[58827] = 12'hfff;
rom[58828] = 12'hfff;
rom[58829] = 12'hfff;
rom[58830] = 12'hfff;
rom[58831] = 12'hfff;
rom[58832] = 12'hfff;
rom[58833] = 12'hfff;
rom[58834] = 12'hfff;
rom[58835] = 12'hfff;
rom[58836] = 12'hfff;
rom[58837] = 12'hfff;
rom[58838] = 12'hfff;
rom[58839] = 12'hfff;
rom[58840] = 12'hfff;
rom[58841] = 12'hfff;
rom[58842] = 12'hfff;
rom[58843] = 12'hfff;
rom[58844] = 12'hfff;
rom[58845] = 12'hfff;
rom[58846] = 12'hfff;
rom[58847] = 12'hfff;
rom[58848] = 12'hfff;
rom[58849] = 12'hfff;
rom[58850] = 12'hfff;
rom[58851] = 12'hfff;
rom[58852] = 12'hfff;
rom[58853] = 12'hfff;
rom[58854] = 12'hfff;
rom[58855] = 12'hfff;
rom[58856] = 12'hfff;
rom[58857] = 12'hfff;
rom[58858] = 12'hfff;
rom[58859] = 12'hfff;
rom[58860] = 12'hfff;
rom[58861] = 12'hfff;
rom[58862] = 12'hfff;
rom[58863] = 12'hfff;
rom[58864] = 12'hfff;
rom[58865] = 12'hfff;
rom[58866] = 12'hfff;
rom[58867] = 12'hfff;
rom[58868] = 12'hfff;
rom[58869] = 12'hfff;
rom[58870] = 12'hfff;
rom[58871] = 12'hfff;
rom[58872] = 12'hfff;
rom[58873] = 12'hfff;
rom[58874] = 12'hfff;
rom[58875] = 12'hfff;
rom[58876] = 12'hfff;
rom[58877] = 12'hfff;
rom[58878] = 12'hfff;
rom[58879] = 12'hfff;
rom[58880] = 12'hfff;
rom[58881] = 12'hfff;
rom[58882] = 12'hfff;
rom[58883] = 12'hfff;
rom[58884] = 12'hfff;
rom[58885] = 12'hfff;
rom[58886] = 12'hfff;
rom[58887] = 12'hfff;
rom[58888] = 12'hfff;
rom[58889] = 12'hfff;
rom[58890] = 12'heee;
rom[58891] = 12'heee;
rom[58892] = 12'heee;
rom[58893] = 12'hddd;
rom[58894] = 12'hddd;
rom[58895] = 12'hddd;
rom[58896] = 12'hddd;
rom[58897] = 12'hddd;
rom[58898] = 12'hccc;
rom[58899] = 12'hccc;
rom[58900] = 12'hccc;
rom[58901] = 12'hccc;
rom[58902] = 12'hccc;
rom[58903] = 12'hccc;
rom[58904] = 12'hbbb;
rom[58905] = 12'hbbb;
rom[58906] = 12'hbbb;
rom[58907] = 12'hccc;
rom[58908] = 12'hccc;
rom[58909] = 12'hddd;
rom[58910] = 12'heee;
rom[58911] = 12'heee;
rom[58912] = 12'heee;
rom[58913] = 12'hddd;
rom[58914] = 12'hddd;
rom[58915] = 12'hccc;
rom[58916] = 12'hccc;
rom[58917] = 12'hccc;
rom[58918] = 12'hbbb;
rom[58919] = 12'hbbb;
rom[58920] = 12'haaa;
rom[58921] = 12'haaa;
rom[58922] = 12'h999;
rom[58923] = 12'h999;
rom[58924] = 12'h999;
rom[58925] = 12'h888;
rom[58926] = 12'h888;
rom[58927] = 12'h888;
rom[58928] = 12'h888;
rom[58929] = 12'h777;
rom[58930] = 12'h777;
rom[58931] = 12'h777;
rom[58932] = 12'h777;
rom[58933] = 12'h777;
rom[58934] = 12'h777;
rom[58935] = 12'h777;
rom[58936] = 12'h777;
rom[58937] = 12'h666;
rom[58938] = 12'h666;
rom[58939] = 12'h555;
rom[58940] = 12'h555;
rom[58941] = 12'h444;
rom[58942] = 12'h444;
rom[58943] = 12'h444;
rom[58944] = 12'h333;
rom[58945] = 12'h333;
rom[58946] = 12'h333;
rom[58947] = 12'h222;
rom[58948] = 12'h222;
rom[58949] = 12'h222;
rom[58950] = 12'h222;
rom[58951] = 12'h222;
rom[58952] = 12'h222;
rom[58953] = 12'h222;
rom[58954] = 12'h222;
rom[58955] = 12'h222;
rom[58956] = 12'h222;
rom[58957] = 12'h222;
rom[58958] = 12'h222;
rom[58959] = 12'h222;
rom[58960] = 12'h111;
rom[58961] = 12'h111;
rom[58962] = 12'h111;
rom[58963] = 12'h111;
rom[58964] = 12'h111;
rom[58965] = 12'h111;
rom[58966] = 12'h111;
rom[58967] = 12'h111;
rom[58968] = 12'h111;
rom[58969] = 12'h111;
rom[58970] = 12'h111;
rom[58971] = 12'h111;
rom[58972] = 12'h111;
rom[58973] = 12'h111;
rom[58974] = 12'h111;
rom[58975] = 12'h111;
rom[58976] = 12'h111;
rom[58977] = 12'h  0;
rom[58978] = 12'h  0;
rom[58979] = 12'h  0;
rom[58980] = 12'h  0;
rom[58981] = 12'h  0;
rom[58982] = 12'h  0;
rom[58983] = 12'h  0;
rom[58984] = 12'h  0;
rom[58985] = 12'h  0;
rom[58986] = 12'h  0;
rom[58987] = 12'h  0;
rom[58988] = 12'h  0;
rom[58989] = 12'h  0;
rom[58990] = 12'h  0;
rom[58991] = 12'h  0;
rom[58992] = 12'h  0;
rom[58993] = 12'h  0;
rom[58994] = 12'h  0;
rom[58995] = 12'h  0;
rom[58996] = 12'h  0;
rom[58997] = 12'h  0;
rom[58998] = 12'h  0;
rom[58999] = 12'h  0;
rom[59000] = 12'h  0;
rom[59001] = 12'h  0;
rom[59002] = 12'h  0;
rom[59003] = 12'h  0;
rom[59004] = 12'h111;
rom[59005] = 12'h111;
rom[59006] = 12'h111;
rom[59007] = 12'h111;
rom[59008] = 12'h  0;
rom[59009] = 12'h111;
rom[59010] = 12'h111;
rom[59011] = 12'h111;
rom[59012] = 12'h111;
rom[59013] = 12'h111;
rom[59014] = 12'h222;
rom[59015] = 12'h222;
rom[59016] = 12'h333;
rom[59017] = 12'h333;
rom[59018] = 12'h222;
rom[59019] = 12'h111;
rom[59020] = 12'h111;
rom[59021] = 12'h111;
rom[59022] = 12'h111;
rom[59023] = 12'h  0;
rom[59024] = 12'h111;
rom[59025] = 12'h111;
rom[59026] = 12'h  0;
rom[59027] = 12'h  0;
rom[59028] = 12'h  0;
rom[59029] = 12'h  0;
rom[59030] = 12'h  0;
rom[59031] = 12'h  0;
rom[59032] = 12'h  0;
rom[59033] = 12'h  0;
rom[59034] = 12'h  0;
rom[59035] = 12'h  0;
rom[59036] = 12'h  0;
rom[59037] = 12'h  0;
rom[59038] = 12'h  0;
rom[59039] = 12'h  0;
rom[59040] = 12'h  0;
rom[59041] = 12'h  0;
rom[59042] = 12'h  0;
rom[59043] = 12'h  0;
rom[59044] = 12'h  0;
rom[59045] = 12'h  0;
rom[59046] = 12'h  0;
rom[59047] = 12'h  0;
rom[59048] = 12'h  0;
rom[59049] = 12'h  0;
rom[59050] = 12'h  0;
rom[59051] = 12'h  0;
rom[59052] = 12'h  0;
rom[59053] = 12'h  0;
rom[59054] = 12'h  0;
rom[59055] = 12'h  0;
rom[59056] = 12'h  0;
rom[59057] = 12'h  0;
rom[59058] = 12'h  0;
rom[59059] = 12'h  0;
rom[59060] = 12'h  0;
rom[59061] = 12'h  0;
rom[59062] = 12'h  0;
rom[59063] = 12'h  0;
rom[59064] = 12'h  0;
rom[59065] = 12'h  0;
rom[59066] = 12'h  0;
rom[59067] = 12'h  0;
rom[59068] = 12'h  0;
rom[59069] = 12'h  0;
rom[59070] = 12'h  0;
rom[59071] = 12'h  0;
rom[59072] = 12'h111;
rom[59073] = 12'h111;
rom[59074] = 12'h111;
rom[59075] = 12'h222;
rom[59076] = 12'h222;
rom[59077] = 12'h222;
rom[59078] = 12'h333;
rom[59079] = 12'h333;
rom[59080] = 12'h333;
rom[59081] = 12'h444;
rom[59082] = 12'h555;
rom[59083] = 12'h555;
rom[59084] = 12'h444;
rom[59085] = 12'h333;
rom[59086] = 12'h222;
rom[59087] = 12'h222;
rom[59088] = 12'h222;
rom[59089] = 12'h222;
rom[59090] = 12'h333;
rom[59091] = 12'h333;
rom[59092] = 12'h333;
rom[59093] = 12'h333;
rom[59094] = 12'h333;
rom[59095] = 12'h333;
rom[59096] = 12'h444;
rom[59097] = 12'h555;
rom[59098] = 12'h666;
rom[59099] = 12'h666;
rom[59100] = 12'h555;
rom[59101] = 12'h555;
rom[59102] = 12'h555;
rom[59103] = 12'h555;
rom[59104] = 12'h555;
rom[59105] = 12'h666;
rom[59106] = 12'h666;
rom[59107] = 12'h666;
rom[59108] = 12'h666;
rom[59109] = 12'h666;
rom[59110] = 12'h555;
rom[59111] = 12'h555;
rom[59112] = 12'h555;
rom[59113] = 12'h555;
rom[59114] = 12'h555;
rom[59115] = 12'h555;
rom[59116] = 12'h555;
rom[59117] = 12'h555;
rom[59118] = 12'h666;
rom[59119] = 12'h666;
rom[59120] = 12'h666;
rom[59121] = 12'h666;
rom[59122] = 12'h666;
rom[59123] = 12'h666;
rom[59124] = 12'h666;
rom[59125] = 12'h666;
rom[59126] = 12'h666;
rom[59127] = 12'h666;
rom[59128] = 12'h666;
rom[59129] = 12'h666;
rom[59130] = 12'h666;
rom[59131] = 12'h666;
rom[59132] = 12'h777;
rom[59133] = 12'h777;
rom[59134] = 12'h777;
rom[59135] = 12'h777;
rom[59136] = 12'h777;
rom[59137] = 12'h777;
rom[59138] = 12'h777;
rom[59139] = 12'h888;
rom[59140] = 12'h888;
rom[59141] = 12'h888;
rom[59142] = 12'h999;
rom[59143] = 12'h999;
rom[59144] = 12'h999;
rom[59145] = 12'h999;
rom[59146] = 12'haaa;
rom[59147] = 12'haaa;
rom[59148] = 12'haaa;
rom[59149] = 12'haaa;
rom[59150] = 12'hbbb;
rom[59151] = 12'hbbb;
rom[59152] = 12'hbbb;
rom[59153] = 12'hccc;
rom[59154] = 12'hccc;
rom[59155] = 12'hccc;
rom[59156] = 12'hddd;
rom[59157] = 12'heee;
rom[59158] = 12'heee;
rom[59159] = 12'hfff;
rom[59160] = 12'heee;
rom[59161] = 12'heee;
rom[59162] = 12'hddd;
rom[59163] = 12'hddd;
rom[59164] = 12'hccc;
rom[59165] = 12'hccc;
rom[59166] = 12'hccc;
rom[59167] = 12'hbbb;
rom[59168] = 12'hbbb;
rom[59169] = 12'hbbb;
rom[59170] = 12'hbbb;
rom[59171] = 12'hbbb;
rom[59172] = 12'haaa;
rom[59173] = 12'haaa;
rom[59174] = 12'haaa;
rom[59175] = 12'haaa;
rom[59176] = 12'haaa;
rom[59177] = 12'haaa;
rom[59178] = 12'h999;
rom[59179] = 12'h999;
rom[59180] = 12'h999;
rom[59181] = 12'h999;
rom[59182] = 12'h999;
rom[59183] = 12'h888;
rom[59184] = 12'h888;
rom[59185] = 12'h888;
rom[59186] = 12'h888;
rom[59187] = 12'h888;
rom[59188] = 12'h888;
rom[59189] = 12'h888;
rom[59190] = 12'h888;
rom[59191] = 12'h888;
rom[59192] = 12'h888;
rom[59193] = 12'h888;
rom[59194] = 12'h888;
rom[59195] = 12'h888;
rom[59196] = 12'h888;
rom[59197] = 12'h888;
rom[59198] = 12'h888;
rom[59199] = 12'h888;
rom[59200] = 12'hfff;
rom[59201] = 12'hfff;
rom[59202] = 12'hfff;
rom[59203] = 12'hfff;
rom[59204] = 12'hfff;
rom[59205] = 12'hfff;
rom[59206] = 12'hfff;
rom[59207] = 12'hfff;
rom[59208] = 12'hfff;
rom[59209] = 12'hfff;
rom[59210] = 12'hfff;
rom[59211] = 12'hfff;
rom[59212] = 12'hfff;
rom[59213] = 12'hfff;
rom[59214] = 12'hfff;
rom[59215] = 12'hfff;
rom[59216] = 12'hfff;
rom[59217] = 12'hfff;
rom[59218] = 12'hfff;
rom[59219] = 12'hfff;
rom[59220] = 12'hfff;
rom[59221] = 12'hfff;
rom[59222] = 12'hfff;
rom[59223] = 12'hfff;
rom[59224] = 12'hfff;
rom[59225] = 12'hfff;
rom[59226] = 12'hfff;
rom[59227] = 12'hfff;
rom[59228] = 12'hfff;
rom[59229] = 12'hfff;
rom[59230] = 12'hfff;
rom[59231] = 12'hfff;
rom[59232] = 12'hfff;
rom[59233] = 12'hfff;
rom[59234] = 12'hfff;
rom[59235] = 12'hfff;
rom[59236] = 12'hfff;
rom[59237] = 12'hfff;
rom[59238] = 12'hfff;
rom[59239] = 12'hfff;
rom[59240] = 12'hfff;
rom[59241] = 12'hfff;
rom[59242] = 12'hfff;
rom[59243] = 12'hfff;
rom[59244] = 12'hfff;
rom[59245] = 12'hfff;
rom[59246] = 12'hfff;
rom[59247] = 12'hfff;
rom[59248] = 12'hfff;
rom[59249] = 12'hfff;
rom[59250] = 12'hfff;
rom[59251] = 12'hfff;
rom[59252] = 12'hfff;
rom[59253] = 12'hfff;
rom[59254] = 12'hfff;
rom[59255] = 12'hfff;
rom[59256] = 12'hfff;
rom[59257] = 12'hfff;
rom[59258] = 12'hfff;
rom[59259] = 12'hfff;
rom[59260] = 12'hfff;
rom[59261] = 12'hfff;
rom[59262] = 12'hfff;
rom[59263] = 12'hfff;
rom[59264] = 12'hfff;
rom[59265] = 12'hfff;
rom[59266] = 12'hfff;
rom[59267] = 12'hfff;
rom[59268] = 12'hfff;
rom[59269] = 12'hfff;
rom[59270] = 12'hfff;
rom[59271] = 12'hfff;
rom[59272] = 12'hfff;
rom[59273] = 12'hfff;
rom[59274] = 12'hfff;
rom[59275] = 12'hfff;
rom[59276] = 12'hfff;
rom[59277] = 12'hfff;
rom[59278] = 12'hfff;
rom[59279] = 12'hfff;
rom[59280] = 12'hfff;
rom[59281] = 12'hfff;
rom[59282] = 12'hfff;
rom[59283] = 12'hfff;
rom[59284] = 12'hfff;
rom[59285] = 12'hfff;
rom[59286] = 12'hfff;
rom[59287] = 12'hfff;
rom[59288] = 12'hfff;
rom[59289] = 12'hfff;
rom[59290] = 12'hfff;
rom[59291] = 12'hfff;
rom[59292] = 12'heee;
rom[59293] = 12'heee;
rom[59294] = 12'hddd;
rom[59295] = 12'hddd;
rom[59296] = 12'hddd;
rom[59297] = 12'hddd;
rom[59298] = 12'hddd;
rom[59299] = 12'hddd;
rom[59300] = 12'hccc;
rom[59301] = 12'hccc;
rom[59302] = 12'hccc;
rom[59303] = 12'hccc;
rom[59304] = 12'hccc;
rom[59305] = 12'hccc;
rom[59306] = 12'hccc;
rom[59307] = 12'hccc;
rom[59308] = 12'hccc;
rom[59309] = 12'hccc;
rom[59310] = 12'hccc;
rom[59311] = 12'hccc;
rom[59312] = 12'hddd;
rom[59313] = 12'hddd;
rom[59314] = 12'hddd;
rom[59315] = 12'hddd;
rom[59316] = 12'hddd;
rom[59317] = 12'hccc;
rom[59318] = 12'hccc;
rom[59319] = 12'hccc;
rom[59320] = 12'hccc;
rom[59321] = 12'hbbb;
rom[59322] = 12'hbbb;
rom[59323] = 12'haaa;
rom[59324] = 12'haaa;
rom[59325] = 12'h999;
rom[59326] = 12'h999;
rom[59327] = 12'h888;
rom[59328] = 12'h777;
rom[59329] = 12'h777;
rom[59330] = 12'h777;
rom[59331] = 12'h777;
rom[59332] = 12'h777;
rom[59333] = 12'h777;
rom[59334] = 12'h777;
rom[59335] = 12'h777;
rom[59336] = 12'h777;
rom[59337] = 12'h777;
rom[59338] = 12'h666;
rom[59339] = 12'h666;
rom[59340] = 12'h555;
rom[59341] = 12'h555;
rom[59342] = 12'h444;
rom[59343] = 12'h444;
rom[59344] = 12'h333;
rom[59345] = 12'h333;
rom[59346] = 12'h333;
rom[59347] = 12'h333;
rom[59348] = 12'h333;
rom[59349] = 12'h333;
rom[59350] = 12'h222;
rom[59351] = 12'h222;
rom[59352] = 12'h222;
rom[59353] = 12'h222;
rom[59354] = 12'h222;
rom[59355] = 12'h222;
rom[59356] = 12'h222;
rom[59357] = 12'h222;
rom[59358] = 12'h222;
rom[59359] = 12'h222;
rom[59360] = 12'h111;
rom[59361] = 12'h111;
rom[59362] = 12'h222;
rom[59363] = 12'h222;
rom[59364] = 12'h222;
rom[59365] = 12'h222;
rom[59366] = 12'h222;
rom[59367] = 12'h222;
rom[59368] = 12'h222;
rom[59369] = 12'h222;
rom[59370] = 12'h222;
rom[59371] = 12'h222;
rom[59372] = 12'h111;
rom[59373] = 12'h111;
rom[59374] = 12'h111;
rom[59375] = 12'h  0;
rom[59376] = 12'h  0;
rom[59377] = 12'h  0;
rom[59378] = 12'h  0;
rom[59379] = 12'h  0;
rom[59380] = 12'h  0;
rom[59381] = 12'h  0;
rom[59382] = 12'h  0;
rom[59383] = 12'h  0;
rom[59384] = 12'h  0;
rom[59385] = 12'h  0;
rom[59386] = 12'h  0;
rom[59387] = 12'h  0;
rom[59388] = 12'h  0;
rom[59389] = 12'h  0;
rom[59390] = 12'h  0;
rom[59391] = 12'h  0;
rom[59392] = 12'h  0;
rom[59393] = 12'h  0;
rom[59394] = 12'h  0;
rom[59395] = 12'h  0;
rom[59396] = 12'h  0;
rom[59397] = 12'h  0;
rom[59398] = 12'h  0;
rom[59399] = 12'h  0;
rom[59400] = 12'h  0;
rom[59401] = 12'h  0;
rom[59402] = 12'h  0;
rom[59403] = 12'h  0;
rom[59404] = 12'h111;
rom[59405] = 12'h111;
rom[59406] = 12'h111;
rom[59407] = 12'h111;
rom[59408] = 12'h  0;
rom[59409] = 12'h111;
rom[59410] = 12'h111;
rom[59411] = 12'h111;
rom[59412] = 12'h111;
rom[59413] = 12'h111;
rom[59414] = 12'h222;
rom[59415] = 12'h222;
rom[59416] = 12'h333;
rom[59417] = 12'h222;
rom[59418] = 12'h111;
rom[59419] = 12'h111;
rom[59420] = 12'h111;
rom[59421] = 12'h111;
rom[59422] = 12'h111;
rom[59423] = 12'h111;
rom[59424] = 12'h111;
rom[59425] = 12'h  0;
rom[59426] = 12'h  0;
rom[59427] = 12'h  0;
rom[59428] = 12'h  0;
rom[59429] = 12'h  0;
rom[59430] = 12'h  0;
rom[59431] = 12'h  0;
rom[59432] = 12'h  0;
rom[59433] = 12'h  0;
rom[59434] = 12'h  0;
rom[59435] = 12'h  0;
rom[59436] = 12'h  0;
rom[59437] = 12'h  0;
rom[59438] = 12'h  0;
rom[59439] = 12'h  0;
rom[59440] = 12'h  0;
rom[59441] = 12'h  0;
rom[59442] = 12'h  0;
rom[59443] = 12'h  0;
rom[59444] = 12'h  0;
rom[59445] = 12'h  0;
rom[59446] = 12'h  0;
rom[59447] = 12'h  0;
rom[59448] = 12'h  0;
rom[59449] = 12'h  0;
rom[59450] = 12'h  0;
rom[59451] = 12'h  0;
rom[59452] = 12'h  0;
rom[59453] = 12'h  0;
rom[59454] = 12'h  0;
rom[59455] = 12'h  0;
rom[59456] = 12'h  0;
rom[59457] = 12'h  0;
rom[59458] = 12'h  0;
rom[59459] = 12'h  0;
rom[59460] = 12'h  0;
rom[59461] = 12'h  0;
rom[59462] = 12'h  0;
rom[59463] = 12'h  0;
rom[59464] = 12'h  0;
rom[59465] = 12'h  0;
rom[59466] = 12'h  0;
rom[59467] = 12'h  0;
rom[59468] = 12'h  0;
rom[59469] = 12'h  0;
rom[59470] = 12'h  0;
rom[59471] = 12'h  0;
rom[59472] = 12'h111;
rom[59473] = 12'h111;
rom[59474] = 12'h111;
rom[59475] = 12'h222;
rom[59476] = 12'h222;
rom[59477] = 12'h333;
rom[59478] = 12'h333;
rom[59479] = 12'h333;
rom[59480] = 12'h444;
rom[59481] = 12'h444;
rom[59482] = 12'h555;
rom[59483] = 12'h555;
rom[59484] = 12'h444;
rom[59485] = 12'h333;
rom[59486] = 12'h222;
rom[59487] = 12'h222;
rom[59488] = 12'h222;
rom[59489] = 12'h222;
rom[59490] = 12'h222;
rom[59491] = 12'h222;
rom[59492] = 12'h222;
rom[59493] = 12'h333;
rom[59494] = 12'h333;
rom[59495] = 12'h333;
rom[59496] = 12'h444;
rom[59497] = 12'h555;
rom[59498] = 12'h666;
rom[59499] = 12'h555;
rom[59500] = 12'h555;
rom[59501] = 12'h555;
rom[59502] = 12'h555;
rom[59503] = 12'h555;
rom[59504] = 12'h666;
rom[59505] = 12'h666;
rom[59506] = 12'h666;
rom[59507] = 12'h666;
rom[59508] = 12'h666;
rom[59509] = 12'h666;
rom[59510] = 12'h555;
rom[59511] = 12'h555;
rom[59512] = 12'h555;
rom[59513] = 12'h555;
rom[59514] = 12'h555;
rom[59515] = 12'h555;
rom[59516] = 12'h555;
rom[59517] = 12'h555;
rom[59518] = 12'h555;
rom[59519] = 12'h555;
rom[59520] = 12'h666;
rom[59521] = 12'h666;
rom[59522] = 12'h666;
rom[59523] = 12'h666;
rom[59524] = 12'h666;
rom[59525] = 12'h666;
rom[59526] = 12'h666;
rom[59527] = 12'h666;
rom[59528] = 12'h777;
rom[59529] = 12'h777;
rom[59530] = 12'h777;
rom[59531] = 12'h777;
rom[59532] = 12'h777;
rom[59533] = 12'h777;
rom[59534] = 12'h777;
rom[59535] = 12'h777;
rom[59536] = 12'h777;
rom[59537] = 12'h777;
rom[59538] = 12'h888;
rom[59539] = 12'h888;
rom[59540] = 12'h888;
rom[59541] = 12'h999;
rom[59542] = 12'h999;
rom[59543] = 12'h999;
rom[59544] = 12'h999;
rom[59545] = 12'haaa;
rom[59546] = 12'haaa;
rom[59547] = 12'haaa;
rom[59548] = 12'haaa;
rom[59549] = 12'hbbb;
rom[59550] = 12'hbbb;
rom[59551] = 12'hbbb;
rom[59552] = 12'hbbb;
rom[59553] = 12'hccc;
rom[59554] = 12'hccc;
rom[59555] = 12'hddd;
rom[59556] = 12'heee;
rom[59557] = 12'heee;
rom[59558] = 12'hfff;
rom[59559] = 12'hfff;
rom[59560] = 12'heee;
rom[59561] = 12'heee;
rom[59562] = 12'hddd;
rom[59563] = 12'hccc;
rom[59564] = 12'hccc;
rom[59565] = 12'hccc;
rom[59566] = 12'hbbb;
rom[59567] = 12'hbbb;
rom[59568] = 12'hbbb;
rom[59569] = 12'hbbb;
rom[59570] = 12'hbbb;
rom[59571] = 12'hbbb;
rom[59572] = 12'haaa;
rom[59573] = 12'haaa;
rom[59574] = 12'haaa;
rom[59575] = 12'haaa;
rom[59576] = 12'haaa;
rom[59577] = 12'h999;
rom[59578] = 12'h999;
rom[59579] = 12'h999;
rom[59580] = 12'h999;
rom[59581] = 12'h999;
rom[59582] = 12'h888;
rom[59583] = 12'h888;
rom[59584] = 12'h888;
rom[59585] = 12'h888;
rom[59586] = 12'h888;
rom[59587] = 12'h888;
rom[59588] = 12'h888;
rom[59589] = 12'h888;
rom[59590] = 12'h888;
rom[59591] = 12'h888;
rom[59592] = 12'h888;
rom[59593] = 12'h888;
rom[59594] = 12'h888;
rom[59595] = 12'h888;
rom[59596] = 12'h888;
rom[59597] = 12'h888;
rom[59598] = 12'h888;
rom[59599] = 12'h888;
rom[59600] = 12'hfff;
rom[59601] = 12'hfff;
rom[59602] = 12'hfff;
rom[59603] = 12'hfff;
rom[59604] = 12'hfff;
rom[59605] = 12'hfff;
rom[59606] = 12'hfff;
rom[59607] = 12'hfff;
rom[59608] = 12'hfff;
rom[59609] = 12'hfff;
rom[59610] = 12'hfff;
rom[59611] = 12'hfff;
rom[59612] = 12'hfff;
rom[59613] = 12'hfff;
rom[59614] = 12'hfff;
rom[59615] = 12'hfff;
rom[59616] = 12'hfff;
rom[59617] = 12'hfff;
rom[59618] = 12'hfff;
rom[59619] = 12'hfff;
rom[59620] = 12'hfff;
rom[59621] = 12'hfff;
rom[59622] = 12'hfff;
rom[59623] = 12'hfff;
rom[59624] = 12'hfff;
rom[59625] = 12'hfff;
rom[59626] = 12'hfff;
rom[59627] = 12'hfff;
rom[59628] = 12'hfff;
rom[59629] = 12'hfff;
rom[59630] = 12'hfff;
rom[59631] = 12'hfff;
rom[59632] = 12'hfff;
rom[59633] = 12'hfff;
rom[59634] = 12'hfff;
rom[59635] = 12'hfff;
rom[59636] = 12'hfff;
rom[59637] = 12'hfff;
rom[59638] = 12'hfff;
rom[59639] = 12'hfff;
rom[59640] = 12'hfff;
rom[59641] = 12'hfff;
rom[59642] = 12'hfff;
rom[59643] = 12'hfff;
rom[59644] = 12'hfff;
rom[59645] = 12'hfff;
rom[59646] = 12'hfff;
rom[59647] = 12'hfff;
rom[59648] = 12'hfff;
rom[59649] = 12'hfff;
rom[59650] = 12'hfff;
rom[59651] = 12'hfff;
rom[59652] = 12'hfff;
rom[59653] = 12'hfff;
rom[59654] = 12'hfff;
rom[59655] = 12'hfff;
rom[59656] = 12'hfff;
rom[59657] = 12'hfff;
rom[59658] = 12'hfff;
rom[59659] = 12'hfff;
rom[59660] = 12'hfff;
rom[59661] = 12'hfff;
rom[59662] = 12'hfff;
rom[59663] = 12'hfff;
rom[59664] = 12'hfff;
rom[59665] = 12'hfff;
rom[59666] = 12'hfff;
rom[59667] = 12'hfff;
rom[59668] = 12'hfff;
rom[59669] = 12'hfff;
rom[59670] = 12'hfff;
rom[59671] = 12'hfff;
rom[59672] = 12'hfff;
rom[59673] = 12'hfff;
rom[59674] = 12'hfff;
rom[59675] = 12'hfff;
rom[59676] = 12'hfff;
rom[59677] = 12'hfff;
rom[59678] = 12'hfff;
rom[59679] = 12'hfff;
rom[59680] = 12'hfff;
rom[59681] = 12'hfff;
rom[59682] = 12'hfff;
rom[59683] = 12'hfff;
rom[59684] = 12'hfff;
rom[59685] = 12'hfff;
rom[59686] = 12'hfff;
rom[59687] = 12'hfff;
rom[59688] = 12'hfff;
rom[59689] = 12'hfff;
rom[59690] = 12'hfff;
rom[59691] = 12'hfff;
rom[59692] = 12'hfff;
rom[59693] = 12'heee;
rom[59694] = 12'heee;
rom[59695] = 12'heee;
rom[59696] = 12'hddd;
rom[59697] = 12'hddd;
rom[59698] = 12'hddd;
rom[59699] = 12'hddd;
rom[59700] = 12'hddd;
rom[59701] = 12'hccc;
rom[59702] = 12'hccc;
rom[59703] = 12'hccc;
rom[59704] = 12'hccc;
rom[59705] = 12'hccc;
rom[59706] = 12'hccc;
rom[59707] = 12'hccc;
rom[59708] = 12'hccc;
rom[59709] = 12'hccc;
rom[59710] = 12'hccc;
rom[59711] = 12'hbbb;
rom[59712] = 12'hbbb;
rom[59713] = 12'hccc;
rom[59714] = 12'hccc;
rom[59715] = 12'hccc;
rom[59716] = 12'hccc;
rom[59717] = 12'hccc;
rom[59718] = 12'hccc;
rom[59719] = 12'hccc;
rom[59720] = 12'hccc;
rom[59721] = 12'hccc;
rom[59722] = 12'hbbb;
rom[59723] = 12'hbbb;
rom[59724] = 12'hbbb;
rom[59725] = 12'haaa;
rom[59726] = 12'haaa;
rom[59727] = 12'haaa;
rom[59728] = 12'h999;
rom[59729] = 12'h888;
rom[59730] = 12'h888;
rom[59731] = 12'h777;
rom[59732] = 12'h777;
rom[59733] = 12'h777;
rom[59734] = 12'h777;
rom[59735] = 12'h777;
rom[59736] = 12'h777;
rom[59737] = 12'h777;
rom[59738] = 12'h666;
rom[59739] = 12'h666;
rom[59740] = 12'h555;
rom[59741] = 12'h555;
rom[59742] = 12'h444;
rom[59743] = 12'h444;
rom[59744] = 12'h444;
rom[59745] = 12'h333;
rom[59746] = 12'h333;
rom[59747] = 12'h333;
rom[59748] = 12'h333;
rom[59749] = 12'h333;
rom[59750] = 12'h333;
rom[59751] = 12'h222;
rom[59752] = 12'h222;
rom[59753] = 12'h222;
rom[59754] = 12'h222;
rom[59755] = 12'h222;
rom[59756] = 12'h222;
rom[59757] = 12'h222;
rom[59758] = 12'h222;
rom[59759] = 12'h222;
rom[59760] = 12'h222;
rom[59761] = 12'h222;
rom[59762] = 12'h222;
rom[59763] = 12'h222;
rom[59764] = 12'h222;
rom[59765] = 12'h222;
rom[59766] = 12'h222;
rom[59767] = 12'h222;
rom[59768] = 12'h222;
rom[59769] = 12'h222;
rom[59770] = 12'h222;
rom[59771] = 12'h222;
rom[59772] = 12'h111;
rom[59773] = 12'h111;
rom[59774] = 12'h  0;
rom[59775] = 12'h  0;
rom[59776] = 12'h  0;
rom[59777] = 12'h  0;
rom[59778] = 12'h  0;
rom[59779] = 12'h  0;
rom[59780] = 12'h  0;
rom[59781] = 12'h  0;
rom[59782] = 12'h  0;
rom[59783] = 12'h  0;
rom[59784] = 12'h  0;
rom[59785] = 12'h  0;
rom[59786] = 12'h  0;
rom[59787] = 12'h  0;
rom[59788] = 12'h  0;
rom[59789] = 12'h  0;
rom[59790] = 12'h  0;
rom[59791] = 12'h  0;
rom[59792] = 12'h  0;
rom[59793] = 12'h  0;
rom[59794] = 12'h  0;
rom[59795] = 12'h  0;
rom[59796] = 12'h  0;
rom[59797] = 12'h  0;
rom[59798] = 12'h  0;
rom[59799] = 12'h  0;
rom[59800] = 12'h  0;
rom[59801] = 12'h  0;
rom[59802] = 12'h  0;
rom[59803] = 12'h  0;
rom[59804] = 12'h111;
rom[59805] = 12'h111;
rom[59806] = 12'h111;
rom[59807] = 12'h111;
rom[59808] = 12'h111;
rom[59809] = 12'h111;
rom[59810] = 12'h111;
rom[59811] = 12'h111;
rom[59812] = 12'h111;
rom[59813] = 12'h111;
rom[59814] = 12'h222;
rom[59815] = 12'h222;
rom[59816] = 12'h222;
rom[59817] = 12'h222;
rom[59818] = 12'h111;
rom[59819] = 12'h111;
rom[59820] = 12'h111;
rom[59821] = 12'h111;
rom[59822] = 12'h111;
rom[59823] = 12'h111;
rom[59824] = 12'h111;
rom[59825] = 12'h  0;
rom[59826] = 12'h  0;
rom[59827] = 12'h  0;
rom[59828] = 12'h  0;
rom[59829] = 12'h  0;
rom[59830] = 12'h  0;
rom[59831] = 12'h  0;
rom[59832] = 12'h  0;
rom[59833] = 12'h  0;
rom[59834] = 12'h  0;
rom[59835] = 12'h  0;
rom[59836] = 12'h  0;
rom[59837] = 12'h  0;
rom[59838] = 12'h  0;
rom[59839] = 12'h  0;
rom[59840] = 12'h  0;
rom[59841] = 12'h  0;
rom[59842] = 12'h  0;
rom[59843] = 12'h  0;
rom[59844] = 12'h  0;
rom[59845] = 12'h  0;
rom[59846] = 12'h  0;
rom[59847] = 12'h  0;
rom[59848] = 12'h  0;
rom[59849] = 12'h  0;
rom[59850] = 12'h  0;
rom[59851] = 12'h  0;
rom[59852] = 12'h  0;
rom[59853] = 12'h  0;
rom[59854] = 12'h  0;
rom[59855] = 12'h  0;
rom[59856] = 12'h  0;
rom[59857] = 12'h  0;
rom[59858] = 12'h  0;
rom[59859] = 12'h  0;
rom[59860] = 12'h  0;
rom[59861] = 12'h  0;
rom[59862] = 12'h  0;
rom[59863] = 12'h  0;
rom[59864] = 12'h  0;
rom[59865] = 12'h  0;
rom[59866] = 12'h  0;
rom[59867] = 12'h  0;
rom[59868] = 12'h  0;
rom[59869] = 12'h  0;
rom[59870] = 12'h  0;
rom[59871] = 12'h  0;
rom[59872] = 12'h111;
rom[59873] = 12'h111;
rom[59874] = 12'h111;
rom[59875] = 12'h222;
rom[59876] = 12'h222;
rom[59877] = 12'h333;
rom[59878] = 12'h333;
rom[59879] = 12'h333;
rom[59880] = 12'h444;
rom[59881] = 12'h444;
rom[59882] = 12'h555;
rom[59883] = 12'h555;
rom[59884] = 12'h333;
rom[59885] = 12'h222;
rom[59886] = 12'h222;
rom[59887] = 12'h222;
rom[59888] = 12'h222;
rom[59889] = 12'h222;
rom[59890] = 12'h222;
rom[59891] = 12'h222;
rom[59892] = 12'h222;
rom[59893] = 12'h222;
rom[59894] = 12'h333;
rom[59895] = 12'h333;
rom[59896] = 12'h333;
rom[59897] = 12'h555;
rom[59898] = 12'h555;
rom[59899] = 12'h555;
rom[59900] = 12'h555;
rom[59901] = 12'h555;
rom[59902] = 12'h555;
rom[59903] = 12'h555;
rom[59904] = 12'h555;
rom[59905] = 12'h666;
rom[59906] = 12'h666;
rom[59907] = 12'h666;
rom[59908] = 12'h666;
rom[59909] = 12'h666;
rom[59910] = 12'h555;
rom[59911] = 12'h555;
rom[59912] = 12'h555;
rom[59913] = 12'h555;
rom[59914] = 12'h555;
rom[59915] = 12'h555;
rom[59916] = 12'h555;
rom[59917] = 12'h555;
rom[59918] = 12'h555;
rom[59919] = 12'h555;
rom[59920] = 12'h666;
rom[59921] = 12'h666;
rom[59922] = 12'h666;
rom[59923] = 12'h666;
rom[59924] = 12'h666;
rom[59925] = 12'h666;
rom[59926] = 12'h777;
rom[59927] = 12'h777;
rom[59928] = 12'h777;
rom[59929] = 12'h777;
rom[59930] = 12'h777;
rom[59931] = 12'h777;
rom[59932] = 12'h777;
rom[59933] = 12'h777;
rom[59934] = 12'h777;
rom[59935] = 12'h777;
rom[59936] = 12'h888;
rom[59937] = 12'h888;
rom[59938] = 12'h888;
rom[59939] = 12'h888;
rom[59940] = 12'h999;
rom[59941] = 12'h999;
rom[59942] = 12'h999;
rom[59943] = 12'h999;
rom[59944] = 12'haaa;
rom[59945] = 12'haaa;
rom[59946] = 12'haaa;
rom[59947] = 12'haaa;
rom[59948] = 12'hbbb;
rom[59949] = 12'hbbb;
rom[59950] = 12'hbbb;
rom[59951] = 12'hbbb;
rom[59952] = 12'hccc;
rom[59953] = 12'hccc;
rom[59954] = 12'hddd;
rom[59955] = 12'hddd;
rom[59956] = 12'heee;
rom[59957] = 12'hfff;
rom[59958] = 12'hfff;
rom[59959] = 12'hfff;
rom[59960] = 12'heee;
rom[59961] = 12'hddd;
rom[59962] = 12'hccc;
rom[59963] = 12'hccc;
rom[59964] = 12'hccc;
rom[59965] = 12'hccc;
rom[59966] = 12'hbbb;
rom[59967] = 12'hbbb;
rom[59968] = 12'hbbb;
rom[59969] = 12'hbbb;
rom[59970] = 12'hbbb;
rom[59971] = 12'hbbb;
rom[59972] = 12'haaa;
rom[59973] = 12'haaa;
rom[59974] = 12'haaa;
rom[59975] = 12'haaa;
rom[59976] = 12'h999;
rom[59977] = 12'h999;
rom[59978] = 12'h999;
rom[59979] = 12'h999;
rom[59980] = 12'h999;
rom[59981] = 12'h999;
rom[59982] = 12'h888;
rom[59983] = 12'h888;
rom[59984] = 12'h888;
rom[59985] = 12'h888;
rom[59986] = 12'h888;
rom[59987] = 12'h888;
rom[59988] = 12'h888;
rom[59989] = 12'h888;
rom[59990] = 12'h888;
rom[59991] = 12'h888;
rom[59992] = 12'h888;
rom[59993] = 12'h888;
rom[59994] = 12'h888;
rom[59995] = 12'h888;
rom[59996] = 12'h888;
rom[59997] = 12'h888;
rom[59998] = 12'h888;
rom[59999] = 12'h888;
rom[60000] = 12'hfff;
rom[60001] = 12'hfff;
rom[60002] = 12'hfff;
rom[60003] = 12'hfff;
rom[60004] = 12'hfff;
rom[60005] = 12'hfff;
rom[60006] = 12'hfff;
rom[60007] = 12'hfff;
rom[60008] = 12'hfff;
rom[60009] = 12'hfff;
rom[60010] = 12'hfff;
rom[60011] = 12'hfff;
rom[60012] = 12'hfff;
rom[60013] = 12'hfff;
rom[60014] = 12'hfff;
rom[60015] = 12'hfff;
rom[60016] = 12'hfff;
rom[60017] = 12'hfff;
rom[60018] = 12'hfff;
rom[60019] = 12'hfff;
rom[60020] = 12'hfff;
rom[60021] = 12'hfff;
rom[60022] = 12'hfff;
rom[60023] = 12'hfff;
rom[60024] = 12'hfff;
rom[60025] = 12'hfff;
rom[60026] = 12'hfff;
rom[60027] = 12'hfff;
rom[60028] = 12'hfff;
rom[60029] = 12'hfff;
rom[60030] = 12'hfff;
rom[60031] = 12'hfff;
rom[60032] = 12'hfff;
rom[60033] = 12'hfff;
rom[60034] = 12'hfff;
rom[60035] = 12'hfff;
rom[60036] = 12'hfff;
rom[60037] = 12'hfff;
rom[60038] = 12'hfff;
rom[60039] = 12'hfff;
rom[60040] = 12'hfff;
rom[60041] = 12'hfff;
rom[60042] = 12'hfff;
rom[60043] = 12'hfff;
rom[60044] = 12'hfff;
rom[60045] = 12'hfff;
rom[60046] = 12'hfff;
rom[60047] = 12'hfff;
rom[60048] = 12'hfff;
rom[60049] = 12'hfff;
rom[60050] = 12'hfff;
rom[60051] = 12'hfff;
rom[60052] = 12'hfff;
rom[60053] = 12'hfff;
rom[60054] = 12'hfff;
rom[60055] = 12'hfff;
rom[60056] = 12'hfff;
rom[60057] = 12'hfff;
rom[60058] = 12'hfff;
rom[60059] = 12'hfff;
rom[60060] = 12'hfff;
rom[60061] = 12'hfff;
rom[60062] = 12'hfff;
rom[60063] = 12'hfff;
rom[60064] = 12'hfff;
rom[60065] = 12'hfff;
rom[60066] = 12'hfff;
rom[60067] = 12'hfff;
rom[60068] = 12'hfff;
rom[60069] = 12'hfff;
rom[60070] = 12'hfff;
rom[60071] = 12'hfff;
rom[60072] = 12'hfff;
rom[60073] = 12'hfff;
rom[60074] = 12'hfff;
rom[60075] = 12'hfff;
rom[60076] = 12'hfff;
rom[60077] = 12'hfff;
rom[60078] = 12'hfff;
rom[60079] = 12'hfff;
rom[60080] = 12'hfff;
rom[60081] = 12'hfff;
rom[60082] = 12'hfff;
rom[60083] = 12'hfff;
rom[60084] = 12'hfff;
rom[60085] = 12'hfff;
rom[60086] = 12'hfff;
rom[60087] = 12'hfff;
rom[60088] = 12'hfff;
rom[60089] = 12'hfff;
rom[60090] = 12'hfff;
rom[60091] = 12'hfff;
rom[60092] = 12'hfff;
rom[60093] = 12'hfff;
rom[60094] = 12'hfff;
rom[60095] = 12'heee;
rom[60096] = 12'heee;
rom[60097] = 12'heee;
rom[60098] = 12'hddd;
rom[60099] = 12'hddd;
rom[60100] = 12'hddd;
rom[60101] = 12'hddd;
rom[60102] = 12'hddd;
rom[60103] = 12'hccc;
rom[60104] = 12'hccc;
rom[60105] = 12'hccc;
rom[60106] = 12'hccc;
rom[60107] = 12'hccc;
rom[60108] = 12'hccc;
rom[60109] = 12'hccc;
rom[60110] = 12'hccc;
rom[60111] = 12'hccc;
rom[60112] = 12'hbbb;
rom[60113] = 12'hbbb;
rom[60114] = 12'hbbb;
rom[60115] = 12'hccc;
rom[60116] = 12'hccc;
rom[60117] = 12'hccc;
rom[60118] = 12'hccc;
rom[60119] = 12'hccc;
rom[60120] = 12'hccc;
rom[60121] = 12'hbbb;
rom[60122] = 12'hbbb;
rom[60123] = 12'hbbb;
rom[60124] = 12'hbbb;
rom[60125] = 12'hbbb;
rom[60126] = 12'hbbb;
rom[60127] = 12'hbbb;
rom[60128] = 12'haaa;
rom[60129] = 12'haaa;
rom[60130] = 12'h999;
rom[60131] = 12'h999;
rom[60132] = 12'h888;
rom[60133] = 12'h888;
rom[60134] = 12'h777;
rom[60135] = 12'h777;
rom[60136] = 12'h777;
rom[60137] = 12'h777;
rom[60138] = 12'h777;
rom[60139] = 12'h666;
rom[60140] = 12'h666;
rom[60141] = 12'h555;
rom[60142] = 12'h555;
rom[60143] = 12'h444;
rom[60144] = 12'h444;
rom[60145] = 12'h444;
rom[60146] = 12'h333;
rom[60147] = 12'h333;
rom[60148] = 12'h333;
rom[60149] = 12'h333;
rom[60150] = 12'h333;
rom[60151] = 12'h333;
rom[60152] = 12'h222;
rom[60153] = 12'h222;
rom[60154] = 12'h222;
rom[60155] = 12'h222;
rom[60156] = 12'h222;
rom[60157] = 12'h222;
rom[60158] = 12'h222;
rom[60159] = 12'h222;
rom[60160] = 12'h222;
rom[60161] = 12'h222;
rom[60162] = 12'h222;
rom[60163] = 12'h222;
rom[60164] = 12'h222;
rom[60165] = 12'h222;
rom[60166] = 12'h222;
rom[60167] = 12'h222;
rom[60168] = 12'h222;
rom[60169] = 12'h222;
rom[60170] = 12'h111;
rom[60171] = 12'h111;
rom[60172] = 12'h111;
rom[60173] = 12'h  0;
rom[60174] = 12'h  0;
rom[60175] = 12'h  0;
rom[60176] = 12'h  0;
rom[60177] = 12'h  0;
rom[60178] = 12'h  0;
rom[60179] = 12'h  0;
rom[60180] = 12'h  0;
rom[60181] = 12'h  0;
rom[60182] = 12'h  0;
rom[60183] = 12'h  0;
rom[60184] = 12'h  0;
rom[60185] = 12'h  0;
rom[60186] = 12'h  0;
rom[60187] = 12'h  0;
rom[60188] = 12'h  0;
rom[60189] = 12'h  0;
rom[60190] = 12'h  0;
rom[60191] = 12'h  0;
rom[60192] = 12'h  0;
rom[60193] = 12'h  0;
rom[60194] = 12'h  0;
rom[60195] = 12'h  0;
rom[60196] = 12'h  0;
rom[60197] = 12'h  0;
rom[60198] = 12'h  0;
rom[60199] = 12'h  0;
rom[60200] = 12'h  0;
rom[60201] = 12'h  0;
rom[60202] = 12'h  0;
rom[60203] = 12'h111;
rom[60204] = 12'h111;
rom[60205] = 12'h111;
rom[60206] = 12'h111;
rom[60207] = 12'h111;
rom[60208] = 12'h111;
rom[60209] = 12'h111;
rom[60210] = 12'h111;
rom[60211] = 12'h111;
rom[60212] = 12'h111;
rom[60213] = 12'h222;
rom[60214] = 12'h222;
rom[60215] = 12'h222;
rom[60216] = 12'h222;
rom[60217] = 12'h222;
rom[60218] = 12'h111;
rom[60219] = 12'h111;
rom[60220] = 12'h111;
rom[60221] = 12'h111;
rom[60222] = 12'h111;
rom[60223] = 12'h111;
rom[60224] = 12'h  0;
rom[60225] = 12'h  0;
rom[60226] = 12'h  0;
rom[60227] = 12'h  0;
rom[60228] = 12'h  0;
rom[60229] = 12'h  0;
rom[60230] = 12'h  0;
rom[60231] = 12'h  0;
rom[60232] = 12'h  0;
rom[60233] = 12'h  0;
rom[60234] = 12'h  0;
rom[60235] = 12'h  0;
rom[60236] = 12'h  0;
rom[60237] = 12'h  0;
rom[60238] = 12'h  0;
rom[60239] = 12'h  0;
rom[60240] = 12'h  0;
rom[60241] = 12'h  0;
rom[60242] = 12'h  0;
rom[60243] = 12'h  0;
rom[60244] = 12'h  0;
rom[60245] = 12'h  0;
rom[60246] = 12'h  0;
rom[60247] = 12'h  0;
rom[60248] = 12'h  0;
rom[60249] = 12'h  0;
rom[60250] = 12'h  0;
rom[60251] = 12'h  0;
rom[60252] = 12'h  0;
rom[60253] = 12'h  0;
rom[60254] = 12'h  0;
rom[60255] = 12'h  0;
rom[60256] = 12'h  0;
rom[60257] = 12'h  0;
rom[60258] = 12'h  0;
rom[60259] = 12'h  0;
rom[60260] = 12'h  0;
rom[60261] = 12'h  0;
rom[60262] = 12'h  0;
rom[60263] = 12'h  0;
rom[60264] = 12'h  0;
rom[60265] = 12'h  0;
rom[60266] = 12'h  0;
rom[60267] = 12'h  0;
rom[60268] = 12'h  0;
rom[60269] = 12'h  0;
rom[60270] = 12'h  0;
rom[60271] = 12'h  0;
rom[60272] = 12'h  0;
rom[60273] = 12'h111;
rom[60274] = 12'h111;
rom[60275] = 12'h222;
rom[60276] = 12'h222;
rom[60277] = 12'h333;
rom[60278] = 12'h333;
rom[60279] = 12'h333;
rom[60280] = 12'h444;
rom[60281] = 12'h444;
rom[60282] = 12'h555;
rom[60283] = 12'h444;
rom[60284] = 12'h333;
rom[60285] = 12'h222;
rom[60286] = 12'h222;
rom[60287] = 12'h222;
rom[60288] = 12'h222;
rom[60289] = 12'h222;
rom[60290] = 12'h222;
rom[60291] = 12'h222;
rom[60292] = 12'h222;
rom[60293] = 12'h222;
rom[60294] = 12'h333;
rom[60295] = 12'h333;
rom[60296] = 12'h333;
rom[60297] = 12'h444;
rom[60298] = 12'h555;
rom[60299] = 12'h555;
rom[60300] = 12'h555;
rom[60301] = 12'h444;
rom[60302] = 12'h555;
rom[60303] = 12'h555;
rom[60304] = 12'h555;
rom[60305] = 12'h555;
rom[60306] = 12'h555;
rom[60307] = 12'h666;
rom[60308] = 12'h666;
rom[60309] = 12'h666;
rom[60310] = 12'h666;
rom[60311] = 12'h666;
rom[60312] = 12'h555;
rom[60313] = 12'h555;
rom[60314] = 12'h555;
rom[60315] = 12'h555;
rom[60316] = 12'h555;
rom[60317] = 12'h555;
rom[60318] = 12'h555;
rom[60319] = 12'h666;
rom[60320] = 12'h666;
rom[60321] = 12'h666;
rom[60322] = 12'h666;
rom[60323] = 12'h666;
rom[60324] = 12'h666;
rom[60325] = 12'h777;
rom[60326] = 12'h777;
rom[60327] = 12'h777;
rom[60328] = 12'h777;
rom[60329] = 12'h777;
rom[60330] = 12'h777;
rom[60331] = 12'h777;
rom[60332] = 12'h777;
rom[60333] = 12'h888;
rom[60334] = 12'h888;
rom[60335] = 12'h888;
rom[60336] = 12'h888;
rom[60337] = 12'h888;
rom[60338] = 12'h888;
rom[60339] = 12'h999;
rom[60340] = 12'h999;
rom[60341] = 12'h999;
rom[60342] = 12'h999;
rom[60343] = 12'haaa;
rom[60344] = 12'haaa;
rom[60345] = 12'haaa;
rom[60346] = 12'haaa;
rom[60347] = 12'hbbb;
rom[60348] = 12'hbbb;
rom[60349] = 12'hbbb;
rom[60350] = 12'hbbb;
rom[60351] = 12'hccc;
rom[60352] = 12'hccc;
rom[60353] = 12'hccc;
rom[60354] = 12'hddd;
rom[60355] = 12'heee;
rom[60356] = 12'hfff;
rom[60357] = 12'hfff;
rom[60358] = 12'hfff;
rom[60359] = 12'heee;
rom[60360] = 12'heee;
rom[60361] = 12'hddd;
rom[60362] = 12'hccc;
rom[60363] = 12'hccc;
rom[60364] = 12'hccc;
rom[60365] = 12'hbbb;
rom[60366] = 12'hbbb;
rom[60367] = 12'hbbb;
rom[60368] = 12'hbbb;
rom[60369] = 12'hbbb;
rom[60370] = 12'hbbb;
rom[60371] = 12'hbbb;
rom[60372] = 12'hbbb;
rom[60373] = 12'haaa;
rom[60374] = 12'haaa;
rom[60375] = 12'haaa;
rom[60376] = 12'h999;
rom[60377] = 12'h999;
rom[60378] = 12'h999;
rom[60379] = 12'h999;
rom[60380] = 12'h999;
rom[60381] = 12'h999;
rom[60382] = 12'h999;
rom[60383] = 12'h999;
rom[60384] = 12'h888;
rom[60385] = 12'h888;
rom[60386] = 12'h888;
rom[60387] = 12'h888;
rom[60388] = 12'h888;
rom[60389] = 12'h888;
rom[60390] = 12'h888;
rom[60391] = 12'h888;
rom[60392] = 12'h888;
rom[60393] = 12'h888;
rom[60394] = 12'h888;
rom[60395] = 12'h888;
rom[60396] = 12'h888;
rom[60397] = 12'h888;
rom[60398] = 12'h888;
rom[60399] = 12'h888;
rom[60400] = 12'hfff;
rom[60401] = 12'hfff;
rom[60402] = 12'hfff;
rom[60403] = 12'hfff;
rom[60404] = 12'hfff;
rom[60405] = 12'hfff;
rom[60406] = 12'hfff;
rom[60407] = 12'hfff;
rom[60408] = 12'hfff;
rom[60409] = 12'hfff;
rom[60410] = 12'hfff;
rom[60411] = 12'hfff;
rom[60412] = 12'hfff;
rom[60413] = 12'hfff;
rom[60414] = 12'hfff;
rom[60415] = 12'hfff;
rom[60416] = 12'hfff;
rom[60417] = 12'hfff;
rom[60418] = 12'hfff;
rom[60419] = 12'hfff;
rom[60420] = 12'hfff;
rom[60421] = 12'hfff;
rom[60422] = 12'hfff;
rom[60423] = 12'hfff;
rom[60424] = 12'hfff;
rom[60425] = 12'hfff;
rom[60426] = 12'hfff;
rom[60427] = 12'hfff;
rom[60428] = 12'hfff;
rom[60429] = 12'hfff;
rom[60430] = 12'hfff;
rom[60431] = 12'hfff;
rom[60432] = 12'hfff;
rom[60433] = 12'hfff;
rom[60434] = 12'hfff;
rom[60435] = 12'hfff;
rom[60436] = 12'hfff;
rom[60437] = 12'hfff;
rom[60438] = 12'hfff;
rom[60439] = 12'hfff;
rom[60440] = 12'hfff;
rom[60441] = 12'hfff;
rom[60442] = 12'hfff;
rom[60443] = 12'hfff;
rom[60444] = 12'hfff;
rom[60445] = 12'hfff;
rom[60446] = 12'hfff;
rom[60447] = 12'hfff;
rom[60448] = 12'hfff;
rom[60449] = 12'hfff;
rom[60450] = 12'hfff;
rom[60451] = 12'hfff;
rom[60452] = 12'hfff;
rom[60453] = 12'hfff;
rom[60454] = 12'hfff;
rom[60455] = 12'hfff;
rom[60456] = 12'hfff;
rom[60457] = 12'hfff;
rom[60458] = 12'hfff;
rom[60459] = 12'hfff;
rom[60460] = 12'hfff;
rom[60461] = 12'hfff;
rom[60462] = 12'hfff;
rom[60463] = 12'hfff;
rom[60464] = 12'hfff;
rom[60465] = 12'hfff;
rom[60466] = 12'hfff;
rom[60467] = 12'hfff;
rom[60468] = 12'hfff;
rom[60469] = 12'hfff;
rom[60470] = 12'hfff;
rom[60471] = 12'hfff;
rom[60472] = 12'hfff;
rom[60473] = 12'hfff;
rom[60474] = 12'hfff;
rom[60475] = 12'hfff;
rom[60476] = 12'hfff;
rom[60477] = 12'hfff;
rom[60478] = 12'hfff;
rom[60479] = 12'hfff;
rom[60480] = 12'hfff;
rom[60481] = 12'hfff;
rom[60482] = 12'hfff;
rom[60483] = 12'hfff;
rom[60484] = 12'hfff;
rom[60485] = 12'hfff;
rom[60486] = 12'hfff;
rom[60487] = 12'hfff;
rom[60488] = 12'hfff;
rom[60489] = 12'hfff;
rom[60490] = 12'hfff;
rom[60491] = 12'hfff;
rom[60492] = 12'hfff;
rom[60493] = 12'hfff;
rom[60494] = 12'hfff;
rom[60495] = 12'hfff;
rom[60496] = 12'heee;
rom[60497] = 12'heee;
rom[60498] = 12'heee;
rom[60499] = 12'heee;
rom[60500] = 12'heee;
rom[60501] = 12'hddd;
rom[60502] = 12'hddd;
rom[60503] = 12'hddd;
rom[60504] = 12'hddd;
rom[60505] = 12'hddd;
rom[60506] = 12'hccc;
rom[60507] = 12'hccc;
rom[60508] = 12'hccc;
rom[60509] = 12'hccc;
rom[60510] = 12'hccc;
rom[60511] = 12'hccc;
rom[60512] = 12'hccc;
rom[60513] = 12'hccc;
rom[60514] = 12'hbbb;
rom[60515] = 12'hbbb;
rom[60516] = 12'hccc;
rom[60517] = 12'hccc;
rom[60518] = 12'hccc;
rom[60519] = 12'hbbb;
rom[60520] = 12'hbbb;
rom[60521] = 12'hbbb;
rom[60522] = 12'hbbb;
rom[60523] = 12'hbbb;
rom[60524] = 12'hbbb;
rom[60525] = 12'hbbb;
rom[60526] = 12'hbbb;
rom[60527] = 12'hbbb;
rom[60528] = 12'hbbb;
rom[60529] = 12'hbbb;
rom[60530] = 12'haaa;
rom[60531] = 12'haaa;
rom[60532] = 12'haaa;
rom[60533] = 12'h999;
rom[60534] = 12'h999;
rom[60535] = 12'h888;
rom[60536] = 12'h777;
rom[60537] = 12'h777;
rom[60538] = 12'h777;
rom[60539] = 12'h777;
rom[60540] = 12'h666;
rom[60541] = 12'h666;
rom[60542] = 12'h555;
rom[60543] = 12'h555;
rom[60544] = 12'h444;
rom[60545] = 12'h444;
rom[60546] = 12'h444;
rom[60547] = 12'h333;
rom[60548] = 12'h333;
rom[60549] = 12'h333;
rom[60550] = 12'h333;
rom[60551] = 12'h333;
rom[60552] = 12'h222;
rom[60553] = 12'h222;
rom[60554] = 12'h222;
rom[60555] = 12'h333;
rom[60556] = 12'h333;
rom[60557] = 12'h333;
rom[60558] = 12'h333;
rom[60559] = 12'h333;
rom[60560] = 12'h222;
rom[60561] = 12'h222;
rom[60562] = 12'h222;
rom[60563] = 12'h222;
rom[60564] = 12'h222;
rom[60565] = 12'h222;
rom[60566] = 12'h222;
rom[60567] = 12'h222;
rom[60568] = 12'h222;
rom[60569] = 12'h111;
rom[60570] = 12'h111;
rom[60571] = 12'h111;
rom[60572] = 12'h  0;
rom[60573] = 12'h  0;
rom[60574] = 12'h  0;
rom[60575] = 12'h  0;
rom[60576] = 12'h  0;
rom[60577] = 12'h  0;
rom[60578] = 12'h  0;
rom[60579] = 12'h  0;
rom[60580] = 12'h  0;
rom[60581] = 12'h  0;
rom[60582] = 12'h  0;
rom[60583] = 12'h  0;
rom[60584] = 12'h  0;
rom[60585] = 12'h  0;
rom[60586] = 12'h  0;
rom[60587] = 12'h  0;
rom[60588] = 12'h  0;
rom[60589] = 12'h  0;
rom[60590] = 12'h  0;
rom[60591] = 12'h  0;
rom[60592] = 12'h  0;
rom[60593] = 12'h  0;
rom[60594] = 12'h  0;
rom[60595] = 12'h  0;
rom[60596] = 12'h  0;
rom[60597] = 12'h  0;
rom[60598] = 12'h  0;
rom[60599] = 12'h  0;
rom[60600] = 12'h  0;
rom[60601] = 12'h  0;
rom[60602] = 12'h111;
rom[60603] = 12'h111;
rom[60604] = 12'h111;
rom[60605] = 12'h111;
rom[60606] = 12'h111;
rom[60607] = 12'h111;
rom[60608] = 12'h111;
rom[60609] = 12'h111;
rom[60610] = 12'h111;
rom[60611] = 12'h111;
rom[60612] = 12'h111;
rom[60613] = 12'h222;
rom[60614] = 12'h222;
rom[60615] = 12'h222;
rom[60616] = 12'h222;
rom[60617] = 12'h111;
rom[60618] = 12'h111;
rom[60619] = 12'h111;
rom[60620] = 12'h111;
rom[60621] = 12'h  0;
rom[60622] = 12'h  0;
rom[60623] = 12'h  0;
rom[60624] = 12'h  0;
rom[60625] = 12'h  0;
rom[60626] = 12'h  0;
rom[60627] = 12'h  0;
rom[60628] = 12'h  0;
rom[60629] = 12'h  0;
rom[60630] = 12'h  0;
rom[60631] = 12'h  0;
rom[60632] = 12'h  0;
rom[60633] = 12'h  0;
rom[60634] = 12'h  0;
rom[60635] = 12'h  0;
rom[60636] = 12'h  0;
rom[60637] = 12'h  0;
rom[60638] = 12'h  0;
rom[60639] = 12'h  0;
rom[60640] = 12'h  0;
rom[60641] = 12'h  0;
rom[60642] = 12'h  0;
rom[60643] = 12'h  0;
rom[60644] = 12'h  0;
rom[60645] = 12'h  0;
rom[60646] = 12'h  0;
rom[60647] = 12'h  0;
rom[60648] = 12'h  0;
rom[60649] = 12'h  0;
rom[60650] = 12'h  0;
rom[60651] = 12'h  0;
rom[60652] = 12'h  0;
rom[60653] = 12'h  0;
rom[60654] = 12'h  0;
rom[60655] = 12'h  0;
rom[60656] = 12'h  0;
rom[60657] = 12'h  0;
rom[60658] = 12'h  0;
rom[60659] = 12'h  0;
rom[60660] = 12'h  0;
rom[60661] = 12'h  0;
rom[60662] = 12'h  0;
rom[60663] = 12'h  0;
rom[60664] = 12'h  0;
rom[60665] = 12'h  0;
rom[60666] = 12'h  0;
rom[60667] = 12'h  0;
rom[60668] = 12'h  0;
rom[60669] = 12'h  0;
rom[60670] = 12'h  0;
rom[60671] = 12'h  0;
rom[60672] = 12'h  0;
rom[60673] = 12'h111;
rom[60674] = 12'h111;
rom[60675] = 12'h222;
rom[60676] = 12'h222;
rom[60677] = 12'h333;
rom[60678] = 12'h333;
rom[60679] = 12'h333;
rom[60680] = 12'h444;
rom[60681] = 12'h444;
rom[60682] = 12'h555;
rom[60683] = 12'h444;
rom[60684] = 12'h333;
rom[60685] = 12'h222;
rom[60686] = 12'h222;
rom[60687] = 12'h222;
rom[60688] = 12'h222;
rom[60689] = 12'h222;
rom[60690] = 12'h222;
rom[60691] = 12'h222;
rom[60692] = 12'h222;
rom[60693] = 12'h222;
rom[60694] = 12'h333;
rom[60695] = 12'h333;
rom[60696] = 12'h333;
rom[60697] = 12'h444;
rom[60698] = 12'h555;
rom[60699] = 12'h555;
rom[60700] = 12'h555;
rom[60701] = 12'h444;
rom[60702] = 12'h444;
rom[60703] = 12'h555;
rom[60704] = 12'h555;
rom[60705] = 12'h555;
rom[60706] = 12'h555;
rom[60707] = 12'h555;
rom[60708] = 12'h666;
rom[60709] = 12'h666;
rom[60710] = 12'h666;
rom[60711] = 12'h666;
rom[60712] = 12'h555;
rom[60713] = 12'h555;
rom[60714] = 12'h555;
rom[60715] = 12'h555;
rom[60716] = 12'h555;
rom[60717] = 12'h555;
rom[60718] = 12'h666;
rom[60719] = 12'h666;
rom[60720] = 12'h666;
rom[60721] = 12'h666;
rom[60722] = 12'h666;
rom[60723] = 12'h666;
rom[60724] = 12'h777;
rom[60725] = 12'h777;
rom[60726] = 12'h777;
rom[60727] = 12'h777;
rom[60728] = 12'h777;
rom[60729] = 12'h777;
rom[60730] = 12'h777;
rom[60731] = 12'h777;
rom[60732] = 12'h888;
rom[60733] = 12'h888;
rom[60734] = 12'h888;
rom[60735] = 12'h888;
rom[60736] = 12'h888;
rom[60737] = 12'h888;
rom[60738] = 12'h999;
rom[60739] = 12'h999;
rom[60740] = 12'h999;
rom[60741] = 12'h999;
rom[60742] = 12'h999;
rom[60743] = 12'haaa;
rom[60744] = 12'haaa;
rom[60745] = 12'haaa;
rom[60746] = 12'hbbb;
rom[60747] = 12'hbbb;
rom[60748] = 12'hbbb;
rom[60749] = 12'hbbb;
rom[60750] = 12'hccc;
rom[60751] = 12'hccc;
rom[60752] = 12'hddd;
rom[60753] = 12'hddd;
rom[60754] = 12'heee;
rom[60755] = 12'heee;
rom[60756] = 12'hfff;
rom[60757] = 12'hfff;
rom[60758] = 12'heee;
rom[60759] = 12'heee;
rom[60760] = 12'hddd;
rom[60761] = 12'hddd;
rom[60762] = 12'hccc;
rom[60763] = 12'hccc;
rom[60764] = 12'hccc;
rom[60765] = 12'hbbb;
rom[60766] = 12'hbbb;
rom[60767] = 12'hbbb;
rom[60768] = 12'hbbb;
rom[60769] = 12'hbbb;
rom[60770] = 12'hbbb;
rom[60771] = 12'hbbb;
rom[60772] = 12'hbbb;
rom[60773] = 12'haaa;
rom[60774] = 12'haaa;
rom[60775] = 12'haaa;
rom[60776] = 12'h999;
rom[60777] = 12'h999;
rom[60778] = 12'h999;
rom[60779] = 12'h888;
rom[60780] = 12'h888;
rom[60781] = 12'h999;
rom[60782] = 12'h999;
rom[60783] = 12'h999;
rom[60784] = 12'h888;
rom[60785] = 12'h888;
rom[60786] = 12'h888;
rom[60787] = 12'h888;
rom[60788] = 12'h888;
rom[60789] = 12'h888;
rom[60790] = 12'h777;
rom[60791] = 12'h777;
rom[60792] = 12'h777;
rom[60793] = 12'h777;
rom[60794] = 12'h777;
rom[60795] = 12'h777;
rom[60796] = 12'h888;
rom[60797] = 12'h888;
rom[60798] = 12'h888;
rom[60799] = 12'h888;
rom[60800] = 12'hfff;
rom[60801] = 12'hfff;
rom[60802] = 12'hfff;
rom[60803] = 12'hfff;
rom[60804] = 12'hfff;
rom[60805] = 12'hfff;
rom[60806] = 12'hfff;
rom[60807] = 12'hfff;
rom[60808] = 12'hfff;
rom[60809] = 12'hfff;
rom[60810] = 12'hfff;
rom[60811] = 12'hfff;
rom[60812] = 12'hfff;
rom[60813] = 12'hfff;
rom[60814] = 12'hfff;
rom[60815] = 12'hfff;
rom[60816] = 12'hfff;
rom[60817] = 12'hfff;
rom[60818] = 12'hfff;
rom[60819] = 12'hfff;
rom[60820] = 12'hfff;
rom[60821] = 12'hfff;
rom[60822] = 12'hfff;
rom[60823] = 12'hfff;
rom[60824] = 12'hfff;
rom[60825] = 12'hfff;
rom[60826] = 12'hfff;
rom[60827] = 12'hfff;
rom[60828] = 12'hfff;
rom[60829] = 12'hfff;
rom[60830] = 12'hfff;
rom[60831] = 12'hfff;
rom[60832] = 12'hfff;
rom[60833] = 12'hfff;
rom[60834] = 12'hfff;
rom[60835] = 12'hfff;
rom[60836] = 12'hfff;
rom[60837] = 12'hfff;
rom[60838] = 12'hfff;
rom[60839] = 12'hfff;
rom[60840] = 12'hfff;
rom[60841] = 12'hfff;
rom[60842] = 12'hfff;
rom[60843] = 12'hfff;
rom[60844] = 12'hfff;
rom[60845] = 12'hfff;
rom[60846] = 12'hfff;
rom[60847] = 12'hfff;
rom[60848] = 12'hfff;
rom[60849] = 12'hfff;
rom[60850] = 12'hfff;
rom[60851] = 12'hfff;
rom[60852] = 12'hfff;
rom[60853] = 12'hfff;
rom[60854] = 12'hfff;
rom[60855] = 12'hfff;
rom[60856] = 12'hfff;
rom[60857] = 12'hfff;
rom[60858] = 12'hfff;
rom[60859] = 12'hfff;
rom[60860] = 12'hfff;
rom[60861] = 12'hfff;
rom[60862] = 12'hfff;
rom[60863] = 12'hfff;
rom[60864] = 12'hfff;
rom[60865] = 12'hfff;
rom[60866] = 12'hfff;
rom[60867] = 12'hfff;
rom[60868] = 12'hfff;
rom[60869] = 12'hfff;
rom[60870] = 12'hfff;
rom[60871] = 12'hfff;
rom[60872] = 12'hfff;
rom[60873] = 12'hfff;
rom[60874] = 12'hfff;
rom[60875] = 12'hfff;
rom[60876] = 12'hfff;
rom[60877] = 12'hfff;
rom[60878] = 12'hfff;
rom[60879] = 12'hfff;
rom[60880] = 12'hfff;
rom[60881] = 12'hfff;
rom[60882] = 12'hfff;
rom[60883] = 12'hfff;
rom[60884] = 12'hfff;
rom[60885] = 12'hfff;
rom[60886] = 12'hfff;
rom[60887] = 12'hfff;
rom[60888] = 12'hfff;
rom[60889] = 12'hfff;
rom[60890] = 12'hfff;
rom[60891] = 12'hfff;
rom[60892] = 12'hfff;
rom[60893] = 12'hfff;
rom[60894] = 12'hfff;
rom[60895] = 12'hfff;
rom[60896] = 12'hfff;
rom[60897] = 12'hfff;
rom[60898] = 12'hfff;
rom[60899] = 12'hfff;
rom[60900] = 12'heee;
rom[60901] = 12'heee;
rom[60902] = 12'hddd;
rom[60903] = 12'hddd;
rom[60904] = 12'hddd;
rom[60905] = 12'hddd;
rom[60906] = 12'hddd;
rom[60907] = 12'hddd;
rom[60908] = 12'hccc;
rom[60909] = 12'hccc;
rom[60910] = 12'hccc;
rom[60911] = 12'hccc;
rom[60912] = 12'hccc;
rom[60913] = 12'hccc;
rom[60914] = 12'hccc;
rom[60915] = 12'hccc;
rom[60916] = 12'hccc;
rom[60917] = 12'hbbb;
rom[60918] = 12'hbbb;
rom[60919] = 12'hbbb;
rom[60920] = 12'hbbb;
rom[60921] = 12'hbbb;
rom[60922] = 12'hbbb;
rom[60923] = 12'haaa;
rom[60924] = 12'haaa;
rom[60925] = 12'haaa;
rom[60926] = 12'haaa;
rom[60927] = 12'haaa;
rom[60928] = 12'haaa;
rom[60929] = 12'haaa;
rom[60930] = 12'haaa;
rom[60931] = 12'haaa;
rom[60932] = 12'haaa;
rom[60933] = 12'haaa;
rom[60934] = 12'h999;
rom[60935] = 12'h999;
rom[60936] = 12'h888;
rom[60937] = 12'h888;
rom[60938] = 12'h888;
rom[60939] = 12'h888;
rom[60940] = 12'h777;
rom[60941] = 12'h666;
rom[60942] = 12'h666;
rom[60943] = 12'h666;
rom[60944] = 12'h555;
rom[60945] = 12'h555;
rom[60946] = 12'h444;
rom[60947] = 12'h333;
rom[60948] = 12'h333;
rom[60949] = 12'h333;
rom[60950] = 12'h333;
rom[60951] = 12'h333;
rom[60952] = 12'h333;
rom[60953] = 12'h333;
rom[60954] = 12'h333;
rom[60955] = 12'h333;
rom[60956] = 12'h333;
rom[60957] = 12'h333;
rom[60958] = 12'h333;
rom[60959] = 12'h333;
rom[60960] = 12'h222;
rom[60961] = 12'h222;
rom[60962] = 12'h222;
rom[60963] = 12'h222;
rom[60964] = 12'h222;
rom[60965] = 12'h222;
rom[60966] = 12'h222;
rom[60967] = 12'h222;
rom[60968] = 12'h111;
rom[60969] = 12'h111;
rom[60970] = 12'h111;
rom[60971] = 12'h  0;
rom[60972] = 12'h  0;
rom[60973] = 12'h  0;
rom[60974] = 12'h  0;
rom[60975] = 12'h  0;
rom[60976] = 12'h  0;
rom[60977] = 12'h  0;
rom[60978] = 12'h  0;
rom[60979] = 12'h  0;
rom[60980] = 12'h  0;
rom[60981] = 12'h  0;
rom[60982] = 12'h  0;
rom[60983] = 12'h  0;
rom[60984] = 12'h  0;
rom[60985] = 12'h  0;
rom[60986] = 12'h  0;
rom[60987] = 12'h  0;
rom[60988] = 12'h  0;
rom[60989] = 12'h  0;
rom[60990] = 12'h  0;
rom[60991] = 12'h  0;
rom[60992] = 12'h  0;
rom[60993] = 12'h  0;
rom[60994] = 12'h  0;
rom[60995] = 12'h  0;
rom[60996] = 12'h  0;
rom[60997] = 12'h  0;
rom[60998] = 12'h  0;
rom[60999] = 12'h  0;
rom[61000] = 12'h  0;
rom[61001] = 12'h  0;
rom[61002] = 12'h111;
rom[61003] = 12'h111;
rom[61004] = 12'h111;
rom[61005] = 12'h111;
rom[61006] = 12'h111;
rom[61007] = 12'h111;
rom[61008] = 12'h111;
rom[61009] = 12'h111;
rom[61010] = 12'h111;
rom[61011] = 12'h111;
rom[61012] = 12'h111;
rom[61013] = 12'h222;
rom[61014] = 12'h222;
rom[61015] = 12'h222;
rom[61016] = 12'h111;
rom[61017] = 12'h111;
rom[61018] = 12'h111;
rom[61019] = 12'h111;
rom[61020] = 12'h111;
rom[61021] = 12'h111;
rom[61022] = 12'h111;
rom[61023] = 12'h  0;
rom[61024] = 12'h  0;
rom[61025] = 12'h  0;
rom[61026] = 12'h  0;
rom[61027] = 12'h  0;
rom[61028] = 12'h  0;
rom[61029] = 12'h  0;
rom[61030] = 12'h  0;
rom[61031] = 12'h  0;
rom[61032] = 12'h  0;
rom[61033] = 12'h  0;
rom[61034] = 12'h  0;
rom[61035] = 12'h  0;
rom[61036] = 12'h  0;
rom[61037] = 12'h  0;
rom[61038] = 12'h  0;
rom[61039] = 12'h  0;
rom[61040] = 12'h  0;
rom[61041] = 12'h  0;
rom[61042] = 12'h  0;
rom[61043] = 12'h  0;
rom[61044] = 12'h  0;
rom[61045] = 12'h  0;
rom[61046] = 12'h  0;
rom[61047] = 12'h  0;
rom[61048] = 12'h  0;
rom[61049] = 12'h  0;
rom[61050] = 12'h  0;
rom[61051] = 12'h  0;
rom[61052] = 12'h  0;
rom[61053] = 12'h  0;
rom[61054] = 12'h  0;
rom[61055] = 12'h  0;
rom[61056] = 12'h  0;
rom[61057] = 12'h  0;
rom[61058] = 12'h  0;
rom[61059] = 12'h  0;
rom[61060] = 12'h  0;
rom[61061] = 12'h  0;
rom[61062] = 12'h  0;
rom[61063] = 12'h  0;
rom[61064] = 12'h  0;
rom[61065] = 12'h  0;
rom[61066] = 12'h  0;
rom[61067] = 12'h  0;
rom[61068] = 12'h  0;
rom[61069] = 12'h  0;
rom[61070] = 12'h  0;
rom[61071] = 12'h  0;
rom[61072] = 12'h  0;
rom[61073] = 12'h111;
rom[61074] = 12'h111;
rom[61075] = 12'h222;
rom[61076] = 12'h222;
rom[61077] = 12'h333;
rom[61078] = 12'h333;
rom[61079] = 12'h444;
rom[61080] = 12'h444;
rom[61081] = 12'h555;
rom[61082] = 12'h555;
rom[61083] = 12'h444;
rom[61084] = 12'h333;
rom[61085] = 12'h222;
rom[61086] = 12'h222;
rom[61087] = 12'h222;
rom[61088] = 12'h222;
rom[61089] = 12'h222;
rom[61090] = 12'h222;
rom[61091] = 12'h222;
rom[61092] = 12'h222;
rom[61093] = 12'h222;
rom[61094] = 12'h222;
rom[61095] = 12'h222;
rom[61096] = 12'h333;
rom[61097] = 12'h444;
rom[61098] = 12'h555;
rom[61099] = 12'h555;
rom[61100] = 12'h444;
rom[61101] = 12'h444;
rom[61102] = 12'h444;
rom[61103] = 12'h444;
rom[61104] = 12'h555;
rom[61105] = 12'h555;
rom[61106] = 12'h555;
rom[61107] = 12'h555;
rom[61108] = 12'h666;
rom[61109] = 12'h666;
rom[61110] = 12'h666;
rom[61111] = 12'h666;
rom[61112] = 12'h666;
rom[61113] = 12'h666;
rom[61114] = 12'h555;
rom[61115] = 12'h555;
rom[61116] = 12'h555;
rom[61117] = 12'h666;
rom[61118] = 12'h666;
rom[61119] = 12'h666;
rom[61120] = 12'h666;
rom[61121] = 12'h666;
rom[61122] = 12'h666;
rom[61123] = 12'h666;
rom[61124] = 12'h777;
rom[61125] = 12'h777;
rom[61126] = 12'h777;
rom[61127] = 12'h777;
rom[61128] = 12'h777;
rom[61129] = 12'h777;
rom[61130] = 12'h777;
rom[61131] = 12'h888;
rom[61132] = 12'h888;
rom[61133] = 12'h888;
rom[61134] = 12'h888;
rom[61135] = 12'h999;
rom[61136] = 12'h999;
rom[61137] = 12'h999;
rom[61138] = 12'h999;
rom[61139] = 12'h999;
rom[61140] = 12'h999;
rom[61141] = 12'h999;
rom[61142] = 12'haaa;
rom[61143] = 12'haaa;
rom[61144] = 12'haaa;
rom[61145] = 12'haaa;
rom[61146] = 12'hbbb;
rom[61147] = 12'hbbb;
rom[61148] = 12'hbbb;
rom[61149] = 12'hccc;
rom[61150] = 12'hccc;
rom[61151] = 12'hccc;
rom[61152] = 12'hddd;
rom[61153] = 12'heee;
rom[61154] = 12'hfff;
rom[61155] = 12'hfff;
rom[61156] = 12'hfff;
rom[61157] = 12'hfff;
rom[61158] = 12'heee;
rom[61159] = 12'hddd;
rom[61160] = 12'hddd;
rom[61161] = 12'hddd;
rom[61162] = 12'hccc;
rom[61163] = 12'hccc;
rom[61164] = 12'hccc;
rom[61165] = 12'hccc;
rom[61166] = 12'hbbb;
rom[61167] = 12'hbbb;
rom[61168] = 12'hbbb;
rom[61169] = 12'hbbb;
rom[61170] = 12'hbbb;
rom[61171] = 12'hbbb;
rom[61172] = 12'hbbb;
rom[61173] = 12'hbbb;
rom[61174] = 12'haaa;
rom[61175] = 12'haaa;
rom[61176] = 12'h999;
rom[61177] = 12'h999;
rom[61178] = 12'h999;
rom[61179] = 12'h888;
rom[61180] = 12'h888;
rom[61181] = 12'h888;
rom[61182] = 12'h888;
rom[61183] = 12'h888;
rom[61184] = 12'h888;
rom[61185] = 12'h888;
rom[61186] = 12'h888;
rom[61187] = 12'h777;
rom[61188] = 12'h777;
rom[61189] = 12'h777;
rom[61190] = 12'h777;
rom[61191] = 12'h777;
rom[61192] = 12'h777;
rom[61193] = 12'h777;
rom[61194] = 12'h777;
rom[61195] = 12'h777;
rom[61196] = 12'h777;
rom[61197] = 12'h777;
rom[61198] = 12'h777;
rom[61199] = 12'h777;
rom[61200] = 12'hfff;
rom[61201] = 12'hfff;
rom[61202] = 12'hfff;
rom[61203] = 12'hfff;
rom[61204] = 12'hfff;
rom[61205] = 12'hfff;
rom[61206] = 12'hfff;
rom[61207] = 12'hfff;
rom[61208] = 12'hfff;
rom[61209] = 12'hfff;
rom[61210] = 12'hfff;
rom[61211] = 12'hfff;
rom[61212] = 12'hfff;
rom[61213] = 12'hfff;
rom[61214] = 12'hfff;
rom[61215] = 12'hfff;
rom[61216] = 12'hfff;
rom[61217] = 12'hfff;
rom[61218] = 12'hfff;
rom[61219] = 12'hfff;
rom[61220] = 12'hfff;
rom[61221] = 12'hfff;
rom[61222] = 12'hfff;
rom[61223] = 12'hfff;
rom[61224] = 12'hfff;
rom[61225] = 12'hfff;
rom[61226] = 12'hfff;
rom[61227] = 12'hfff;
rom[61228] = 12'hfff;
rom[61229] = 12'hfff;
rom[61230] = 12'hfff;
rom[61231] = 12'hfff;
rom[61232] = 12'hfff;
rom[61233] = 12'hfff;
rom[61234] = 12'hfff;
rom[61235] = 12'hfff;
rom[61236] = 12'hfff;
rom[61237] = 12'hfff;
rom[61238] = 12'hfff;
rom[61239] = 12'hfff;
rom[61240] = 12'hfff;
rom[61241] = 12'hfff;
rom[61242] = 12'hfff;
rom[61243] = 12'hfff;
rom[61244] = 12'hfff;
rom[61245] = 12'hfff;
rom[61246] = 12'hfff;
rom[61247] = 12'hfff;
rom[61248] = 12'hfff;
rom[61249] = 12'hfff;
rom[61250] = 12'hfff;
rom[61251] = 12'hfff;
rom[61252] = 12'hfff;
rom[61253] = 12'hfff;
rom[61254] = 12'hfff;
rom[61255] = 12'hfff;
rom[61256] = 12'hfff;
rom[61257] = 12'hfff;
rom[61258] = 12'hfff;
rom[61259] = 12'hfff;
rom[61260] = 12'hfff;
rom[61261] = 12'hfff;
rom[61262] = 12'hfff;
rom[61263] = 12'hfff;
rom[61264] = 12'hfff;
rom[61265] = 12'hfff;
rom[61266] = 12'hfff;
rom[61267] = 12'hfff;
rom[61268] = 12'hfff;
rom[61269] = 12'hfff;
rom[61270] = 12'hfff;
rom[61271] = 12'hfff;
rom[61272] = 12'hfff;
rom[61273] = 12'hfff;
rom[61274] = 12'hfff;
rom[61275] = 12'hfff;
rom[61276] = 12'hfff;
rom[61277] = 12'hfff;
rom[61278] = 12'hfff;
rom[61279] = 12'hfff;
rom[61280] = 12'hfff;
rom[61281] = 12'hfff;
rom[61282] = 12'hfff;
rom[61283] = 12'hfff;
rom[61284] = 12'hfff;
rom[61285] = 12'hfff;
rom[61286] = 12'hfff;
rom[61287] = 12'hfff;
rom[61288] = 12'hfff;
rom[61289] = 12'hfff;
rom[61290] = 12'hfff;
rom[61291] = 12'hfff;
rom[61292] = 12'hfff;
rom[61293] = 12'hfff;
rom[61294] = 12'hfff;
rom[61295] = 12'hfff;
rom[61296] = 12'hfff;
rom[61297] = 12'hfff;
rom[61298] = 12'hfff;
rom[61299] = 12'hfff;
rom[61300] = 12'hfff;
rom[61301] = 12'heee;
rom[61302] = 12'heee;
rom[61303] = 12'heee;
rom[61304] = 12'hddd;
rom[61305] = 12'hddd;
rom[61306] = 12'hddd;
rom[61307] = 12'hddd;
rom[61308] = 12'hddd;
rom[61309] = 12'hccc;
rom[61310] = 12'hccc;
rom[61311] = 12'hccc;
rom[61312] = 12'hccc;
rom[61313] = 12'hccc;
rom[61314] = 12'hccc;
rom[61315] = 12'hccc;
rom[61316] = 12'hccc;
rom[61317] = 12'hccc;
rom[61318] = 12'hccc;
rom[61319] = 12'hccc;
rom[61320] = 12'hbbb;
rom[61321] = 12'hbbb;
rom[61322] = 12'hbbb;
rom[61323] = 12'haaa;
rom[61324] = 12'haaa;
rom[61325] = 12'haaa;
rom[61326] = 12'haaa;
rom[61327] = 12'haaa;
rom[61328] = 12'haaa;
rom[61329] = 12'h999;
rom[61330] = 12'h999;
rom[61331] = 12'h999;
rom[61332] = 12'h999;
rom[61333] = 12'h999;
rom[61334] = 12'h999;
rom[61335] = 12'h999;
rom[61336] = 12'h999;
rom[61337] = 12'h999;
rom[61338] = 12'h999;
rom[61339] = 12'h888;
rom[61340] = 12'h888;
rom[61341] = 12'h777;
rom[61342] = 12'h777;
rom[61343] = 12'h666;
rom[61344] = 12'h666;
rom[61345] = 12'h666;
rom[61346] = 12'h555;
rom[61347] = 12'h444;
rom[61348] = 12'h444;
rom[61349] = 12'h444;
rom[61350] = 12'h444;
rom[61351] = 12'h444;
rom[61352] = 12'h444;
rom[61353] = 12'h444;
rom[61354] = 12'h333;
rom[61355] = 12'h333;
rom[61356] = 12'h333;
rom[61357] = 12'h333;
rom[61358] = 12'h222;
rom[61359] = 12'h222;
rom[61360] = 12'h222;
rom[61361] = 12'h222;
rom[61362] = 12'h333;
rom[61363] = 12'h333;
rom[61364] = 12'h222;
rom[61365] = 12'h222;
rom[61366] = 12'h222;
rom[61367] = 12'h222;
rom[61368] = 12'h111;
rom[61369] = 12'h111;
rom[61370] = 12'h111;
rom[61371] = 12'h  0;
rom[61372] = 12'h111;
rom[61373] = 12'h111;
rom[61374] = 12'h  0;
rom[61375] = 12'h  0;
rom[61376] = 12'h  0;
rom[61377] = 12'h  0;
rom[61378] = 12'h  0;
rom[61379] = 12'h  0;
rom[61380] = 12'h  0;
rom[61381] = 12'h  0;
rom[61382] = 12'h  0;
rom[61383] = 12'h  0;
rom[61384] = 12'h  0;
rom[61385] = 12'h  0;
rom[61386] = 12'h  0;
rom[61387] = 12'h  0;
rom[61388] = 12'h  0;
rom[61389] = 12'h  0;
rom[61390] = 12'h  0;
rom[61391] = 12'h  0;
rom[61392] = 12'h  0;
rom[61393] = 12'h  0;
rom[61394] = 12'h  0;
rom[61395] = 12'h  0;
rom[61396] = 12'h  0;
rom[61397] = 12'h  0;
rom[61398] = 12'h  0;
rom[61399] = 12'h  0;
rom[61400] = 12'h  0;
rom[61401] = 12'h  0;
rom[61402] = 12'h111;
rom[61403] = 12'h111;
rom[61404] = 12'h111;
rom[61405] = 12'h111;
rom[61406] = 12'h111;
rom[61407] = 12'h  0;
rom[61408] = 12'h  0;
rom[61409] = 12'h111;
rom[61410] = 12'h111;
rom[61411] = 12'h111;
rom[61412] = 12'h111;
rom[61413] = 12'h222;
rom[61414] = 12'h222;
rom[61415] = 12'h222;
rom[61416] = 12'h111;
rom[61417] = 12'h111;
rom[61418] = 12'h111;
rom[61419] = 12'h111;
rom[61420] = 12'h111;
rom[61421] = 12'h111;
rom[61422] = 12'h111;
rom[61423] = 12'h  0;
rom[61424] = 12'h  0;
rom[61425] = 12'h  0;
rom[61426] = 12'h  0;
rom[61427] = 12'h  0;
rom[61428] = 12'h  0;
rom[61429] = 12'h  0;
rom[61430] = 12'h  0;
rom[61431] = 12'h  0;
rom[61432] = 12'h  0;
rom[61433] = 12'h  0;
rom[61434] = 12'h  0;
rom[61435] = 12'h  0;
rom[61436] = 12'h  0;
rom[61437] = 12'h  0;
rom[61438] = 12'h  0;
rom[61439] = 12'h  0;
rom[61440] = 12'h  0;
rom[61441] = 12'h  0;
rom[61442] = 12'h  0;
rom[61443] = 12'h  0;
rom[61444] = 12'h  0;
rom[61445] = 12'h  0;
rom[61446] = 12'h  0;
rom[61447] = 12'h  0;
rom[61448] = 12'h  0;
rom[61449] = 12'h  0;
rom[61450] = 12'h  0;
rom[61451] = 12'h  0;
rom[61452] = 12'h  0;
rom[61453] = 12'h  0;
rom[61454] = 12'h  0;
rom[61455] = 12'h  0;
rom[61456] = 12'h  0;
rom[61457] = 12'h  0;
rom[61458] = 12'h  0;
rom[61459] = 12'h  0;
rom[61460] = 12'h  0;
rom[61461] = 12'h  0;
rom[61462] = 12'h  0;
rom[61463] = 12'h  0;
rom[61464] = 12'h  0;
rom[61465] = 12'h  0;
rom[61466] = 12'h  0;
rom[61467] = 12'h  0;
rom[61468] = 12'h  0;
rom[61469] = 12'h  0;
rom[61470] = 12'h  0;
rom[61471] = 12'h  0;
rom[61472] = 12'h  0;
rom[61473] = 12'h111;
rom[61474] = 12'h111;
rom[61475] = 12'h222;
rom[61476] = 12'h222;
rom[61477] = 12'h333;
rom[61478] = 12'h333;
rom[61479] = 12'h444;
rom[61480] = 12'h444;
rom[61481] = 12'h555;
rom[61482] = 12'h555;
rom[61483] = 12'h444;
rom[61484] = 12'h333;
rom[61485] = 12'h222;
rom[61486] = 12'h222;
rom[61487] = 12'h222;
rom[61488] = 12'h222;
rom[61489] = 12'h222;
rom[61490] = 12'h222;
rom[61491] = 12'h222;
rom[61492] = 12'h222;
rom[61493] = 12'h222;
rom[61494] = 12'h222;
rom[61495] = 12'h222;
rom[61496] = 12'h333;
rom[61497] = 12'h444;
rom[61498] = 12'h555;
rom[61499] = 12'h555;
rom[61500] = 12'h555;
rom[61501] = 12'h444;
rom[61502] = 12'h444;
rom[61503] = 12'h444;
rom[61504] = 12'h444;
rom[61505] = 12'h444;
rom[61506] = 12'h555;
rom[61507] = 12'h555;
rom[61508] = 12'h666;
rom[61509] = 12'h666;
rom[61510] = 12'h666;
rom[61511] = 12'h666;
rom[61512] = 12'h666;
rom[61513] = 12'h666;
rom[61514] = 12'h666;
rom[61515] = 12'h666;
rom[61516] = 12'h666;
rom[61517] = 12'h666;
rom[61518] = 12'h666;
rom[61519] = 12'h666;
rom[61520] = 12'h666;
rom[61521] = 12'h666;
rom[61522] = 12'h666;
rom[61523] = 12'h666;
rom[61524] = 12'h777;
rom[61525] = 12'h777;
rom[61526] = 12'h777;
rom[61527] = 12'h777;
rom[61528] = 12'h777;
rom[61529] = 12'h777;
rom[61530] = 12'h888;
rom[61531] = 12'h888;
rom[61532] = 12'h888;
rom[61533] = 12'h888;
rom[61534] = 12'h999;
rom[61535] = 12'h999;
rom[61536] = 12'h999;
rom[61537] = 12'h999;
rom[61538] = 12'h999;
rom[61539] = 12'h999;
rom[61540] = 12'haaa;
rom[61541] = 12'haaa;
rom[61542] = 12'haaa;
rom[61543] = 12'haaa;
rom[61544] = 12'haaa;
rom[61545] = 12'hbbb;
rom[61546] = 12'hbbb;
rom[61547] = 12'hbbb;
rom[61548] = 12'hccc;
rom[61549] = 12'hccc;
rom[61550] = 12'hccc;
rom[61551] = 12'hddd;
rom[61552] = 12'heee;
rom[61553] = 12'heee;
rom[61554] = 12'hfff;
rom[61555] = 12'hfff;
rom[61556] = 12'hfff;
rom[61557] = 12'heee;
rom[61558] = 12'heee;
rom[61559] = 12'hddd;
rom[61560] = 12'hddd;
rom[61561] = 12'hddd;
rom[61562] = 12'hccc;
rom[61563] = 12'hccc;
rom[61564] = 12'hccc;
rom[61565] = 12'hccc;
rom[61566] = 12'hbbb;
rom[61567] = 12'hbbb;
rom[61568] = 12'hbbb;
rom[61569] = 12'hbbb;
rom[61570] = 12'hbbb;
rom[61571] = 12'hbbb;
rom[61572] = 12'hbbb;
rom[61573] = 12'hbbb;
rom[61574] = 12'haaa;
rom[61575] = 12'haaa;
rom[61576] = 12'h999;
rom[61577] = 12'h999;
rom[61578] = 12'h999;
rom[61579] = 12'h888;
rom[61580] = 12'h888;
rom[61581] = 12'h888;
rom[61582] = 12'h888;
rom[61583] = 12'h888;
rom[61584] = 12'h888;
rom[61585] = 12'h777;
rom[61586] = 12'h777;
rom[61587] = 12'h777;
rom[61588] = 12'h777;
rom[61589] = 12'h777;
rom[61590] = 12'h777;
rom[61591] = 12'h777;
rom[61592] = 12'h777;
rom[61593] = 12'h777;
rom[61594] = 12'h777;
rom[61595] = 12'h777;
rom[61596] = 12'h777;
rom[61597] = 12'h777;
rom[61598] = 12'h777;
rom[61599] = 12'h777;
rom[61600] = 12'hfff;
rom[61601] = 12'hfff;
rom[61602] = 12'hfff;
rom[61603] = 12'hfff;
rom[61604] = 12'hfff;
rom[61605] = 12'hfff;
rom[61606] = 12'hfff;
rom[61607] = 12'hfff;
rom[61608] = 12'hfff;
rom[61609] = 12'hfff;
rom[61610] = 12'hfff;
rom[61611] = 12'hfff;
rom[61612] = 12'hfff;
rom[61613] = 12'hfff;
rom[61614] = 12'hfff;
rom[61615] = 12'hfff;
rom[61616] = 12'hfff;
rom[61617] = 12'hfff;
rom[61618] = 12'hfff;
rom[61619] = 12'hfff;
rom[61620] = 12'hfff;
rom[61621] = 12'hfff;
rom[61622] = 12'hfff;
rom[61623] = 12'hfff;
rom[61624] = 12'hfff;
rom[61625] = 12'hfff;
rom[61626] = 12'hfff;
rom[61627] = 12'hfff;
rom[61628] = 12'hfff;
rom[61629] = 12'hfff;
rom[61630] = 12'hfff;
rom[61631] = 12'hfff;
rom[61632] = 12'hfff;
rom[61633] = 12'hfff;
rom[61634] = 12'hfff;
rom[61635] = 12'hfff;
rom[61636] = 12'hfff;
rom[61637] = 12'hfff;
rom[61638] = 12'hfff;
rom[61639] = 12'hfff;
rom[61640] = 12'hfff;
rom[61641] = 12'hfff;
rom[61642] = 12'hfff;
rom[61643] = 12'hfff;
rom[61644] = 12'hfff;
rom[61645] = 12'hfff;
rom[61646] = 12'hfff;
rom[61647] = 12'hfff;
rom[61648] = 12'hfff;
rom[61649] = 12'hfff;
rom[61650] = 12'hfff;
rom[61651] = 12'hfff;
rom[61652] = 12'hfff;
rom[61653] = 12'hfff;
rom[61654] = 12'hfff;
rom[61655] = 12'hfff;
rom[61656] = 12'hfff;
rom[61657] = 12'hfff;
rom[61658] = 12'hfff;
rom[61659] = 12'hfff;
rom[61660] = 12'hfff;
rom[61661] = 12'hfff;
rom[61662] = 12'hfff;
rom[61663] = 12'hfff;
rom[61664] = 12'hfff;
rom[61665] = 12'hfff;
rom[61666] = 12'hfff;
rom[61667] = 12'hfff;
rom[61668] = 12'hfff;
rom[61669] = 12'hfff;
rom[61670] = 12'hfff;
rom[61671] = 12'hfff;
rom[61672] = 12'hfff;
rom[61673] = 12'hfff;
rom[61674] = 12'hfff;
rom[61675] = 12'hfff;
rom[61676] = 12'hfff;
rom[61677] = 12'hfff;
rom[61678] = 12'hfff;
rom[61679] = 12'hfff;
rom[61680] = 12'hfff;
rom[61681] = 12'hfff;
rom[61682] = 12'hfff;
rom[61683] = 12'hfff;
rom[61684] = 12'hfff;
rom[61685] = 12'hfff;
rom[61686] = 12'hfff;
rom[61687] = 12'hfff;
rom[61688] = 12'hfff;
rom[61689] = 12'hfff;
rom[61690] = 12'hfff;
rom[61691] = 12'hfff;
rom[61692] = 12'hfff;
rom[61693] = 12'hfff;
rom[61694] = 12'hfff;
rom[61695] = 12'hfff;
rom[61696] = 12'hfff;
rom[61697] = 12'hfff;
rom[61698] = 12'hfff;
rom[61699] = 12'hfff;
rom[61700] = 12'hfff;
rom[61701] = 12'hfff;
rom[61702] = 12'hfff;
rom[61703] = 12'heee;
rom[61704] = 12'heee;
rom[61705] = 12'heee;
rom[61706] = 12'heee;
rom[61707] = 12'hddd;
rom[61708] = 12'hddd;
rom[61709] = 12'hddd;
rom[61710] = 12'hddd;
rom[61711] = 12'hddd;
rom[61712] = 12'hccc;
rom[61713] = 12'hccc;
rom[61714] = 12'hccc;
rom[61715] = 12'hccc;
rom[61716] = 12'hccc;
rom[61717] = 12'hccc;
rom[61718] = 12'hccc;
rom[61719] = 12'hccc;
rom[61720] = 12'hbbb;
rom[61721] = 12'hbbb;
rom[61722] = 12'hbbb;
rom[61723] = 12'hbbb;
rom[61724] = 12'haaa;
rom[61725] = 12'haaa;
rom[61726] = 12'haaa;
rom[61727] = 12'h999;
rom[61728] = 12'h999;
rom[61729] = 12'h999;
rom[61730] = 12'h888;
rom[61731] = 12'h888;
rom[61732] = 12'h888;
rom[61733] = 12'h999;
rom[61734] = 12'h999;
rom[61735] = 12'h999;
rom[61736] = 12'h999;
rom[61737] = 12'h999;
rom[61738] = 12'h999;
rom[61739] = 12'h999;
rom[61740] = 12'h888;
rom[61741] = 12'h888;
rom[61742] = 12'h888;
rom[61743] = 12'h777;
rom[61744] = 12'h777;
rom[61745] = 12'h777;
rom[61746] = 12'h666;
rom[61747] = 12'h666;
rom[61748] = 12'h555;
rom[61749] = 12'h555;
rom[61750] = 12'h444;
rom[61751] = 12'h444;
rom[61752] = 12'h444;
rom[61753] = 12'h444;
rom[61754] = 12'h444;
rom[61755] = 12'h333;
rom[61756] = 12'h333;
rom[61757] = 12'h333;
rom[61758] = 12'h333;
rom[61759] = 12'h222;
rom[61760] = 12'h333;
rom[61761] = 12'h333;
rom[61762] = 12'h333;
rom[61763] = 12'h333;
rom[61764] = 12'h222;
rom[61765] = 12'h222;
rom[61766] = 12'h222;
rom[61767] = 12'h222;
rom[61768] = 12'h111;
rom[61769] = 12'h111;
rom[61770] = 12'h111;
rom[61771] = 12'h111;
rom[61772] = 12'h111;
rom[61773] = 12'h111;
rom[61774] = 12'h111;
rom[61775] = 12'h111;
rom[61776] = 12'h  0;
rom[61777] = 12'h  0;
rom[61778] = 12'h  0;
rom[61779] = 12'h  0;
rom[61780] = 12'h  0;
rom[61781] = 12'h  0;
rom[61782] = 12'h  0;
rom[61783] = 12'h  0;
rom[61784] = 12'h  0;
rom[61785] = 12'h  0;
rom[61786] = 12'h  0;
rom[61787] = 12'h  0;
rom[61788] = 12'h  0;
rom[61789] = 12'h  0;
rom[61790] = 12'h  0;
rom[61791] = 12'h  0;
rom[61792] = 12'h  0;
rom[61793] = 12'h  0;
rom[61794] = 12'h  0;
rom[61795] = 12'h  0;
rom[61796] = 12'h  0;
rom[61797] = 12'h  0;
rom[61798] = 12'h  0;
rom[61799] = 12'h  0;
rom[61800] = 12'h  0;
rom[61801] = 12'h  0;
rom[61802] = 12'h  0;
rom[61803] = 12'h  0;
rom[61804] = 12'h  0;
rom[61805] = 12'h  0;
rom[61806] = 12'h  0;
rom[61807] = 12'h  0;
rom[61808] = 12'h  0;
rom[61809] = 12'h111;
rom[61810] = 12'h111;
rom[61811] = 12'h111;
rom[61812] = 12'h222;
rom[61813] = 12'h222;
rom[61814] = 12'h222;
rom[61815] = 12'h222;
rom[61816] = 12'h111;
rom[61817] = 12'h111;
rom[61818] = 12'h111;
rom[61819] = 12'h111;
rom[61820] = 12'h111;
rom[61821] = 12'h111;
rom[61822] = 12'h111;
rom[61823] = 12'h  0;
rom[61824] = 12'h  0;
rom[61825] = 12'h  0;
rom[61826] = 12'h  0;
rom[61827] = 12'h  0;
rom[61828] = 12'h  0;
rom[61829] = 12'h  0;
rom[61830] = 12'h  0;
rom[61831] = 12'h  0;
rom[61832] = 12'h  0;
rom[61833] = 12'h  0;
rom[61834] = 12'h  0;
rom[61835] = 12'h  0;
rom[61836] = 12'h  0;
rom[61837] = 12'h  0;
rom[61838] = 12'h  0;
rom[61839] = 12'h  0;
rom[61840] = 12'h  0;
rom[61841] = 12'h  0;
rom[61842] = 12'h  0;
rom[61843] = 12'h  0;
rom[61844] = 12'h  0;
rom[61845] = 12'h  0;
rom[61846] = 12'h  0;
rom[61847] = 12'h  0;
rom[61848] = 12'h  0;
rom[61849] = 12'h  0;
rom[61850] = 12'h  0;
rom[61851] = 12'h  0;
rom[61852] = 12'h  0;
rom[61853] = 12'h  0;
rom[61854] = 12'h  0;
rom[61855] = 12'h  0;
rom[61856] = 12'h  0;
rom[61857] = 12'h  0;
rom[61858] = 12'h  0;
rom[61859] = 12'h  0;
rom[61860] = 12'h  0;
rom[61861] = 12'h  0;
rom[61862] = 12'h  0;
rom[61863] = 12'h  0;
rom[61864] = 12'h  0;
rom[61865] = 12'h  0;
rom[61866] = 12'h  0;
rom[61867] = 12'h  0;
rom[61868] = 12'h  0;
rom[61869] = 12'h  0;
rom[61870] = 12'h  0;
rom[61871] = 12'h  0;
rom[61872] = 12'h  0;
rom[61873] = 12'h111;
rom[61874] = 12'h111;
rom[61875] = 12'h222;
rom[61876] = 12'h222;
rom[61877] = 12'h333;
rom[61878] = 12'h444;
rom[61879] = 12'h444;
rom[61880] = 12'h444;
rom[61881] = 12'h555;
rom[61882] = 12'h555;
rom[61883] = 12'h444;
rom[61884] = 12'h333;
rom[61885] = 12'h222;
rom[61886] = 12'h222;
rom[61887] = 12'h222;
rom[61888] = 12'h222;
rom[61889] = 12'h222;
rom[61890] = 12'h222;
rom[61891] = 12'h222;
rom[61892] = 12'h222;
rom[61893] = 12'h222;
rom[61894] = 12'h222;
rom[61895] = 12'h222;
rom[61896] = 12'h222;
rom[61897] = 12'h444;
rom[61898] = 12'h555;
rom[61899] = 12'h555;
rom[61900] = 12'h555;
rom[61901] = 12'h444;
rom[61902] = 12'h444;
rom[61903] = 12'h444;
rom[61904] = 12'h444;
rom[61905] = 12'h444;
rom[61906] = 12'h444;
rom[61907] = 12'h555;
rom[61908] = 12'h555;
rom[61909] = 12'h666;
rom[61910] = 12'h666;
rom[61911] = 12'h777;
rom[61912] = 12'h777;
rom[61913] = 12'h666;
rom[61914] = 12'h666;
rom[61915] = 12'h666;
rom[61916] = 12'h666;
rom[61917] = 12'h666;
rom[61918] = 12'h666;
rom[61919] = 12'h666;
rom[61920] = 12'h666;
rom[61921] = 12'h666;
rom[61922] = 12'h666;
rom[61923] = 12'h666;
rom[61924] = 12'h777;
rom[61925] = 12'h777;
rom[61926] = 12'h777;
rom[61927] = 12'h777;
rom[61928] = 12'h888;
rom[61929] = 12'h888;
rom[61930] = 12'h888;
rom[61931] = 12'h888;
rom[61932] = 12'h888;
rom[61933] = 12'h999;
rom[61934] = 12'h999;
rom[61935] = 12'h999;
rom[61936] = 12'h999;
rom[61937] = 12'h999;
rom[61938] = 12'h999;
rom[61939] = 12'haaa;
rom[61940] = 12'haaa;
rom[61941] = 12'haaa;
rom[61942] = 12'haaa;
rom[61943] = 12'haaa;
rom[61944] = 12'hbbb;
rom[61945] = 12'hbbb;
rom[61946] = 12'hbbb;
rom[61947] = 12'hccc;
rom[61948] = 12'hccc;
rom[61949] = 12'hccc;
rom[61950] = 12'hddd;
rom[61951] = 12'hddd;
rom[61952] = 12'heee;
rom[61953] = 12'hfff;
rom[61954] = 12'hfff;
rom[61955] = 12'hfff;
rom[61956] = 12'hfff;
rom[61957] = 12'heee;
rom[61958] = 12'hddd;
rom[61959] = 12'hddd;
rom[61960] = 12'hccc;
rom[61961] = 12'hccc;
rom[61962] = 12'hccc;
rom[61963] = 12'hccc;
rom[61964] = 12'hbbb;
rom[61965] = 12'hbbb;
rom[61966] = 12'hbbb;
rom[61967] = 12'hbbb;
rom[61968] = 12'hbbb;
rom[61969] = 12'hbbb;
rom[61970] = 12'hbbb;
rom[61971] = 12'hbbb;
rom[61972] = 12'hbbb;
rom[61973] = 12'hbbb;
rom[61974] = 12'hbbb;
rom[61975] = 12'haaa;
rom[61976] = 12'h999;
rom[61977] = 12'h999;
rom[61978] = 12'h999;
rom[61979] = 12'h888;
rom[61980] = 12'h888;
rom[61981] = 12'h888;
rom[61982] = 12'h888;
rom[61983] = 12'h888;
rom[61984] = 12'h777;
rom[61985] = 12'h777;
rom[61986] = 12'h777;
rom[61987] = 12'h777;
rom[61988] = 12'h777;
rom[61989] = 12'h777;
rom[61990] = 12'h777;
rom[61991] = 12'h777;
rom[61992] = 12'h777;
rom[61993] = 12'h777;
rom[61994] = 12'h777;
rom[61995] = 12'h777;
rom[61996] = 12'h777;
rom[61997] = 12'h777;
rom[61998] = 12'h777;
rom[61999] = 12'h777;
rom[62000] = 12'hfff;
rom[62001] = 12'hfff;
rom[62002] = 12'hfff;
rom[62003] = 12'hfff;
rom[62004] = 12'hfff;
rom[62005] = 12'hfff;
rom[62006] = 12'hfff;
rom[62007] = 12'hfff;
rom[62008] = 12'hfff;
rom[62009] = 12'hfff;
rom[62010] = 12'hfff;
rom[62011] = 12'hfff;
rom[62012] = 12'hfff;
rom[62013] = 12'hfff;
rom[62014] = 12'hfff;
rom[62015] = 12'hfff;
rom[62016] = 12'hfff;
rom[62017] = 12'hfff;
rom[62018] = 12'hfff;
rom[62019] = 12'hfff;
rom[62020] = 12'hfff;
rom[62021] = 12'hfff;
rom[62022] = 12'hfff;
rom[62023] = 12'hfff;
rom[62024] = 12'hfff;
rom[62025] = 12'hfff;
rom[62026] = 12'hfff;
rom[62027] = 12'hfff;
rom[62028] = 12'hfff;
rom[62029] = 12'hfff;
rom[62030] = 12'hfff;
rom[62031] = 12'hfff;
rom[62032] = 12'hfff;
rom[62033] = 12'hfff;
rom[62034] = 12'hfff;
rom[62035] = 12'hfff;
rom[62036] = 12'hfff;
rom[62037] = 12'hfff;
rom[62038] = 12'hfff;
rom[62039] = 12'hfff;
rom[62040] = 12'hfff;
rom[62041] = 12'hfff;
rom[62042] = 12'hfff;
rom[62043] = 12'hfff;
rom[62044] = 12'hfff;
rom[62045] = 12'hfff;
rom[62046] = 12'hfff;
rom[62047] = 12'hfff;
rom[62048] = 12'hfff;
rom[62049] = 12'hfff;
rom[62050] = 12'hfff;
rom[62051] = 12'hfff;
rom[62052] = 12'hfff;
rom[62053] = 12'hfff;
rom[62054] = 12'hfff;
rom[62055] = 12'hfff;
rom[62056] = 12'hfff;
rom[62057] = 12'hfff;
rom[62058] = 12'hfff;
rom[62059] = 12'hfff;
rom[62060] = 12'hfff;
rom[62061] = 12'hfff;
rom[62062] = 12'hfff;
rom[62063] = 12'hfff;
rom[62064] = 12'hfff;
rom[62065] = 12'hfff;
rom[62066] = 12'hfff;
rom[62067] = 12'hfff;
rom[62068] = 12'hfff;
rom[62069] = 12'hfff;
rom[62070] = 12'hfff;
rom[62071] = 12'hfff;
rom[62072] = 12'hfff;
rom[62073] = 12'hfff;
rom[62074] = 12'hfff;
rom[62075] = 12'hfff;
rom[62076] = 12'hfff;
rom[62077] = 12'hfff;
rom[62078] = 12'hfff;
rom[62079] = 12'hfff;
rom[62080] = 12'hfff;
rom[62081] = 12'hfff;
rom[62082] = 12'hfff;
rom[62083] = 12'hfff;
rom[62084] = 12'hfff;
rom[62085] = 12'hfff;
rom[62086] = 12'hfff;
rom[62087] = 12'hfff;
rom[62088] = 12'hfff;
rom[62089] = 12'hfff;
rom[62090] = 12'hfff;
rom[62091] = 12'hfff;
rom[62092] = 12'hfff;
rom[62093] = 12'hfff;
rom[62094] = 12'hfff;
rom[62095] = 12'hfff;
rom[62096] = 12'hfff;
rom[62097] = 12'hfff;
rom[62098] = 12'hfff;
rom[62099] = 12'hfff;
rom[62100] = 12'hfff;
rom[62101] = 12'hfff;
rom[62102] = 12'hfff;
rom[62103] = 12'hfff;
rom[62104] = 12'hfff;
rom[62105] = 12'hfff;
rom[62106] = 12'heee;
rom[62107] = 12'heee;
rom[62108] = 12'heee;
rom[62109] = 12'hddd;
rom[62110] = 12'hddd;
rom[62111] = 12'hddd;
rom[62112] = 12'hddd;
rom[62113] = 12'hddd;
rom[62114] = 12'hddd;
rom[62115] = 12'hddd;
rom[62116] = 12'hddd;
rom[62117] = 12'hccc;
rom[62118] = 12'hccc;
rom[62119] = 12'hccc;
rom[62120] = 12'hbbb;
rom[62121] = 12'hbbb;
rom[62122] = 12'hbbb;
rom[62123] = 12'haaa;
rom[62124] = 12'haaa;
rom[62125] = 12'h999;
rom[62126] = 12'h999;
rom[62127] = 12'h999;
rom[62128] = 12'h999;
rom[62129] = 12'h999;
rom[62130] = 12'h888;
rom[62131] = 12'h888;
rom[62132] = 12'h888;
rom[62133] = 12'h888;
rom[62134] = 12'h888;
rom[62135] = 12'h888;
rom[62136] = 12'h888;
rom[62137] = 12'h888;
rom[62138] = 12'h888;
rom[62139] = 12'h888;
rom[62140] = 12'h888;
rom[62141] = 12'h888;
rom[62142] = 12'h888;
rom[62143] = 12'h888;
rom[62144] = 12'h888;
rom[62145] = 12'h888;
rom[62146] = 12'h777;
rom[62147] = 12'h777;
rom[62148] = 12'h666;
rom[62149] = 12'h666;
rom[62150] = 12'h666;
rom[62151] = 12'h555;
rom[62152] = 12'h444;
rom[62153] = 12'h444;
rom[62154] = 12'h444;
rom[62155] = 12'h444;
rom[62156] = 12'h444;
rom[62157] = 12'h444;
rom[62158] = 12'h444;
rom[62159] = 12'h333;
rom[62160] = 12'h333;
rom[62161] = 12'h333;
rom[62162] = 12'h333;
rom[62163] = 12'h222;
rom[62164] = 12'h222;
rom[62165] = 12'h222;
rom[62166] = 12'h222;
rom[62167] = 12'h222;
rom[62168] = 12'h111;
rom[62169] = 12'h111;
rom[62170] = 12'h111;
rom[62171] = 12'h111;
rom[62172] = 12'h111;
rom[62173] = 12'h111;
rom[62174] = 12'h111;
rom[62175] = 12'h111;
rom[62176] = 12'h  0;
rom[62177] = 12'h  0;
rom[62178] = 12'h  0;
rom[62179] = 12'h  0;
rom[62180] = 12'h  0;
rom[62181] = 12'h  0;
rom[62182] = 12'h  0;
rom[62183] = 12'h  0;
rom[62184] = 12'h  0;
rom[62185] = 12'h  0;
rom[62186] = 12'h  0;
rom[62187] = 12'h  0;
rom[62188] = 12'h  0;
rom[62189] = 12'h  0;
rom[62190] = 12'h  0;
rom[62191] = 12'h  0;
rom[62192] = 12'h  0;
rom[62193] = 12'h  0;
rom[62194] = 12'h  0;
rom[62195] = 12'h  0;
rom[62196] = 12'h  0;
rom[62197] = 12'h  0;
rom[62198] = 12'h  0;
rom[62199] = 12'h  0;
rom[62200] = 12'h  0;
rom[62201] = 12'h  0;
rom[62202] = 12'h  0;
rom[62203] = 12'h  0;
rom[62204] = 12'h  0;
rom[62205] = 12'h  0;
rom[62206] = 12'h  0;
rom[62207] = 12'h  0;
rom[62208] = 12'h  0;
rom[62209] = 12'h  0;
rom[62210] = 12'h111;
rom[62211] = 12'h111;
rom[62212] = 12'h222;
rom[62213] = 12'h222;
rom[62214] = 12'h222;
rom[62215] = 12'h111;
rom[62216] = 12'h111;
rom[62217] = 12'h111;
rom[62218] = 12'h111;
rom[62219] = 12'h111;
rom[62220] = 12'h111;
rom[62221] = 12'h111;
rom[62222] = 12'h111;
rom[62223] = 12'h  0;
rom[62224] = 12'h  0;
rom[62225] = 12'h  0;
rom[62226] = 12'h  0;
rom[62227] = 12'h  0;
rom[62228] = 12'h  0;
rom[62229] = 12'h  0;
rom[62230] = 12'h  0;
rom[62231] = 12'h  0;
rom[62232] = 12'h  0;
rom[62233] = 12'h  0;
rom[62234] = 12'h  0;
rom[62235] = 12'h  0;
rom[62236] = 12'h  0;
rom[62237] = 12'h  0;
rom[62238] = 12'h  0;
rom[62239] = 12'h  0;
rom[62240] = 12'h  0;
rom[62241] = 12'h  0;
rom[62242] = 12'h  0;
rom[62243] = 12'h  0;
rom[62244] = 12'h  0;
rom[62245] = 12'h  0;
rom[62246] = 12'h  0;
rom[62247] = 12'h  0;
rom[62248] = 12'h  0;
rom[62249] = 12'h  0;
rom[62250] = 12'h  0;
rom[62251] = 12'h  0;
rom[62252] = 12'h  0;
rom[62253] = 12'h  0;
rom[62254] = 12'h  0;
rom[62255] = 12'h  0;
rom[62256] = 12'h  0;
rom[62257] = 12'h  0;
rom[62258] = 12'h  0;
rom[62259] = 12'h  0;
rom[62260] = 12'h  0;
rom[62261] = 12'h  0;
rom[62262] = 12'h  0;
rom[62263] = 12'h  0;
rom[62264] = 12'h  0;
rom[62265] = 12'h  0;
rom[62266] = 12'h  0;
rom[62267] = 12'h  0;
rom[62268] = 12'h  0;
rom[62269] = 12'h  0;
rom[62270] = 12'h  0;
rom[62271] = 12'h  0;
rom[62272] = 12'h  0;
rom[62273] = 12'h111;
rom[62274] = 12'h111;
rom[62275] = 12'h222;
rom[62276] = 12'h222;
rom[62277] = 12'h333;
rom[62278] = 12'h444;
rom[62279] = 12'h444;
rom[62280] = 12'h444;
rom[62281] = 12'h555;
rom[62282] = 12'h555;
rom[62283] = 12'h444;
rom[62284] = 12'h333;
rom[62285] = 12'h222;
rom[62286] = 12'h222;
rom[62287] = 12'h222;
rom[62288] = 12'h222;
rom[62289] = 12'h222;
rom[62290] = 12'h222;
rom[62291] = 12'h222;
rom[62292] = 12'h222;
rom[62293] = 12'h222;
rom[62294] = 12'h222;
rom[62295] = 12'h222;
rom[62296] = 12'h222;
rom[62297] = 12'h333;
rom[62298] = 12'h555;
rom[62299] = 12'h555;
rom[62300] = 12'h555;
rom[62301] = 12'h444;
rom[62302] = 12'h444;
rom[62303] = 12'h333;
rom[62304] = 12'h444;
rom[62305] = 12'h444;
rom[62306] = 12'h444;
rom[62307] = 12'h555;
rom[62308] = 12'h555;
rom[62309] = 12'h666;
rom[62310] = 12'h666;
rom[62311] = 12'h666;
rom[62312] = 12'h777;
rom[62313] = 12'h777;
rom[62314] = 12'h777;
rom[62315] = 12'h666;
rom[62316] = 12'h666;
rom[62317] = 12'h666;
rom[62318] = 12'h666;
rom[62319] = 12'h666;
rom[62320] = 12'h666;
rom[62321] = 12'h666;
rom[62322] = 12'h666;
rom[62323] = 12'h777;
rom[62324] = 12'h777;
rom[62325] = 12'h777;
rom[62326] = 12'h777;
rom[62327] = 12'h777;
rom[62328] = 12'h888;
rom[62329] = 12'h888;
rom[62330] = 12'h888;
rom[62331] = 12'h888;
rom[62332] = 12'h888;
rom[62333] = 12'h999;
rom[62334] = 12'h999;
rom[62335] = 12'h999;
rom[62336] = 12'h999;
rom[62337] = 12'h999;
rom[62338] = 12'haaa;
rom[62339] = 12'haaa;
rom[62340] = 12'haaa;
rom[62341] = 12'haaa;
rom[62342] = 12'haaa;
rom[62343] = 12'hbbb;
rom[62344] = 12'hbbb;
rom[62345] = 12'hbbb;
rom[62346] = 12'hccc;
rom[62347] = 12'hccc;
rom[62348] = 12'hddd;
rom[62349] = 12'hddd;
rom[62350] = 12'hddd;
rom[62351] = 12'heee;
rom[62352] = 12'hfff;
rom[62353] = 12'hfff;
rom[62354] = 12'hfff;
rom[62355] = 12'hfff;
rom[62356] = 12'heee;
rom[62357] = 12'heee;
rom[62358] = 12'hddd;
rom[62359] = 12'hddd;
rom[62360] = 12'hccc;
rom[62361] = 12'hccc;
rom[62362] = 12'hccc;
rom[62363] = 12'hbbb;
rom[62364] = 12'hbbb;
rom[62365] = 12'hbbb;
rom[62366] = 12'hbbb;
rom[62367] = 12'hbbb;
rom[62368] = 12'hbbb;
rom[62369] = 12'hbbb;
rom[62370] = 12'hbbb;
rom[62371] = 12'hbbb;
rom[62372] = 12'hbbb;
rom[62373] = 12'hbbb;
rom[62374] = 12'hbbb;
rom[62375] = 12'haaa;
rom[62376] = 12'h999;
rom[62377] = 12'h999;
rom[62378] = 12'h999;
rom[62379] = 12'h888;
rom[62380] = 12'h888;
rom[62381] = 12'h888;
rom[62382] = 12'h888;
rom[62383] = 12'h777;
rom[62384] = 12'h777;
rom[62385] = 12'h777;
rom[62386] = 12'h777;
rom[62387] = 12'h777;
rom[62388] = 12'h777;
rom[62389] = 12'h777;
rom[62390] = 12'h666;
rom[62391] = 12'h666;
rom[62392] = 12'h777;
rom[62393] = 12'h777;
rom[62394] = 12'h777;
rom[62395] = 12'h777;
rom[62396] = 12'h777;
rom[62397] = 12'h777;
rom[62398] = 12'h777;
rom[62399] = 12'h777;
rom[62400] = 12'hfff;
rom[62401] = 12'hfff;
rom[62402] = 12'hfff;
rom[62403] = 12'hfff;
rom[62404] = 12'hfff;
rom[62405] = 12'hfff;
rom[62406] = 12'hfff;
rom[62407] = 12'hfff;
rom[62408] = 12'hfff;
rom[62409] = 12'hfff;
rom[62410] = 12'hfff;
rom[62411] = 12'hfff;
rom[62412] = 12'hfff;
rom[62413] = 12'hfff;
rom[62414] = 12'hfff;
rom[62415] = 12'hfff;
rom[62416] = 12'hfff;
rom[62417] = 12'hfff;
rom[62418] = 12'hfff;
rom[62419] = 12'hfff;
rom[62420] = 12'hfff;
rom[62421] = 12'hfff;
rom[62422] = 12'hfff;
rom[62423] = 12'hfff;
rom[62424] = 12'hfff;
rom[62425] = 12'hfff;
rom[62426] = 12'hfff;
rom[62427] = 12'hfff;
rom[62428] = 12'hfff;
rom[62429] = 12'hfff;
rom[62430] = 12'hfff;
rom[62431] = 12'hfff;
rom[62432] = 12'hfff;
rom[62433] = 12'hfff;
rom[62434] = 12'hfff;
rom[62435] = 12'hfff;
rom[62436] = 12'hfff;
rom[62437] = 12'hfff;
rom[62438] = 12'hfff;
rom[62439] = 12'hfff;
rom[62440] = 12'hfff;
rom[62441] = 12'hfff;
rom[62442] = 12'hfff;
rom[62443] = 12'hfff;
rom[62444] = 12'hfff;
rom[62445] = 12'hfff;
rom[62446] = 12'hfff;
rom[62447] = 12'hfff;
rom[62448] = 12'hfff;
rom[62449] = 12'hfff;
rom[62450] = 12'hfff;
rom[62451] = 12'hfff;
rom[62452] = 12'hfff;
rom[62453] = 12'hfff;
rom[62454] = 12'hfff;
rom[62455] = 12'hfff;
rom[62456] = 12'hfff;
rom[62457] = 12'hfff;
rom[62458] = 12'hfff;
rom[62459] = 12'hfff;
rom[62460] = 12'hfff;
rom[62461] = 12'hfff;
rom[62462] = 12'hfff;
rom[62463] = 12'hfff;
rom[62464] = 12'hfff;
rom[62465] = 12'hfff;
rom[62466] = 12'hfff;
rom[62467] = 12'hfff;
rom[62468] = 12'hfff;
rom[62469] = 12'hfff;
rom[62470] = 12'hfff;
rom[62471] = 12'hfff;
rom[62472] = 12'hfff;
rom[62473] = 12'hfff;
rom[62474] = 12'hfff;
rom[62475] = 12'hfff;
rom[62476] = 12'hfff;
rom[62477] = 12'hfff;
rom[62478] = 12'hfff;
rom[62479] = 12'hfff;
rom[62480] = 12'hfff;
rom[62481] = 12'hfff;
rom[62482] = 12'hfff;
rom[62483] = 12'hfff;
rom[62484] = 12'hfff;
rom[62485] = 12'hfff;
rom[62486] = 12'hfff;
rom[62487] = 12'hfff;
rom[62488] = 12'hfff;
rom[62489] = 12'hfff;
rom[62490] = 12'hfff;
rom[62491] = 12'hfff;
rom[62492] = 12'hfff;
rom[62493] = 12'hfff;
rom[62494] = 12'hfff;
rom[62495] = 12'hfff;
rom[62496] = 12'hfff;
rom[62497] = 12'hfff;
rom[62498] = 12'hfff;
rom[62499] = 12'hfff;
rom[62500] = 12'hfff;
rom[62501] = 12'hfff;
rom[62502] = 12'hfff;
rom[62503] = 12'hfff;
rom[62504] = 12'hfff;
rom[62505] = 12'hfff;
rom[62506] = 12'hfff;
rom[62507] = 12'hfff;
rom[62508] = 12'heee;
rom[62509] = 12'heee;
rom[62510] = 12'heee;
rom[62511] = 12'heee;
rom[62512] = 12'heee;
rom[62513] = 12'heee;
rom[62514] = 12'hddd;
rom[62515] = 12'hddd;
rom[62516] = 12'hddd;
rom[62517] = 12'hddd;
rom[62518] = 12'hccc;
rom[62519] = 12'hccc;
rom[62520] = 12'hbbb;
rom[62521] = 12'hbbb;
rom[62522] = 12'hbbb;
rom[62523] = 12'haaa;
rom[62524] = 12'haaa;
rom[62525] = 12'h999;
rom[62526] = 12'h999;
rom[62527] = 12'h999;
rom[62528] = 12'h999;
rom[62529] = 12'h999;
rom[62530] = 12'h888;
rom[62531] = 12'h888;
rom[62532] = 12'h888;
rom[62533] = 12'h888;
rom[62534] = 12'h888;
rom[62535] = 12'h777;
rom[62536] = 12'h777;
rom[62537] = 12'h777;
rom[62538] = 12'h777;
rom[62539] = 12'h777;
rom[62540] = 12'h888;
rom[62541] = 12'h777;
rom[62542] = 12'h777;
rom[62543] = 12'h777;
rom[62544] = 12'h777;
rom[62545] = 12'h777;
rom[62546] = 12'h777;
rom[62547] = 12'h777;
rom[62548] = 12'h777;
rom[62549] = 12'h777;
rom[62550] = 12'h777;
rom[62551] = 12'h666;
rom[62552] = 12'h555;
rom[62553] = 12'h555;
rom[62554] = 12'h555;
rom[62555] = 12'h444;
rom[62556] = 12'h444;
rom[62557] = 12'h444;
rom[62558] = 12'h444;
rom[62559] = 12'h444;
rom[62560] = 12'h333;
rom[62561] = 12'h333;
rom[62562] = 12'h333;
rom[62563] = 12'h222;
rom[62564] = 12'h222;
rom[62565] = 12'h222;
rom[62566] = 12'h222;
rom[62567] = 12'h222;
rom[62568] = 12'h111;
rom[62569] = 12'h111;
rom[62570] = 12'h111;
rom[62571] = 12'h111;
rom[62572] = 12'h111;
rom[62573] = 12'h111;
rom[62574] = 12'h111;
rom[62575] = 12'h111;
rom[62576] = 12'h111;
rom[62577] = 12'h111;
rom[62578] = 12'h  0;
rom[62579] = 12'h  0;
rom[62580] = 12'h  0;
rom[62581] = 12'h  0;
rom[62582] = 12'h  0;
rom[62583] = 12'h  0;
rom[62584] = 12'h  0;
rom[62585] = 12'h  0;
rom[62586] = 12'h  0;
rom[62587] = 12'h  0;
rom[62588] = 12'h  0;
rom[62589] = 12'h  0;
rom[62590] = 12'h  0;
rom[62591] = 12'h  0;
rom[62592] = 12'h  0;
rom[62593] = 12'h  0;
rom[62594] = 12'h  0;
rom[62595] = 12'h  0;
rom[62596] = 12'h  0;
rom[62597] = 12'h  0;
rom[62598] = 12'h  0;
rom[62599] = 12'h  0;
rom[62600] = 12'h  0;
rom[62601] = 12'h  0;
rom[62602] = 12'h  0;
rom[62603] = 12'h  0;
rom[62604] = 12'h  0;
rom[62605] = 12'h  0;
rom[62606] = 12'h  0;
rom[62607] = 12'h  0;
rom[62608] = 12'h  0;
rom[62609] = 12'h  0;
rom[62610] = 12'h111;
rom[62611] = 12'h111;
rom[62612] = 12'h222;
rom[62613] = 12'h222;
rom[62614] = 12'h111;
rom[62615] = 12'h111;
rom[62616] = 12'h111;
rom[62617] = 12'h111;
rom[62618] = 12'h111;
rom[62619] = 12'h111;
rom[62620] = 12'h111;
rom[62621] = 12'h111;
rom[62622] = 12'h111;
rom[62623] = 12'h  0;
rom[62624] = 12'h  0;
rom[62625] = 12'h  0;
rom[62626] = 12'h  0;
rom[62627] = 12'h  0;
rom[62628] = 12'h  0;
rom[62629] = 12'h  0;
rom[62630] = 12'h  0;
rom[62631] = 12'h  0;
rom[62632] = 12'h  0;
rom[62633] = 12'h  0;
rom[62634] = 12'h  0;
rom[62635] = 12'h  0;
rom[62636] = 12'h  0;
rom[62637] = 12'h  0;
rom[62638] = 12'h  0;
rom[62639] = 12'h  0;
rom[62640] = 12'h  0;
rom[62641] = 12'h  0;
rom[62642] = 12'h  0;
rom[62643] = 12'h  0;
rom[62644] = 12'h  0;
rom[62645] = 12'h  0;
rom[62646] = 12'h  0;
rom[62647] = 12'h  0;
rom[62648] = 12'h  0;
rom[62649] = 12'h  0;
rom[62650] = 12'h  0;
rom[62651] = 12'h  0;
rom[62652] = 12'h  0;
rom[62653] = 12'h  0;
rom[62654] = 12'h  0;
rom[62655] = 12'h  0;
rom[62656] = 12'h  0;
rom[62657] = 12'h  0;
rom[62658] = 12'h  0;
rom[62659] = 12'h  0;
rom[62660] = 12'h  0;
rom[62661] = 12'h  0;
rom[62662] = 12'h  0;
rom[62663] = 12'h  0;
rom[62664] = 12'h  0;
rom[62665] = 12'h  0;
rom[62666] = 12'h  0;
rom[62667] = 12'h  0;
rom[62668] = 12'h  0;
rom[62669] = 12'h  0;
rom[62670] = 12'h  0;
rom[62671] = 12'h  0;
rom[62672] = 12'h  0;
rom[62673] = 12'h111;
rom[62674] = 12'h111;
rom[62675] = 12'h222;
rom[62676] = 12'h222;
rom[62677] = 12'h333;
rom[62678] = 12'h444;
rom[62679] = 12'h444;
rom[62680] = 12'h555;
rom[62681] = 12'h555;
rom[62682] = 12'h444;
rom[62683] = 12'h444;
rom[62684] = 12'h333;
rom[62685] = 12'h222;
rom[62686] = 12'h222;
rom[62687] = 12'h222;
rom[62688] = 12'h222;
rom[62689] = 12'h222;
rom[62690] = 12'h222;
rom[62691] = 12'h111;
rom[62692] = 12'h222;
rom[62693] = 12'h222;
rom[62694] = 12'h222;
rom[62695] = 12'h222;
rom[62696] = 12'h222;
rom[62697] = 12'h333;
rom[62698] = 12'h444;
rom[62699] = 12'h555;
rom[62700] = 12'h555;
rom[62701] = 12'h444;
rom[62702] = 12'h444;
rom[62703] = 12'h333;
rom[62704] = 12'h444;
rom[62705] = 12'h444;
rom[62706] = 12'h444;
rom[62707] = 12'h444;
rom[62708] = 12'h555;
rom[62709] = 12'h555;
rom[62710] = 12'h666;
rom[62711] = 12'h666;
rom[62712] = 12'h777;
rom[62713] = 12'h777;
rom[62714] = 12'h777;
rom[62715] = 12'h777;
rom[62716] = 12'h777;
rom[62717] = 12'h777;
rom[62718] = 12'h666;
rom[62719] = 12'h666;
rom[62720] = 12'h666;
rom[62721] = 12'h666;
rom[62722] = 12'h777;
rom[62723] = 12'h777;
rom[62724] = 12'h777;
rom[62725] = 12'h777;
rom[62726] = 12'h777;
rom[62727] = 12'h888;
rom[62728] = 12'h888;
rom[62729] = 12'h888;
rom[62730] = 12'h888;
rom[62731] = 12'h888;
rom[62732] = 12'h999;
rom[62733] = 12'h999;
rom[62734] = 12'h999;
rom[62735] = 12'h999;
rom[62736] = 12'h999;
rom[62737] = 12'haaa;
rom[62738] = 12'haaa;
rom[62739] = 12'haaa;
rom[62740] = 12'haaa;
rom[62741] = 12'haaa;
rom[62742] = 12'hbbb;
rom[62743] = 12'hbbb;
rom[62744] = 12'hbbb;
rom[62745] = 12'hccc;
rom[62746] = 12'hccc;
rom[62747] = 12'hccc;
rom[62748] = 12'hddd;
rom[62749] = 12'hddd;
rom[62750] = 12'heee;
rom[62751] = 12'heee;
rom[62752] = 12'hfff;
rom[62753] = 12'hfff;
rom[62754] = 12'hfff;
rom[62755] = 12'hfff;
rom[62756] = 12'heee;
rom[62757] = 12'hddd;
rom[62758] = 12'hddd;
rom[62759] = 12'hccc;
rom[62760] = 12'hccc;
rom[62761] = 12'hccc;
rom[62762] = 12'hbbb;
rom[62763] = 12'hbbb;
rom[62764] = 12'hbbb;
rom[62765] = 12'hbbb;
rom[62766] = 12'hbbb;
rom[62767] = 12'hbbb;
rom[62768] = 12'hbbb;
rom[62769] = 12'hbbb;
rom[62770] = 12'hbbb;
rom[62771] = 12'hbbb;
rom[62772] = 12'hccc;
rom[62773] = 12'hbbb;
rom[62774] = 12'hbbb;
rom[62775] = 12'hbbb;
rom[62776] = 12'haaa;
rom[62777] = 12'h999;
rom[62778] = 12'h999;
rom[62779] = 12'h999;
rom[62780] = 12'h888;
rom[62781] = 12'h888;
rom[62782] = 12'h777;
rom[62783] = 12'h777;
rom[62784] = 12'h777;
rom[62785] = 12'h777;
rom[62786] = 12'h777;
rom[62787] = 12'h777;
rom[62788] = 12'h777;
rom[62789] = 12'h777;
rom[62790] = 12'h777;
rom[62791] = 12'h777;
rom[62792] = 12'h777;
rom[62793] = 12'h777;
rom[62794] = 12'h777;
rom[62795] = 12'h777;
rom[62796] = 12'h777;
rom[62797] = 12'h777;
rom[62798] = 12'h777;
rom[62799] = 12'h777;
rom[62800] = 12'hfff;
rom[62801] = 12'hfff;
rom[62802] = 12'hfff;
rom[62803] = 12'hfff;
rom[62804] = 12'hfff;
rom[62805] = 12'hfff;
rom[62806] = 12'hfff;
rom[62807] = 12'hfff;
rom[62808] = 12'hfff;
rom[62809] = 12'hfff;
rom[62810] = 12'hfff;
rom[62811] = 12'hfff;
rom[62812] = 12'hfff;
rom[62813] = 12'hfff;
rom[62814] = 12'hfff;
rom[62815] = 12'hfff;
rom[62816] = 12'hfff;
rom[62817] = 12'hfff;
rom[62818] = 12'hfff;
rom[62819] = 12'hfff;
rom[62820] = 12'hfff;
rom[62821] = 12'hfff;
rom[62822] = 12'hfff;
rom[62823] = 12'hfff;
rom[62824] = 12'hfff;
rom[62825] = 12'hfff;
rom[62826] = 12'hfff;
rom[62827] = 12'hfff;
rom[62828] = 12'hfff;
rom[62829] = 12'hfff;
rom[62830] = 12'hfff;
rom[62831] = 12'hfff;
rom[62832] = 12'hfff;
rom[62833] = 12'hfff;
rom[62834] = 12'hfff;
rom[62835] = 12'hfff;
rom[62836] = 12'hfff;
rom[62837] = 12'hfff;
rom[62838] = 12'hfff;
rom[62839] = 12'hfff;
rom[62840] = 12'hfff;
rom[62841] = 12'hfff;
rom[62842] = 12'hfff;
rom[62843] = 12'hfff;
rom[62844] = 12'hfff;
rom[62845] = 12'hfff;
rom[62846] = 12'hfff;
rom[62847] = 12'hfff;
rom[62848] = 12'hfff;
rom[62849] = 12'hfff;
rom[62850] = 12'hfff;
rom[62851] = 12'hfff;
rom[62852] = 12'hfff;
rom[62853] = 12'hfff;
rom[62854] = 12'hfff;
rom[62855] = 12'hfff;
rom[62856] = 12'hfff;
rom[62857] = 12'hfff;
rom[62858] = 12'hfff;
rom[62859] = 12'hfff;
rom[62860] = 12'hfff;
rom[62861] = 12'hfff;
rom[62862] = 12'hfff;
rom[62863] = 12'hfff;
rom[62864] = 12'hfff;
rom[62865] = 12'hfff;
rom[62866] = 12'hfff;
rom[62867] = 12'hfff;
rom[62868] = 12'hfff;
rom[62869] = 12'hfff;
rom[62870] = 12'hfff;
rom[62871] = 12'hfff;
rom[62872] = 12'hfff;
rom[62873] = 12'hfff;
rom[62874] = 12'hfff;
rom[62875] = 12'hfff;
rom[62876] = 12'hfff;
rom[62877] = 12'hfff;
rom[62878] = 12'hfff;
rom[62879] = 12'hfff;
rom[62880] = 12'hfff;
rom[62881] = 12'hfff;
rom[62882] = 12'hfff;
rom[62883] = 12'hfff;
rom[62884] = 12'hfff;
rom[62885] = 12'hfff;
rom[62886] = 12'hfff;
rom[62887] = 12'hfff;
rom[62888] = 12'hfff;
rom[62889] = 12'hfff;
rom[62890] = 12'hfff;
rom[62891] = 12'hfff;
rom[62892] = 12'hfff;
rom[62893] = 12'hfff;
rom[62894] = 12'hfff;
rom[62895] = 12'hfff;
rom[62896] = 12'hfff;
rom[62897] = 12'hfff;
rom[62898] = 12'hfff;
rom[62899] = 12'hfff;
rom[62900] = 12'hfff;
rom[62901] = 12'hfff;
rom[62902] = 12'hfff;
rom[62903] = 12'hfff;
rom[62904] = 12'hfff;
rom[62905] = 12'hfff;
rom[62906] = 12'hfff;
rom[62907] = 12'hfff;
rom[62908] = 12'hfff;
rom[62909] = 12'hfff;
rom[62910] = 12'heee;
rom[62911] = 12'heee;
rom[62912] = 12'heee;
rom[62913] = 12'heee;
rom[62914] = 12'heee;
rom[62915] = 12'hddd;
rom[62916] = 12'hddd;
rom[62917] = 12'hddd;
rom[62918] = 12'hddd;
rom[62919] = 12'hddd;
rom[62920] = 12'hccc;
rom[62921] = 12'hccc;
rom[62922] = 12'hbbb;
rom[62923] = 12'hbbb;
rom[62924] = 12'hbbb;
rom[62925] = 12'haaa;
rom[62926] = 12'haaa;
rom[62927] = 12'haaa;
rom[62928] = 12'h999;
rom[62929] = 12'h999;
rom[62930] = 12'h888;
rom[62931] = 12'h888;
rom[62932] = 12'h888;
rom[62933] = 12'h888;
rom[62934] = 12'h888;
rom[62935] = 12'h777;
rom[62936] = 12'h777;
rom[62937] = 12'h777;
rom[62938] = 12'h777;
rom[62939] = 12'h777;
rom[62940] = 12'h777;
rom[62941] = 12'h777;
rom[62942] = 12'h777;
rom[62943] = 12'h777;
rom[62944] = 12'h777;
rom[62945] = 12'h777;
rom[62946] = 12'h777;
rom[62947] = 12'h777;
rom[62948] = 12'h777;
rom[62949] = 12'h777;
rom[62950] = 12'h777;
rom[62951] = 12'h666;
rom[62952] = 12'h666;
rom[62953] = 12'h666;
rom[62954] = 12'h555;
rom[62955] = 12'h555;
rom[62956] = 12'h555;
rom[62957] = 12'h444;
rom[62958] = 12'h444;
rom[62959] = 12'h444;
rom[62960] = 12'h333;
rom[62961] = 12'h333;
rom[62962] = 12'h333;
rom[62963] = 12'h222;
rom[62964] = 12'h222;
rom[62965] = 12'h222;
rom[62966] = 12'h222;
rom[62967] = 12'h222;
rom[62968] = 12'h111;
rom[62969] = 12'h111;
rom[62970] = 12'h111;
rom[62971] = 12'h111;
rom[62972] = 12'h111;
rom[62973] = 12'h111;
rom[62974] = 12'h111;
rom[62975] = 12'h111;
rom[62976] = 12'h111;
rom[62977] = 12'h111;
rom[62978] = 12'h  0;
rom[62979] = 12'h  0;
rom[62980] = 12'h  0;
rom[62981] = 12'h  0;
rom[62982] = 12'h  0;
rom[62983] = 12'h  0;
rom[62984] = 12'h  0;
rom[62985] = 12'h  0;
rom[62986] = 12'h  0;
rom[62987] = 12'h  0;
rom[62988] = 12'h  0;
rom[62989] = 12'h  0;
rom[62990] = 12'h  0;
rom[62991] = 12'h  0;
rom[62992] = 12'h  0;
rom[62993] = 12'h  0;
rom[62994] = 12'h  0;
rom[62995] = 12'h  0;
rom[62996] = 12'h  0;
rom[62997] = 12'h  0;
rom[62998] = 12'h  0;
rom[62999] = 12'h  0;
rom[63000] = 12'h  0;
rom[63001] = 12'h  0;
rom[63002] = 12'h  0;
rom[63003] = 12'h  0;
rom[63004] = 12'h  0;
rom[63005] = 12'h  0;
rom[63006] = 12'h  0;
rom[63007] = 12'h  0;
rom[63008] = 12'h  0;
rom[63009] = 12'h  0;
rom[63010] = 12'h111;
rom[63011] = 12'h111;
rom[63012] = 12'h222;
rom[63013] = 12'h222;
rom[63014] = 12'h111;
rom[63015] = 12'h111;
rom[63016] = 12'h111;
rom[63017] = 12'h111;
rom[63018] = 12'h111;
rom[63019] = 12'h  0;
rom[63020] = 12'h111;
rom[63021] = 12'h111;
rom[63022] = 12'h  0;
rom[63023] = 12'h  0;
rom[63024] = 12'h  0;
rom[63025] = 12'h  0;
rom[63026] = 12'h  0;
rom[63027] = 12'h  0;
rom[63028] = 12'h  0;
rom[63029] = 12'h  0;
rom[63030] = 12'h  0;
rom[63031] = 12'h  0;
rom[63032] = 12'h  0;
rom[63033] = 12'h  0;
rom[63034] = 12'h  0;
rom[63035] = 12'h  0;
rom[63036] = 12'h  0;
rom[63037] = 12'h  0;
rom[63038] = 12'h  0;
rom[63039] = 12'h  0;
rom[63040] = 12'h  0;
rom[63041] = 12'h  0;
rom[63042] = 12'h  0;
rom[63043] = 12'h  0;
rom[63044] = 12'h  0;
rom[63045] = 12'h  0;
rom[63046] = 12'h  0;
rom[63047] = 12'h  0;
rom[63048] = 12'h  0;
rom[63049] = 12'h  0;
rom[63050] = 12'h  0;
rom[63051] = 12'h  0;
rom[63052] = 12'h  0;
rom[63053] = 12'h  0;
rom[63054] = 12'h  0;
rom[63055] = 12'h  0;
rom[63056] = 12'h  0;
rom[63057] = 12'h  0;
rom[63058] = 12'h  0;
rom[63059] = 12'h  0;
rom[63060] = 12'h  0;
rom[63061] = 12'h  0;
rom[63062] = 12'h  0;
rom[63063] = 12'h  0;
rom[63064] = 12'h  0;
rom[63065] = 12'h  0;
rom[63066] = 12'h  0;
rom[63067] = 12'h  0;
rom[63068] = 12'h  0;
rom[63069] = 12'h  0;
rom[63070] = 12'h  0;
rom[63071] = 12'h  0;
rom[63072] = 12'h  0;
rom[63073] = 12'h111;
rom[63074] = 12'h111;
rom[63075] = 12'h222;
rom[63076] = 12'h222;
rom[63077] = 12'h333;
rom[63078] = 12'h444;
rom[63079] = 12'h444;
rom[63080] = 12'h555;
rom[63081] = 12'h555;
rom[63082] = 12'h444;
rom[63083] = 12'h333;
rom[63084] = 12'h222;
rom[63085] = 12'h222;
rom[63086] = 12'h222;
rom[63087] = 12'h222;
rom[63088] = 12'h111;
rom[63089] = 12'h222;
rom[63090] = 12'h111;
rom[63091] = 12'h111;
rom[63092] = 12'h111;
rom[63093] = 12'h222;
rom[63094] = 12'h222;
rom[63095] = 12'h111;
rom[63096] = 12'h222;
rom[63097] = 12'h333;
rom[63098] = 12'h444;
rom[63099] = 12'h555;
rom[63100] = 12'h555;
rom[63101] = 12'h444;
rom[63102] = 12'h444;
rom[63103] = 12'h333;
rom[63104] = 12'h444;
rom[63105] = 12'h444;
rom[63106] = 12'h444;
rom[63107] = 12'h444;
rom[63108] = 12'h444;
rom[63109] = 12'h555;
rom[63110] = 12'h555;
rom[63111] = 12'h666;
rom[63112] = 12'h666;
rom[63113] = 12'h777;
rom[63114] = 12'h777;
rom[63115] = 12'h777;
rom[63116] = 12'h777;
rom[63117] = 12'h777;
rom[63118] = 12'h777;
rom[63119] = 12'h777;
rom[63120] = 12'h777;
rom[63121] = 12'h777;
rom[63122] = 12'h777;
rom[63123] = 12'h777;
rom[63124] = 12'h777;
rom[63125] = 12'h777;
rom[63126] = 12'h888;
rom[63127] = 12'h888;
rom[63128] = 12'h888;
rom[63129] = 12'h888;
rom[63130] = 12'h888;
rom[63131] = 12'h888;
rom[63132] = 12'h999;
rom[63133] = 12'h999;
rom[63134] = 12'h999;
rom[63135] = 12'h999;
rom[63136] = 12'h999;
rom[63137] = 12'haaa;
rom[63138] = 12'haaa;
rom[63139] = 12'haaa;
rom[63140] = 12'haaa;
rom[63141] = 12'hbbb;
rom[63142] = 12'hbbb;
rom[63143] = 12'hbbb;
rom[63144] = 12'hbbb;
rom[63145] = 12'hccc;
rom[63146] = 12'hccc;
rom[63147] = 12'hddd;
rom[63148] = 12'hddd;
rom[63149] = 12'heee;
rom[63150] = 12'heee;
rom[63151] = 12'hfff;
rom[63152] = 12'hfff;
rom[63153] = 12'hfff;
rom[63154] = 12'hfff;
rom[63155] = 12'heee;
rom[63156] = 12'heee;
rom[63157] = 12'hddd;
rom[63158] = 12'hccc;
rom[63159] = 12'hccc;
rom[63160] = 12'hccc;
rom[63161] = 12'hccc;
rom[63162] = 12'hbbb;
rom[63163] = 12'hbbb;
rom[63164] = 12'hbbb;
rom[63165] = 12'hbbb;
rom[63166] = 12'hbbb;
rom[63167] = 12'hbbb;
rom[63168] = 12'hbbb;
rom[63169] = 12'hbbb;
rom[63170] = 12'hbbb;
rom[63171] = 12'hbbb;
rom[63172] = 12'hccc;
rom[63173] = 12'hbbb;
rom[63174] = 12'hbbb;
rom[63175] = 12'hbbb;
rom[63176] = 12'haaa;
rom[63177] = 12'haaa;
rom[63178] = 12'h999;
rom[63179] = 12'h999;
rom[63180] = 12'h888;
rom[63181] = 12'h888;
rom[63182] = 12'h777;
rom[63183] = 12'h777;
rom[63184] = 12'h777;
rom[63185] = 12'h777;
rom[63186] = 12'h777;
rom[63187] = 12'h777;
rom[63188] = 12'h777;
rom[63189] = 12'h777;
rom[63190] = 12'h777;
rom[63191] = 12'h777;
rom[63192] = 12'h777;
rom[63193] = 12'h777;
rom[63194] = 12'h777;
rom[63195] = 12'h777;
rom[63196] = 12'h777;
rom[63197] = 12'h777;
rom[63198] = 12'h777;
rom[63199] = 12'h777;
rom[63200] = 12'hfff;
rom[63201] = 12'hfff;
rom[63202] = 12'hfff;
rom[63203] = 12'hfff;
rom[63204] = 12'hfff;
rom[63205] = 12'hfff;
rom[63206] = 12'hfff;
rom[63207] = 12'hfff;
rom[63208] = 12'hfff;
rom[63209] = 12'hfff;
rom[63210] = 12'hfff;
rom[63211] = 12'hfff;
rom[63212] = 12'hfff;
rom[63213] = 12'hfff;
rom[63214] = 12'hfff;
rom[63215] = 12'hfff;
rom[63216] = 12'hfff;
rom[63217] = 12'hfff;
rom[63218] = 12'hfff;
rom[63219] = 12'hfff;
rom[63220] = 12'hfff;
rom[63221] = 12'hfff;
rom[63222] = 12'hfff;
rom[63223] = 12'hfff;
rom[63224] = 12'hfff;
rom[63225] = 12'hfff;
rom[63226] = 12'hfff;
rom[63227] = 12'hfff;
rom[63228] = 12'hfff;
rom[63229] = 12'hfff;
rom[63230] = 12'hfff;
rom[63231] = 12'hfff;
rom[63232] = 12'hfff;
rom[63233] = 12'hfff;
rom[63234] = 12'hfff;
rom[63235] = 12'hfff;
rom[63236] = 12'hfff;
rom[63237] = 12'hfff;
rom[63238] = 12'hfff;
rom[63239] = 12'hfff;
rom[63240] = 12'hfff;
rom[63241] = 12'hfff;
rom[63242] = 12'hfff;
rom[63243] = 12'hfff;
rom[63244] = 12'hfff;
rom[63245] = 12'hfff;
rom[63246] = 12'hfff;
rom[63247] = 12'hfff;
rom[63248] = 12'hfff;
rom[63249] = 12'hfff;
rom[63250] = 12'hfff;
rom[63251] = 12'hfff;
rom[63252] = 12'hfff;
rom[63253] = 12'hfff;
rom[63254] = 12'hfff;
rom[63255] = 12'hfff;
rom[63256] = 12'hfff;
rom[63257] = 12'hfff;
rom[63258] = 12'hfff;
rom[63259] = 12'hfff;
rom[63260] = 12'hfff;
rom[63261] = 12'hfff;
rom[63262] = 12'hfff;
rom[63263] = 12'hfff;
rom[63264] = 12'hfff;
rom[63265] = 12'hfff;
rom[63266] = 12'hfff;
rom[63267] = 12'hfff;
rom[63268] = 12'hfff;
rom[63269] = 12'hfff;
rom[63270] = 12'hfff;
rom[63271] = 12'hfff;
rom[63272] = 12'hfff;
rom[63273] = 12'hfff;
rom[63274] = 12'hfff;
rom[63275] = 12'hfff;
rom[63276] = 12'hfff;
rom[63277] = 12'hfff;
rom[63278] = 12'hfff;
rom[63279] = 12'hfff;
rom[63280] = 12'hfff;
rom[63281] = 12'hfff;
rom[63282] = 12'hfff;
rom[63283] = 12'hfff;
rom[63284] = 12'hfff;
rom[63285] = 12'hfff;
rom[63286] = 12'hfff;
rom[63287] = 12'hfff;
rom[63288] = 12'hfff;
rom[63289] = 12'hfff;
rom[63290] = 12'hfff;
rom[63291] = 12'hfff;
rom[63292] = 12'hfff;
rom[63293] = 12'hfff;
rom[63294] = 12'hfff;
rom[63295] = 12'hfff;
rom[63296] = 12'hfff;
rom[63297] = 12'hfff;
rom[63298] = 12'hfff;
rom[63299] = 12'hfff;
rom[63300] = 12'hfff;
rom[63301] = 12'hfff;
rom[63302] = 12'hfff;
rom[63303] = 12'hfff;
rom[63304] = 12'hfff;
rom[63305] = 12'hfff;
rom[63306] = 12'hfff;
rom[63307] = 12'hfff;
rom[63308] = 12'hfff;
rom[63309] = 12'hfff;
rom[63310] = 12'hfff;
rom[63311] = 12'heee;
rom[63312] = 12'heee;
rom[63313] = 12'heee;
rom[63314] = 12'heee;
rom[63315] = 12'hddd;
rom[63316] = 12'hddd;
rom[63317] = 12'hddd;
rom[63318] = 12'hddd;
rom[63319] = 12'hccc;
rom[63320] = 12'hccc;
rom[63321] = 12'hccc;
rom[63322] = 12'hccc;
rom[63323] = 12'hccc;
rom[63324] = 12'hbbb;
rom[63325] = 12'hbbb;
rom[63326] = 12'hbbb;
rom[63327] = 12'hbbb;
rom[63328] = 12'h999;
rom[63329] = 12'h999;
rom[63330] = 12'h999;
rom[63331] = 12'h999;
rom[63332] = 12'h999;
rom[63333] = 12'h888;
rom[63334] = 12'h888;
rom[63335] = 12'h888;
rom[63336] = 12'h888;
rom[63337] = 12'h888;
rom[63338] = 12'h888;
rom[63339] = 12'h777;
rom[63340] = 12'h777;
rom[63341] = 12'h777;
rom[63342] = 12'h666;
rom[63343] = 12'h666;
rom[63344] = 12'h666;
rom[63345] = 12'h666;
rom[63346] = 12'h666;
rom[63347] = 12'h666;
rom[63348] = 12'h666;
rom[63349] = 12'h666;
rom[63350] = 12'h666;
rom[63351] = 12'h555;
rom[63352] = 12'h555;
rom[63353] = 12'h555;
rom[63354] = 12'h555;
rom[63355] = 12'h555;
rom[63356] = 12'h444;
rom[63357] = 12'h444;
rom[63358] = 12'h444;
rom[63359] = 12'h333;
rom[63360] = 12'h333;
rom[63361] = 12'h333;
rom[63362] = 12'h333;
rom[63363] = 12'h222;
rom[63364] = 12'h222;
rom[63365] = 12'h222;
rom[63366] = 12'h222;
rom[63367] = 12'h222;
rom[63368] = 12'h111;
rom[63369] = 12'h111;
rom[63370] = 12'h111;
rom[63371] = 12'h111;
rom[63372] = 12'h111;
rom[63373] = 12'h  0;
rom[63374] = 12'h  0;
rom[63375] = 12'h  0;
rom[63376] = 12'h111;
rom[63377] = 12'h111;
rom[63378] = 12'h  0;
rom[63379] = 12'h  0;
rom[63380] = 12'h  0;
rom[63381] = 12'h  0;
rom[63382] = 12'h  0;
rom[63383] = 12'h  0;
rom[63384] = 12'h  0;
rom[63385] = 12'h  0;
rom[63386] = 12'h  0;
rom[63387] = 12'h  0;
rom[63388] = 12'h  0;
rom[63389] = 12'h  0;
rom[63390] = 12'h  0;
rom[63391] = 12'h  0;
rom[63392] = 12'h  0;
rom[63393] = 12'h  0;
rom[63394] = 12'h  0;
rom[63395] = 12'h  0;
rom[63396] = 12'h  0;
rom[63397] = 12'h  0;
rom[63398] = 12'h  0;
rom[63399] = 12'h  0;
rom[63400] = 12'h  0;
rom[63401] = 12'h  0;
rom[63402] = 12'h  0;
rom[63403] = 12'h  0;
rom[63404] = 12'h  0;
rom[63405] = 12'h  0;
rom[63406] = 12'h  0;
rom[63407] = 12'h  0;
rom[63408] = 12'h111;
rom[63409] = 12'h  0;
rom[63410] = 12'h111;
rom[63411] = 12'h111;
rom[63412] = 12'h222;
rom[63413] = 12'h111;
rom[63414] = 12'h111;
rom[63415] = 12'h111;
rom[63416] = 12'h111;
rom[63417] = 12'h111;
rom[63418] = 12'h111;
rom[63419] = 12'h  0;
rom[63420] = 12'h  0;
rom[63421] = 12'h  0;
rom[63422] = 12'h  0;
rom[63423] = 12'h  0;
rom[63424] = 12'h  0;
rom[63425] = 12'h  0;
rom[63426] = 12'h  0;
rom[63427] = 12'h  0;
rom[63428] = 12'h  0;
rom[63429] = 12'h  0;
rom[63430] = 12'h  0;
rom[63431] = 12'h  0;
rom[63432] = 12'h  0;
rom[63433] = 12'h  0;
rom[63434] = 12'h  0;
rom[63435] = 12'h  0;
rom[63436] = 12'h  0;
rom[63437] = 12'h  0;
rom[63438] = 12'h  0;
rom[63439] = 12'h  0;
rom[63440] = 12'h  0;
rom[63441] = 12'h  0;
rom[63442] = 12'h  0;
rom[63443] = 12'h  0;
rom[63444] = 12'h  0;
rom[63445] = 12'h  0;
rom[63446] = 12'h  0;
rom[63447] = 12'h  0;
rom[63448] = 12'h  0;
rom[63449] = 12'h  0;
rom[63450] = 12'h  0;
rom[63451] = 12'h  0;
rom[63452] = 12'h  0;
rom[63453] = 12'h  0;
rom[63454] = 12'h  0;
rom[63455] = 12'h  0;
rom[63456] = 12'h  0;
rom[63457] = 12'h  0;
rom[63458] = 12'h  0;
rom[63459] = 12'h  0;
rom[63460] = 12'h  0;
rom[63461] = 12'h  0;
rom[63462] = 12'h  0;
rom[63463] = 12'h  0;
rom[63464] = 12'h  0;
rom[63465] = 12'h  0;
rom[63466] = 12'h  0;
rom[63467] = 12'h  0;
rom[63468] = 12'h  0;
rom[63469] = 12'h  0;
rom[63470] = 12'h  0;
rom[63471] = 12'h  0;
rom[63472] = 12'h  0;
rom[63473] = 12'h111;
rom[63474] = 12'h111;
rom[63475] = 12'h222;
rom[63476] = 12'h222;
rom[63477] = 12'h333;
rom[63478] = 12'h444;
rom[63479] = 12'h444;
rom[63480] = 12'h555;
rom[63481] = 12'h555;
rom[63482] = 12'h444;
rom[63483] = 12'h333;
rom[63484] = 12'h222;
rom[63485] = 12'h222;
rom[63486] = 12'h111;
rom[63487] = 12'h111;
rom[63488] = 12'h111;
rom[63489] = 12'h111;
rom[63490] = 12'h111;
rom[63491] = 12'h111;
rom[63492] = 12'h111;
rom[63493] = 12'h111;
rom[63494] = 12'h111;
rom[63495] = 12'h111;
rom[63496] = 12'h111;
rom[63497] = 12'h222;
rom[63498] = 12'h444;
rom[63499] = 12'h444;
rom[63500] = 12'h444;
rom[63501] = 12'h444;
rom[63502] = 12'h444;
rom[63503] = 12'h444;
rom[63504] = 12'h333;
rom[63505] = 12'h333;
rom[63506] = 12'h444;
rom[63507] = 12'h444;
rom[63508] = 12'h444;
rom[63509] = 12'h555;
rom[63510] = 12'h555;
rom[63511] = 12'h555;
rom[63512] = 12'h666;
rom[63513] = 12'h777;
rom[63514] = 12'h777;
rom[63515] = 12'h777;
rom[63516] = 12'h777;
rom[63517] = 12'h777;
rom[63518] = 12'h777;
rom[63519] = 12'h777;
rom[63520] = 12'h777;
rom[63521] = 12'h777;
rom[63522] = 12'h777;
rom[63523] = 12'h777;
rom[63524] = 12'h777;
rom[63525] = 12'h888;
rom[63526] = 12'h888;
rom[63527] = 12'h888;
rom[63528] = 12'h888;
rom[63529] = 12'h888;
rom[63530] = 12'h888;
rom[63531] = 12'h999;
rom[63532] = 12'h999;
rom[63533] = 12'h999;
rom[63534] = 12'h999;
rom[63535] = 12'h999;
rom[63536] = 12'haaa;
rom[63537] = 12'haaa;
rom[63538] = 12'haaa;
rom[63539] = 12'haaa;
rom[63540] = 12'hbbb;
rom[63541] = 12'hbbb;
rom[63542] = 12'hbbb;
rom[63543] = 12'hbbb;
rom[63544] = 12'hccc;
rom[63545] = 12'hccc;
rom[63546] = 12'hddd;
rom[63547] = 12'hddd;
rom[63548] = 12'heee;
rom[63549] = 12'heee;
rom[63550] = 12'hfff;
rom[63551] = 12'hfff;
rom[63552] = 12'hfff;
rom[63553] = 12'hfff;
rom[63554] = 12'hfff;
rom[63555] = 12'heee;
rom[63556] = 12'hddd;
rom[63557] = 12'hddd;
rom[63558] = 12'hccc;
rom[63559] = 12'hccc;
rom[63560] = 12'hccc;
rom[63561] = 12'hccc;
rom[63562] = 12'hbbb;
rom[63563] = 12'hbbb;
rom[63564] = 12'hbbb;
rom[63565] = 12'hbbb;
rom[63566] = 12'hbbb;
rom[63567] = 12'hbbb;
rom[63568] = 12'hbbb;
rom[63569] = 12'hbbb;
rom[63570] = 12'hbbb;
rom[63571] = 12'hbbb;
rom[63572] = 12'hbbb;
rom[63573] = 12'hbbb;
rom[63574] = 12'hbbb;
rom[63575] = 12'hbbb;
rom[63576] = 12'hbbb;
rom[63577] = 12'haaa;
rom[63578] = 12'h999;
rom[63579] = 12'h999;
rom[63580] = 12'h888;
rom[63581] = 12'h888;
rom[63582] = 12'h888;
rom[63583] = 12'h777;
rom[63584] = 12'h777;
rom[63585] = 12'h777;
rom[63586] = 12'h777;
rom[63587] = 12'h777;
rom[63588] = 12'h777;
rom[63589] = 12'h666;
rom[63590] = 12'h666;
rom[63591] = 12'h666;
rom[63592] = 12'h777;
rom[63593] = 12'h777;
rom[63594] = 12'h777;
rom[63595] = 12'h777;
rom[63596] = 12'h777;
rom[63597] = 12'h777;
rom[63598] = 12'h777;
rom[63599] = 12'h777;
rom[63600] = 12'hfff;
rom[63601] = 12'hfff;
rom[63602] = 12'hfff;
rom[63603] = 12'hfff;
rom[63604] = 12'hfff;
rom[63605] = 12'hfff;
rom[63606] = 12'hfff;
rom[63607] = 12'hfff;
rom[63608] = 12'hfff;
rom[63609] = 12'hfff;
rom[63610] = 12'hfff;
rom[63611] = 12'hfff;
rom[63612] = 12'hfff;
rom[63613] = 12'hfff;
rom[63614] = 12'hfff;
rom[63615] = 12'hfff;
rom[63616] = 12'hfff;
rom[63617] = 12'hfff;
rom[63618] = 12'hfff;
rom[63619] = 12'hfff;
rom[63620] = 12'hfff;
rom[63621] = 12'hfff;
rom[63622] = 12'hfff;
rom[63623] = 12'hfff;
rom[63624] = 12'hfff;
rom[63625] = 12'hfff;
rom[63626] = 12'hfff;
rom[63627] = 12'hfff;
rom[63628] = 12'hfff;
rom[63629] = 12'hfff;
rom[63630] = 12'hfff;
rom[63631] = 12'hfff;
rom[63632] = 12'hfff;
rom[63633] = 12'hfff;
rom[63634] = 12'hfff;
rom[63635] = 12'hfff;
rom[63636] = 12'hfff;
rom[63637] = 12'hfff;
rom[63638] = 12'hfff;
rom[63639] = 12'hfff;
rom[63640] = 12'hfff;
rom[63641] = 12'hfff;
rom[63642] = 12'hfff;
rom[63643] = 12'hfff;
rom[63644] = 12'hfff;
rom[63645] = 12'hfff;
rom[63646] = 12'hfff;
rom[63647] = 12'hfff;
rom[63648] = 12'hfff;
rom[63649] = 12'hfff;
rom[63650] = 12'hfff;
rom[63651] = 12'hfff;
rom[63652] = 12'hfff;
rom[63653] = 12'hfff;
rom[63654] = 12'hfff;
rom[63655] = 12'hfff;
rom[63656] = 12'hfff;
rom[63657] = 12'hfff;
rom[63658] = 12'hfff;
rom[63659] = 12'hfff;
rom[63660] = 12'hfff;
rom[63661] = 12'hfff;
rom[63662] = 12'hfff;
rom[63663] = 12'hfff;
rom[63664] = 12'hfff;
rom[63665] = 12'hfff;
rom[63666] = 12'hfff;
rom[63667] = 12'hfff;
rom[63668] = 12'hfff;
rom[63669] = 12'hfff;
rom[63670] = 12'hfff;
rom[63671] = 12'hfff;
rom[63672] = 12'hfff;
rom[63673] = 12'hfff;
rom[63674] = 12'hfff;
rom[63675] = 12'hfff;
rom[63676] = 12'hfff;
rom[63677] = 12'hfff;
rom[63678] = 12'hfff;
rom[63679] = 12'hfff;
rom[63680] = 12'hfff;
rom[63681] = 12'hfff;
rom[63682] = 12'hfff;
rom[63683] = 12'hfff;
rom[63684] = 12'hfff;
rom[63685] = 12'hfff;
rom[63686] = 12'hfff;
rom[63687] = 12'hfff;
rom[63688] = 12'hfff;
rom[63689] = 12'hfff;
rom[63690] = 12'hfff;
rom[63691] = 12'hfff;
rom[63692] = 12'hfff;
rom[63693] = 12'hfff;
rom[63694] = 12'hfff;
rom[63695] = 12'hfff;
rom[63696] = 12'hfff;
rom[63697] = 12'hfff;
rom[63698] = 12'hfff;
rom[63699] = 12'hfff;
rom[63700] = 12'hfff;
rom[63701] = 12'hfff;
rom[63702] = 12'hfff;
rom[63703] = 12'hfff;
rom[63704] = 12'hfff;
rom[63705] = 12'hfff;
rom[63706] = 12'hfff;
rom[63707] = 12'hfff;
rom[63708] = 12'hfff;
rom[63709] = 12'hfff;
rom[63710] = 12'hfff;
rom[63711] = 12'hfff;
rom[63712] = 12'hfff;
rom[63713] = 12'heee;
rom[63714] = 12'hddd;
rom[63715] = 12'hddd;
rom[63716] = 12'hccc;
rom[63717] = 12'hccc;
rom[63718] = 12'hccc;
rom[63719] = 12'hccc;
rom[63720] = 12'hccc;
rom[63721] = 12'hbbb;
rom[63722] = 12'hbbb;
rom[63723] = 12'hbbb;
rom[63724] = 12'hbbb;
rom[63725] = 12'hbbb;
rom[63726] = 12'hbbb;
rom[63727] = 12'hbbb;
rom[63728] = 12'haaa;
rom[63729] = 12'haaa;
rom[63730] = 12'haaa;
rom[63731] = 12'h999;
rom[63732] = 12'h999;
rom[63733] = 12'h999;
rom[63734] = 12'h999;
rom[63735] = 12'h888;
rom[63736] = 12'h888;
rom[63737] = 12'h888;
rom[63738] = 12'h888;
rom[63739] = 12'h888;
rom[63740] = 12'h888;
rom[63741] = 12'h777;
rom[63742] = 12'h777;
rom[63743] = 12'h666;
rom[63744] = 12'h666;
rom[63745] = 12'h666;
rom[63746] = 12'h666;
rom[63747] = 12'h666;
rom[63748] = 12'h555;
rom[63749] = 12'h555;
rom[63750] = 12'h555;
rom[63751] = 12'h444;
rom[63752] = 12'h444;
rom[63753] = 12'h444;
rom[63754] = 12'h444;
rom[63755] = 12'h444;
rom[63756] = 12'h444;
rom[63757] = 12'h444;
rom[63758] = 12'h444;
rom[63759] = 12'h333;
rom[63760] = 12'h333;
rom[63761] = 12'h333;
rom[63762] = 12'h333;
rom[63763] = 12'h222;
rom[63764] = 12'h222;
rom[63765] = 12'h222;
rom[63766] = 12'h222;
rom[63767] = 12'h222;
rom[63768] = 12'h111;
rom[63769] = 12'h111;
rom[63770] = 12'h111;
rom[63771] = 12'h111;
rom[63772] = 12'h111;
rom[63773] = 12'h  0;
rom[63774] = 12'h  0;
rom[63775] = 12'h  0;
rom[63776] = 12'h111;
rom[63777] = 12'h111;
rom[63778] = 12'h  0;
rom[63779] = 12'h  0;
rom[63780] = 12'h  0;
rom[63781] = 12'h  0;
rom[63782] = 12'h  0;
rom[63783] = 12'h  0;
rom[63784] = 12'h  0;
rom[63785] = 12'h  0;
rom[63786] = 12'h  0;
rom[63787] = 12'h  0;
rom[63788] = 12'h  0;
rom[63789] = 12'h  0;
rom[63790] = 12'h  0;
rom[63791] = 12'h  0;
rom[63792] = 12'h  0;
rom[63793] = 12'h  0;
rom[63794] = 12'h  0;
rom[63795] = 12'h  0;
rom[63796] = 12'h  0;
rom[63797] = 12'h  0;
rom[63798] = 12'h  0;
rom[63799] = 12'h  0;
rom[63800] = 12'h  0;
rom[63801] = 12'h  0;
rom[63802] = 12'h  0;
rom[63803] = 12'h  0;
rom[63804] = 12'h  0;
rom[63805] = 12'h  0;
rom[63806] = 12'h  0;
rom[63807] = 12'h  0;
rom[63808] = 12'h111;
rom[63809] = 12'h  0;
rom[63810] = 12'h111;
rom[63811] = 12'h111;
rom[63812] = 12'h222;
rom[63813] = 12'h111;
rom[63814] = 12'h111;
rom[63815] = 12'h111;
rom[63816] = 12'h111;
rom[63817] = 12'h111;
rom[63818] = 12'h111;
rom[63819] = 12'h  0;
rom[63820] = 12'h  0;
rom[63821] = 12'h  0;
rom[63822] = 12'h  0;
rom[63823] = 12'h  0;
rom[63824] = 12'h  0;
rom[63825] = 12'h  0;
rom[63826] = 12'h  0;
rom[63827] = 12'h  0;
rom[63828] = 12'h  0;
rom[63829] = 12'h  0;
rom[63830] = 12'h  0;
rom[63831] = 12'h  0;
rom[63832] = 12'h  0;
rom[63833] = 12'h  0;
rom[63834] = 12'h  0;
rom[63835] = 12'h  0;
rom[63836] = 12'h  0;
rom[63837] = 12'h  0;
rom[63838] = 12'h  0;
rom[63839] = 12'h  0;
rom[63840] = 12'h  0;
rom[63841] = 12'h  0;
rom[63842] = 12'h  0;
rom[63843] = 12'h  0;
rom[63844] = 12'h  0;
rom[63845] = 12'h  0;
rom[63846] = 12'h  0;
rom[63847] = 12'h  0;
rom[63848] = 12'h  0;
rom[63849] = 12'h  0;
rom[63850] = 12'h  0;
rom[63851] = 12'h  0;
rom[63852] = 12'h  0;
rom[63853] = 12'h  0;
rom[63854] = 12'h  0;
rom[63855] = 12'h  0;
rom[63856] = 12'h  0;
rom[63857] = 12'h  0;
rom[63858] = 12'h  0;
rom[63859] = 12'h  0;
rom[63860] = 12'h  0;
rom[63861] = 12'h  0;
rom[63862] = 12'h  0;
rom[63863] = 12'h  0;
rom[63864] = 12'h  0;
rom[63865] = 12'h  0;
rom[63866] = 12'h  0;
rom[63867] = 12'h  0;
rom[63868] = 12'h  0;
rom[63869] = 12'h  0;
rom[63870] = 12'h  0;
rom[63871] = 12'h  0;
rom[63872] = 12'h111;
rom[63873] = 12'h111;
rom[63874] = 12'h111;
rom[63875] = 12'h222;
rom[63876] = 12'h222;
rom[63877] = 12'h333;
rom[63878] = 12'h444;
rom[63879] = 12'h555;
rom[63880] = 12'h555;
rom[63881] = 12'h555;
rom[63882] = 12'h444;
rom[63883] = 12'h333;
rom[63884] = 12'h222;
rom[63885] = 12'h222;
rom[63886] = 12'h111;
rom[63887] = 12'h111;
rom[63888] = 12'h111;
rom[63889] = 12'h111;
rom[63890] = 12'h111;
rom[63891] = 12'h111;
rom[63892] = 12'h111;
rom[63893] = 12'h111;
rom[63894] = 12'h111;
rom[63895] = 12'h111;
rom[63896] = 12'h111;
rom[63897] = 12'h222;
rom[63898] = 12'h333;
rom[63899] = 12'h444;
rom[63900] = 12'h444;
rom[63901] = 12'h444;
rom[63902] = 12'h444;
rom[63903] = 12'h444;
rom[63904] = 12'h333;
rom[63905] = 12'h333;
rom[63906] = 12'h333;
rom[63907] = 12'h444;
rom[63908] = 12'h444;
rom[63909] = 12'h555;
rom[63910] = 12'h555;
rom[63911] = 12'h555;
rom[63912] = 12'h666;
rom[63913] = 12'h777;
rom[63914] = 12'h777;
rom[63915] = 12'h888;
rom[63916] = 12'h888;
rom[63917] = 12'h777;
rom[63918] = 12'h777;
rom[63919] = 12'h777;
rom[63920] = 12'h777;
rom[63921] = 12'h777;
rom[63922] = 12'h777;
rom[63923] = 12'h777;
rom[63924] = 12'h888;
rom[63925] = 12'h888;
rom[63926] = 12'h888;
rom[63927] = 12'h888;
rom[63928] = 12'h888;
rom[63929] = 12'h888;
rom[63930] = 12'h999;
rom[63931] = 12'h999;
rom[63932] = 12'h999;
rom[63933] = 12'h999;
rom[63934] = 12'haaa;
rom[63935] = 12'haaa;
rom[63936] = 12'haaa;
rom[63937] = 12'haaa;
rom[63938] = 12'haaa;
rom[63939] = 12'hbbb;
rom[63940] = 12'hbbb;
rom[63941] = 12'hbbb;
rom[63942] = 12'hbbb;
rom[63943] = 12'hccc;
rom[63944] = 12'hccc;
rom[63945] = 12'hccc;
rom[63946] = 12'hddd;
rom[63947] = 12'heee;
rom[63948] = 12'heee;
rom[63949] = 12'hfff;
rom[63950] = 12'hfff;
rom[63951] = 12'hfff;
rom[63952] = 12'hfff;
rom[63953] = 12'hfff;
rom[63954] = 12'heee;
rom[63955] = 12'heee;
rom[63956] = 12'hddd;
rom[63957] = 12'hddd;
rom[63958] = 12'hccc;
rom[63959] = 12'hccc;
rom[63960] = 12'hccc;
rom[63961] = 12'hccc;
rom[63962] = 12'hbbb;
rom[63963] = 12'hbbb;
rom[63964] = 12'hbbb;
rom[63965] = 12'hbbb;
rom[63966] = 12'hbbb;
rom[63967] = 12'hbbb;
rom[63968] = 12'hbbb;
rom[63969] = 12'hbbb;
rom[63970] = 12'hbbb;
rom[63971] = 12'hbbb;
rom[63972] = 12'hbbb;
rom[63973] = 12'hccc;
rom[63974] = 12'hbbb;
rom[63975] = 12'hbbb;
rom[63976] = 12'hbbb;
rom[63977] = 12'haaa;
rom[63978] = 12'haaa;
rom[63979] = 12'h999;
rom[63980] = 12'h888;
rom[63981] = 12'h888;
rom[63982] = 12'h888;
rom[63983] = 12'h888;
rom[63984] = 12'h777;
rom[63985] = 12'h777;
rom[63986] = 12'h777;
rom[63987] = 12'h777;
rom[63988] = 12'h666;
rom[63989] = 12'h666;
rom[63990] = 12'h666;
rom[63991] = 12'h666;
rom[63992] = 12'h666;
rom[63993] = 12'h666;
rom[63994] = 12'h666;
rom[63995] = 12'h666;
rom[63996] = 12'h666;
rom[63997] = 12'h666;
rom[63998] = 12'h666;
rom[63999] = 12'h666;
rom[64000] = 12'hfff;
rom[64001] = 12'hfff;
rom[64002] = 12'hfff;
rom[64003] = 12'hfff;
rom[64004] = 12'hfff;
rom[64005] = 12'hfff;
rom[64006] = 12'hfff;
rom[64007] = 12'hfff;
rom[64008] = 12'hfff;
rom[64009] = 12'hfff;
rom[64010] = 12'hfff;
rom[64011] = 12'hfff;
rom[64012] = 12'hfff;
rom[64013] = 12'hfff;
rom[64014] = 12'hfff;
rom[64015] = 12'hfff;
rom[64016] = 12'hfff;
rom[64017] = 12'hfff;
rom[64018] = 12'hfff;
rom[64019] = 12'hfff;
rom[64020] = 12'hfff;
rom[64021] = 12'hfff;
rom[64022] = 12'hfff;
rom[64023] = 12'hfff;
rom[64024] = 12'hfff;
rom[64025] = 12'hfff;
rom[64026] = 12'hfff;
rom[64027] = 12'hfff;
rom[64028] = 12'hfff;
rom[64029] = 12'hfff;
rom[64030] = 12'hfff;
rom[64031] = 12'hfff;
rom[64032] = 12'hfff;
rom[64033] = 12'hfff;
rom[64034] = 12'hfff;
rom[64035] = 12'hfff;
rom[64036] = 12'hfff;
rom[64037] = 12'hfff;
rom[64038] = 12'hfff;
rom[64039] = 12'hfff;
rom[64040] = 12'hfff;
rom[64041] = 12'hfff;
rom[64042] = 12'hfff;
rom[64043] = 12'hfff;
rom[64044] = 12'hfff;
rom[64045] = 12'hfff;
rom[64046] = 12'hfff;
rom[64047] = 12'hfff;
rom[64048] = 12'hfff;
rom[64049] = 12'hfff;
rom[64050] = 12'hfff;
rom[64051] = 12'hfff;
rom[64052] = 12'hfff;
rom[64053] = 12'hfff;
rom[64054] = 12'hfff;
rom[64055] = 12'hfff;
rom[64056] = 12'hfff;
rom[64057] = 12'hfff;
rom[64058] = 12'hfff;
rom[64059] = 12'hfff;
rom[64060] = 12'hfff;
rom[64061] = 12'hfff;
rom[64062] = 12'hfff;
rom[64063] = 12'hfff;
rom[64064] = 12'hfff;
rom[64065] = 12'hfff;
rom[64066] = 12'hfff;
rom[64067] = 12'hfff;
rom[64068] = 12'hfff;
rom[64069] = 12'hfff;
rom[64070] = 12'hfff;
rom[64071] = 12'hfff;
rom[64072] = 12'hfff;
rom[64073] = 12'hfff;
rom[64074] = 12'hfff;
rom[64075] = 12'hfff;
rom[64076] = 12'hfff;
rom[64077] = 12'hfff;
rom[64078] = 12'hfff;
rom[64079] = 12'hfff;
rom[64080] = 12'hfff;
rom[64081] = 12'hfff;
rom[64082] = 12'hfff;
rom[64083] = 12'hfff;
rom[64084] = 12'hfff;
rom[64085] = 12'hfff;
rom[64086] = 12'hfff;
rom[64087] = 12'hfff;
rom[64088] = 12'hfff;
rom[64089] = 12'hfff;
rom[64090] = 12'hfff;
rom[64091] = 12'hfff;
rom[64092] = 12'hfff;
rom[64093] = 12'hfff;
rom[64094] = 12'hfff;
rom[64095] = 12'hfff;
rom[64096] = 12'hfff;
rom[64097] = 12'hfff;
rom[64098] = 12'hfff;
rom[64099] = 12'hfff;
rom[64100] = 12'hfff;
rom[64101] = 12'hfff;
rom[64102] = 12'hfff;
rom[64103] = 12'hfff;
rom[64104] = 12'hfff;
rom[64105] = 12'hfff;
rom[64106] = 12'hfff;
rom[64107] = 12'hfff;
rom[64108] = 12'hfff;
rom[64109] = 12'hfff;
rom[64110] = 12'hfff;
rom[64111] = 12'heee;
rom[64112] = 12'heee;
rom[64113] = 12'heee;
rom[64114] = 12'heee;
rom[64115] = 12'heee;
rom[64116] = 12'hddd;
rom[64117] = 12'hddd;
rom[64118] = 12'hccc;
rom[64119] = 12'hccc;
rom[64120] = 12'hbbb;
rom[64121] = 12'hbbb;
rom[64122] = 12'hbbb;
rom[64123] = 12'haaa;
rom[64124] = 12'haaa;
rom[64125] = 12'haaa;
rom[64126] = 12'haaa;
rom[64127] = 12'haaa;
rom[64128] = 12'haaa;
rom[64129] = 12'haaa;
rom[64130] = 12'h999;
rom[64131] = 12'h999;
rom[64132] = 12'h999;
rom[64133] = 12'h999;
rom[64134] = 12'h888;
rom[64135] = 12'h888;
rom[64136] = 12'h888;
rom[64137] = 12'h888;
rom[64138] = 12'h888;
rom[64139] = 12'h888;
rom[64140] = 12'h777;
rom[64141] = 12'h777;
rom[64142] = 12'h666;
rom[64143] = 12'h666;
rom[64144] = 12'h666;
rom[64145] = 12'h666;
rom[64146] = 12'h666;
rom[64147] = 12'h555;
rom[64148] = 12'h555;
rom[64149] = 12'h555;
rom[64150] = 12'h444;
rom[64151] = 12'h444;
rom[64152] = 12'h444;
rom[64153] = 12'h333;
rom[64154] = 12'h333;
rom[64155] = 12'h333;
rom[64156] = 12'h333;
rom[64157] = 12'h333;
rom[64158] = 12'h333;
rom[64159] = 12'h333;
rom[64160] = 12'h222;
rom[64161] = 12'h222;
rom[64162] = 12'h222;
rom[64163] = 12'h222;
rom[64164] = 12'h222;
rom[64165] = 12'h222;
rom[64166] = 12'h111;
rom[64167] = 12'h111;
rom[64168] = 12'h111;
rom[64169] = 12'h111;
rom[64170] = 12'h111;
rom[64171] = 12'h111;
rom[64172] = 12'h111;
rom[64173] = 12'h111;
rom[64174] = 12'h111;
rom[64175] = 12'h  0;
rom[64176] = 12'h111;
rom[64177] = 12'h111;
rom[64178] = 12'h  0;
rom[64179] = 12'h  0;
rom[64180] = 12'h  0;
rom[64181] = 12'h  0;
rom[64182] = 12'h  0;
rom[64183] = 12'h  0;
rom[64184] = 12'h111;
rom[64185] = 12'h  0;
rom[64186] = 12'h  0;
rom[64187] = 12'h  0;
rom[64188] = 12'h  0;
rom[64189] = 12'h111;
rom[64190] = 12'h  0;
rom[64191] = 12'h  0;
rom[64192] = 12'h  0;
rom[64193] = 12'h  0;
rom[64194] = 12'h  0;
rom[64195] = 12'h  0;
rom[64196] = 12'h  0;
rom[64197] = 12'h  0;
rom[64198] = 12'h  0;
rom[64199] = 12'h  0;
rom[64200] = 12'h  0;
rom[64201] = 12'h  0;
rom[64202] = 12'h  0;
rom[64203] = 12'h  0;
rom[64204] = 12'h  0;
rom[64205] = 12'h  0;
rom[64206] = 12'h  0;
rom[64207] = 12'h  0;
rom[64208] = 12'h  0;
rom[64209] = 12'h111;
rom[64210] = 12'h111;
rom[64211] = 12'h111;
rom[64212] = 12'h111;
rom[64213] = 12'h111;
rom[64214] = 12'h111;
rom[64215] = 12'h111;
rom[64216] = 12'h111;
rom[64217] = 12'h111;
rom[64218] = 12'h  0;
rom[64219] = 12'h  0;
rom[64220] = 12'h  0;
rom[64221] = 12'h  0;
rom[64222] = 12'h  0;
rom[64223] = 12'h  0;
rom[64224] = 12'h  0;
rom[64225] = 12'h  0;
rom[64226] = 12'h  0;
rom[64227] = 12'h  0;
rom[64228] = 12'h  0;
rom[64229] = 12'h  0;
rom[64230] = 12'h  0;
rom[64231] = 12'h  0;
rom[64232] = 12'h  0;
rom[64233] = 12'h  0;
rom[64234] = 12'h  0;
rom[64235] = 12'h  0;
rom[64236] = 12'h  0;
rom[64237] = 12'h  0;
rom[64238] = 12'h  0;
rom[64239] = 12'h  0;
rom[64240] = 12'h  0;
rom[64241] = 12'h  0;
rom[64242] = 12'h  0;
rom[64243] = 12'h  0;
rom[64244] = 12'h  0;
rom[64245] = 12'h  0;
rom[64246] = 12'h  0;
rom[64247] = 12'h  0;
rom[64248] = 12'h  0;
rom[64249] = 12'h  0;
rom[64250] = 12'h  0;
rom[64251] = 12'h  0;
rom[64252] = 12'h  0;
rom[64253] = 12'h  0;
rom[64254] = 12'h  0;
rom[64255] = 12'h  0;
rom[64256] = 12'h  0;
rom[64257] = 12'h  0;
rom[64258] = 12'h  0;
rom[64259] = 12'h  0;
rom[64260] = 12'h  0;
rom[64261] = 12'h  0;
rom[64262] = 12'h  0;
rom[64263] = 12'h  0;
rom[64264] = 12'h  0;
rom[64265] = 12'h  0;
rom[64266] = 12'h  0;
rom[64267] = 12'h  0;
rom[64268] = 12'h  0;
rom[64269] = 12'h  0;
rom[64270] = 12'h  0;
rom[64271] = 12'h  0;
rom[64272] = 12'h111;
rom[64273] = 12'h111;
rom[64274] = 12'h111;
rom[64275] = 12'h222;
rom[64276] = 12'h222;
rom[64277] = 12'h333;
rom[64278] = 12'h444;
rom[64279] = 12'h555;
rom[64280] = 12'h444;
rom[64281] = 12'h444;
rom[64282] = 12'h444;
rom[64283] = 12'h444;
rom[64284] = 12'h222;
rom[64285] = 12'h111;
rom[64286] = 12'h111;
rom[64287] = 12'h111;
rom[64288] = 12'h111;
rom[64289] = 12'h111;
rom[64290] = 12'h111;
rom[64291] = 12'h111;
rom[64292] = 12'h111;
rom[64293] = 12'h111;
rom[64294] = 12'h111;
rom[64295] = 12'h111;
rom[64296] = 12'h222;
rom[64297] = 12'h222;
rom[64298] = 12'h333;
rom[64299] = 12'h444;
rom[64300] = 12'h444;
rom[64301] = 12'h444;
rom[64302] = 12'h444;
rom[64303] = 12'h444;
rom[64304] = 12'h333;
rom[64305] = 12'h444;
rom[64306] = 12'h444;
rom[64307] = 12'h444;
rom[64308] = 12'h444;
rom[64309] = 12'h444;
rom[64310] = 12'h555;
rom[64311] = 12'h555;
rom[64312] = 12'h666;
rom[64313] = 12'h666;
rom[64314] = 12'h777;
rom[64315] = 12'h888;
rom[64316] = 12'h888;
rom[64317] = 12'h888;
rom[64318] = 12'h777;
rom[64319] = 12'h777;
rom[64320] = 12'h777;
rom[64321] = 12'h777;
rom[64322] = 12'h888;
rom[64323] = 12'h888;
rom[64324] = 12'h888;
rom[64325] = 12'h888;
rom[64326] = 12'h888;
rom[64327] = 12'h888;
rom[64328] = 12'h999;
rom[64329] = 12'h999;
rom[64330] = 12'h999;
rom[64331] = 12'h999;
rom[64332] = 12'h999;
rom[64333] = 12'haaa;
rom[64334] = 12'haaa;
rom[64335] = 12'haaa;
rom[64336] = 12'haaa;
rom[64337] = 12'haaa;
rom[64338] = 12'hbbb;
rom[64339] = 12'hbbb;
rom[64340] = 12'hbbb;
rom[64341] = 12'hbbb;
rom[64342] = 12'hccc;
rom[64343] = 12'hccc;
rom[64344] = 12'hccc;
rom[64345] = 12'hddd;
rom[64346] = 12'hddd;
rom[64347] = 12'heee;
rom[64348] = 12'hfff;
rom[64349] = 12'hfff;
rom[64350] = 12'hfff;
rom[64351] = 12'hfff;
rom[64352] = 12'hfff;
rom[64353] = 12'heee;
rom[64354] = 12'heee;
rom[64355] = 12'hddd;
rom[64356] = 12'hddd;
rom[64357] = 12'hddd;
rom[64358] = 12'hccc;
rom[64359] = 12'hccc;
rom[64360] = 12'hccc;
rom[64361] = 12'hbbb;
rom[64362] = 12'hbbb;
rom[64363] = 12'hbbb;
rom[64364] = 12'hbbb;
rom[64365] = 12'hbbb;
rom[64366] = 12'hbbb;
rom[64367] = 12'haaa;
rom[64368] = 12'haaa;
rom[64369] = 12'haaa;
rom[64370] = 12'hbbb;
rom[64371] = 12'hbbb;
rom[64372] = 12'hbbb;
rom[64373] = 12'hbbb;
rom[64374] = 12'hbbb;
rom[64375] = 12'hbbb;
rom[64376] = 12'hccc;
rom[64377] = 12'hbbb;
rom[64378] = 12'haaa;
rom[64379] = 12'h999;
rom[64380] = 12'h999;
rom[64381] = 12'h888;
rom[64382] = 12'h888;
rom[64383] = 12'h888;
rom[64384] = 12'h777;
rom[64385] = 12'h777;
rom[64386] = 12'h777;
rom[64387] = 12'h666;
rom[64388] = 12'h666;
rom[64389] = 12'h777;
rom[64390] = 12'h777;
rom[64391] = 12'h777;
rom[64392] = 12'h666;
rom[64393] = 12'h666;
rom[64394] = 12'h666;
rom[64395] = 12'h666;
rom[64396] = 12'h666;
rom[64397] = 12'h666;
rom[64398] = 12'h777;
rom[64399] = 12'h777;
rom[64400] = 12'hfff;
rom[64401] = 12'hfff;
rom[64402] = 12'hfff;
rom[64403] = 12'hfff;
rom[64404] = 12'hfff;
rom[64405] = 12'hfff;
rom[64406] = 12'hfff;
rom[64407] = 12'hfff;
rom[64408] = 12'hfff;
rom[64409] = 12'hfff;
rom[64410] = 12'hfff;
rom[64411] = 12'hfff;
rom[64412] = 12'hfff;
rom[64413] = 12'hfff;
rom[64414] = 12'hfff;
rom[64415] = 12'hfff;
rom[64416] = 12'hfff;
rom[64417] = 12'hfff;
rom[64418] = 12'hfff;
rom[64419] = 12'hfff;
rom[64420] = 12'hfff;
rom[64421] = 12'hfff;
rom[64422] = 12'hfff;
rom[64423] = 12'hfff;
rom[64424] = 12'hfff;
rom[64425] = 12'hfff;
rom[64426] = 12'hfff;
rom[64427] = 12'hfff;
rom[64428] = 12'hfff;
rom[64429] = 12'hfff;
rom[64430] = 12'hfff;
rom[64431] = 12'hfff;
rom[64432] = 12'hfff;
rom[64433] = 12'hfff;
rom[64434] = 12'hfff;
rom[64435] = 12'hfff;
rom[64436] = 12'hfff;
rom[64437] = 12'hfff;
rom[64438] = 12'hfff;
rom[64439] = 12'hfff;
rom[64440] = 12'hfff;
rom[64441] = 12'hfff;
rom[64442] = 12'hfff;
rom[64443] = 12'hfff;
rom[64444] = 12'hfff;
rom[64445] = 12'hfff;
rom[64446] = 12'hfff;
rom[64447] = 12'hfff;
rom[64448] = 12'hfff;
rom[64449] = 12'hfff;
rom[64450] = 12'hfff;
rom[64451] = 12'hfff;
rom[64452] = 12'hfff;
rom[64453] = 12'hfff;
rom[64454] = 12'hfff;
rom[64455] = 12'hfff;
rom[64456] = 12'hfff;
rom[64457] = 12'hfff;
rom[64458] = 12'hfff;
rom[64459] = 12'hfff;
rom[64460] = 12'hfff;
rom[64461] = 12'hfff;
rom[64462] = 12'hfff;
rom[64463] = 12'hfff;
rom[64464] = 12'hfff;
rom[64465] = 12'hfff;
rom[64466] = 12'hfff;
rom[64467] = 12'hfff;
rom[64468] = 12'hfff;
rom[64469] = 12'hfff;
rom[64470] = 12'hfff;
rom[64471] = 12'hfff;
rom[64472] = 12'hfff;
rom[64473] = 12'hfff;
rom[64474] = 12'hfff;
rom[64475] = 12'hfff;
rom[64476] = 12'hfff;
rom[64477] = 12'hfff;
rom[64478] = 12'hfff;
rom[64479] = 12'hfff;
rom[64480] = 12'hfff;
rom[64481] = 12'hfff;
rom[64482] = 12'hfff;
rom[64483] = 12'hfff;
rom[64484] = 12'hfff;
rom[64485] = 12'hfff;
rom[64486] = 12'hfff;
rom[64487] = 12'hfff;
rom[64488] = 12'hfff;
rom[64489] = 12'hfff;
rom[64490] = 12'hfff;
rom[64491] = 12'hfff;
rom[64492] = 12'hfff;
rom[64493] = 12'hfff;
rom[64494] = 12'hfff;
rom[64495] = 12'hfff;
rom[64496] = 12'hfff;
rom[64497] = 12'hfff;
rom[64498] = 12'hfff;
rom[64499] = 12'hfff;
rom[64500] = 12'hfff;
rom[64501] = 12'hfff;
rom[64502] = 12'hfff;
rom[64503] = 12'hfff;
rom[64504] = 12'hfff;
rom[64505] = 12'hfff;
rom[64506] = 12'hfff;
rom[64507] = 12'hfff;
rom[64508] = 12'hfff;
rom[64509] = 12'hfff;
rom[64510] = 12'hfff;
rom[64511] = 12'heee;
rom[64512] = 12'heee;
rom[64513] = 12'heee;
rom[64514] = 12'heee;
rom[64515] = 12'heee;
rom[64516] = 12'heee;
rom[64517] = 12'hddd;
rom[64518] = 12'hddd;
rom[64519] = 12'hddd;
rom[64520] = 12'hccc;
rom[64521] = 12'hccc;
rom[64522] = 12'hbbb;
rom[64523] = 12'hbbb;
rom[64524] = 12'hbbb;
rom[64525] = 12'haaa;
rom[64526] = 12'haaa;
rom[64527] = 12'haaa;
rom[64528] = 12'h999;
rom[64529] = 12'h999;
rom[64530] = 12'h999;
rom[64531] = 12'h999;
rom[64532] = 12'h888;
rom[64533] = 12'h888;
rom[64534] = 12'h888;
rom[64535] = 12'h888;
rom[64536] = 12'h777;
rom[64537] = 12'h777;
rom[64538] = 12'h777;
rom[64539] = 12'h666;
rom[64540] = 12'h666;
rom[64541] = 12'h666;
rom[64542] = 12'h666;
rom[64543] = 12'h666;
rom[64544] = 12'h777;
rom[64545] = 12'h666;
rom[64546] = 12'h666;
rom[64547] = 12'h666;
rom[64548] = 12'h555;
rom[64549] = 12'h555;
rom[64550] = 12'h444;
rom[64551] = 12'h444;
rom[64552] = 12'h444;
rom[64553] = 12'h333;
rom[64554] = 12'h333;
rom[64555] = 12'h333;
rom[64556] = 12'h333;
rom[64557] = 12'h333;
rom[64558] = 12'h333;
rom[64559] = 12'h333;
rom[64560] = 12'h222;
rom[64561] = 12'h222;
rom[64562] = 12'h222;
rom[64563] = 12'h222;
rom[64564] = 12'h222;
rom[64565] = 12'h222;
rom[64566] = 12'h111;
rom[64567] = 12'h111;
rom[64568] = 12'h111;
rom[64569] = 12'h111;
rom[64570] = 12'h111;
rom[64571] = 12'h111;
rom[64572] = 12'h111;
rom[64573] = 12'h111;
rom[64574] = 12'h111;
rom[64575] = 12'h111;
rom[64576] = 12'h111;
rom[64577] = 12'h111;
rom[64578] = 12'h  0;
rom[64579] = 12'h  0;
rom[64580] = 12'h  0;
rom[64581] = 12'h  0;
rom[64582] = 12'h  0;
rom[64583] = 12'h  0;
rom[64584] = 12'h111;
rom[64585] = 12'h  0;
rom[64586] = 12'h  0;
rom[64587] = 12'h  0;
rom[64588] = 12'h  0;
rom[64589] = 12'h111;
rom[64590] = 12'h  0;
rom[64591] = 12'h  0;
rom[64592] = 12'h  0;
rom[64593] = 12'h  0;
rom[64594] = 12'h  0;
rom[64595] = 12'h  0;
rom[64596] = 12'h  0;
rom[64597] = 12'h  0;
rom[64598] = 12'h  0;
rom[64599] = 12'h  0;
rom[64600] = 12'h  0;
rom[64601] = 12'h  0;
rom[64602] = 12'h  0;
rom[64603] = 12'h  0;
rom[64604] = 12'h  0;
rom[64605] = 12'h  0;
rom[64606] = 12'h  0;
rom[64607] = 12'h  0;
rom[64608] = 12'h  0;
rom[64609] = 12'h111;
rom[64610] = 12'h111;
rom[64611] = 12'h111;
rom[64612] = 12'h111;
rom[64613] = 12'h111;
rom[64614] = 12'h111;
rom[64615] = 12'h111;
rom[64616] = 12'h111;
rom[64617] = 12'h111;
rom[64618] = 12'h  0;
rom[64619] = 12'h  0;
rom[64620] = 12'h  0;
rom[64621] = 12'h  0;
rom[64622] = 12'h  0;
rom[64623] = 12'h  0;
rom[64624] = 12'h  0;
rom[64625] = 12'h  0;
rom[64626] = 12'h  0;
rom[64627] = 12'h  0;
rom[64628] = 12'h  0;
rom[64629] = 12'h  0;
rom[64630] = 12'h  0;
rom[64631] = 12'h  0;
rom[64632] = 12'h  0;
rom[64633] = 12'h  0;
rom[64634] = 12'h  0;
rom[64635] = 12'h  0;
rom[64636] = 12'h  0;
rom[64637] = 12'h  0;
rom[64638] = 12'h  0;
rom[64639] = 12'h  0;
rom[64640] = 12'h  0;
rom[64641] = 12'h  0;
rom[64642] = 12'h  0;
rom[64643] = 12'h  0;
rom[64644] = 12'h  0;
rom[64645] = 12'h  0;
rom[64646] = 12'h  0;
rom[64647] = 12'h  0;
rom[64648] = 12'h  0;
rom[64649] = 12'h  0;
rom[64650] = 12'h  0;
rom[64651] = 12'h  0;
rom[64652] = 12'h  0;
rom[64653] = 12'h  0;
rom[64654] = 12'h  0;
rom[64655] = 12'h  0;
rom[64656] = 12'h  0;
rom[64657] = 12'h  0;
rom[64658] = 12'h  0;
rom[64659] = 12'h  0;
rom[64660] = 12'h  0;
rom[64661] = 12'h  0;
rom[64662] = 12'h  0;
rom[64663] = 12'h  0;
rom[64664] = 12'h  0;
rom[64665] = 12'h  0;
rom[64666] = 12'h  0;
rom[64667] = 12'h  0;
rom[64668] = 12'h  0;
rom[64669] = 12'h  0;
rom[64670] = 12'h  0;
rom[64671] = 12'h  0;
rom[64672] = 12'h111;
rom[64673] = 12'h111;
rom[64674] = 12'h111;
rom[64675] = 12'h222;
rom[64676] = 12'h222;
rom[64677] = 12'h333;
rom[64678] = 12'h444;
rom[64679] = 12'h555;
rom[64680] = 12'h444;
rom[64681] = 12'h444;
rom[64682] = 12'h444;
rom[64683] = 12'h444;
rom[64684] = 12'h222;
rom[64685] = 12'h111;
rom[64686] = 12'h111;
rom[64687] = 12'h111;
rom[64688] = 12'h111;
rom[64689] = 12'h111;
rom[64690] = 12'h111;
rom[64691] = 12'h111;
rom[64692] = 12'h111;
rom[64693] = 12'h111;
rom[64694] = 12'h111;
rom[64695] = 12'h111;
rom[64696] = 12'h222;
rom[64697] = 12'h222;
rom[64698] = 12'h333;
rom[64699] = 12'h444;
rom[64700] = 12'h444;
rom[64701] = 12'h444;
rom[64702] = 12'h444;
rom[64703] = 12'h444;
rom[64704] = 12'h333;
rom[64705] = 12'h444;
rom[64706] = 12'h444;
rom[64707] = 12'h444;
rom[64708] = 12'h444;
rom[64709] = 12'h444;
rom[64710] = 12'h555;
rom[64711] = 12'h555;
rom[64712] = 12'h666;
rom[64713] = 12'h666;
rom[64714] = 12'h777;
rom[64715] = 12'h888;
rom[64716] = 12'h888;
rom[64717] = 12'h888;
rom[64718] = 12'h888;
rom[64719] = 12'h777;
rom[64720] = 12'h888;
rom[64721] = 12'h888;
rom[64722] = 12'h888;
rom[64723] = 12'h888;
rom[64724] = 12'h888;
rom[64725] = 12'h888;
rom[64726] = 12'h888;
rom[64727] = 12'h999;
rom[64728] = 12'h999;
rom[64729] = 12'h999;
rom[64730] = 12'h999;
rom[64731] = 12'h999;
rom[64732] = 12'h999;
rom[64733] = 12'haaa;
rom[64734] = 12'haaa;
rom[64735] = 12'haaa;
rom[64736] = 12'haaa;
rom[64737] = 12'hbbb;
rom[64738] = 12'hbbb;
rom[64739] = 12'hbbb;
rom[64740] = 12'hbbb;
rom[64741] = 12'hccc;
rom[64742] = 12'hccc;
rom[64743] = 12'hccc;
rom[64744] = 12'hddd;
rom[64745] = 12'hddd;
rom[64746] = 12'heee;
rom[64747] = 12'hfff;
rom[64748] = 12'hfff;
rom[64749] = 12'hfff;
rom[64750] = 12'hfff;
rom[64751] = 12'hfff;
rom[64752] = 12'hfff;
rom[64753] = 12'heee;
rom[64754] = 12'heee;
rom[64755] = 12'hddd;
rom[64756] = 12'hddd;
rom[64757] = 12'hddd;
rom[64758] = 12'hccc;
rom[64759] = 12'hccc;
rom[64760] = 12'hbbb;
rom[64761] = 12'hbbb;
rom[64762] = 12'hbbb;
rom[64763] = 12'hbbb;
rom[64764] = 12'hbbb;
rom[64765] = 12'haaa;
rom[64766] = 12'haaa;
rom[64767] = 12'haaa;
rom[64768] = 12'haaa;
rom[64769] = 12'haaa;
rom[64770] = 12'haaa;
rom[64771] = 12'hbbb;
rom[64772] = 12'hbbb;
rom[64773] = 12'hbbb;
rom[64774] = 12'hbbb;
rom[64775] = 12'hbbb;
rom[64776] = 12'hccc;
rom[64777] = 12'hccc;
rom[64778] = 12'hbbb;
rom[64779] = 12'haaa;
rom[64780] = 12'h999;
rom[64781] = 12'h888;
rom[64782] = 12'h888;
rom[64783] = 12'h888;
rom[64784] = 12'h777;
rom[64785] = 12'h777;
rom[64786] = 12'h777;
rom[64787] = 12'h777;
rom[64788] = 12'h777;
rom[64789] = 12'h777;
rom[64790] = 12'h777;
rom[64791] = 12'h777;
rom[64792] = 12'h666;
rom[64793] = 12'h666;
rom[64794] = 12'h666;
rom[64795] = 12'h666;
rom[64796] = 12'h666;
rom[64797] = 12'h777;
rom[64798] = 12'h777;
rom[64799] = 12'h777;
rom[64800] = 12'hfff;
rom[64801] = 12'hfff;
rom[64802] = 12'hfff;
rom[64803] = 12'hfff;
rom[64804] = 12'hfff;
rom[64805] = 12'hfff;
rom[64806] = 12'hfff;
rom[64807] = 12'hfff;
rom[64808] = 12'hfff;
rom[64809] = 12'hfff;
rom[64810] = 12'hfff;
rom[64811] = 12'hfff;
rom[64812] = 12'hfff;
rom[64813] = 12'hfff;
rom[64814] = 12'hfff;
rom[64815] = 12'hfff;
rom[64816] = 12'hfff;
rom[64817] = 12'hfff;
rom[64818] = 12'hfff;
rom[64819] = 12'hfff;
rom[64820] = 12'hfff;
rom[64821] = 12'hfff;
rom[64822] = 12'hfff;
rom[64823] = 12'hfff;
rom[64824] = 12'hfff;
rom[64825] = 12'hfff;
rom[64826] = 12'hfff;
rom[64827] = 12'hfff;
rom[64828] = 12'hfff;
rom[64829] = 12'hfff;
rom[64830] = 12'hfff;
rom[64831] = 12'hfff;
rom[64832] = 12'hfff;
rom[64833] = 12'hfff;
rom[64834] = 12'hfff;
rom[64835] = 12'hfff;
rom[64836] = 12'hfff;
rom[64837] = 12'hfff;
rom[64838] = 12'hfff;
rom[64839] = 12'hfff;
rom[64840] = 12'hfff;
rom[64841] = 12'hfff;
rom[64842] = 12'hfff;
rom[64843] = 12'hfff;
rom[64844] = 12'hfff;
rom[64845] = 12'hfff;
rom[64846] = 12'hfff;
rom[64847] = 12'hfff;
rom[64848] = 12'hfff;
rom[64849] = 12'hfff;
rom[64850] = 12'hfff;
rom[64851] = 12'hfff;
rom[64852] = 12'hfff;
rom[64853] = 12'hfff;
rom[64854] = 12'hfff;
rom[64855] = 12'hfff;
rom[64856] = 12'hfff;
rom[64857] = 12'hfff;
rom[64858] = 12'hfff;
rom[64859] = 12'hfff;
rom[64860] = 12'hfff;
rom[64861] = 12'hfff;
rom[64862] = 12'hfff;
rom[64863] = 12'hfff;
rom[64864] = 12'hfff;
rom[64865] = 12'hfff;
rom[64866] = 12'hfff;
rom[64867] = 12'hfff;
rom[64868] = 12'hfff;
rom[64869] = 12'hfff;
rom[64870] = 12'hfff;
rom[64871] = 12'hfff;
rom[64872] = 12'hfff;
rom[64873] = 12'hfff;
rom[64874] = 12'hfff;
rom[64875] = 12'hfff;
rom[64876] = 12'hfff;
rom[64877] = 12'hfff;
rom[64878] = 12'hfff;
rom[64879] = 12'hfff;
rom[64880] = 12'hfff;
rom[64881] = 12'hfff;
rom[64882] = 12'hfff;
rom[64883] = 12'hfff;
rom[64884] = 12'hfff;
rom[64885] = 12'hfff;
rom[64886] = 12'hfff;
rom[64887] = 12'hfff;
rom[64888] = 12'hfff;
rom[64889] = 12'hfff;
rom[64890] = 12'hfff;
rom[64891] = 12'hfff;
rom[64892] = 12'hfff;
rom[64893] = 12'hfff;
rom[64894] = 12'hfff;
rom[64895] = 12'hfff;
rom[64896] = 12'hfff;
rom[64897] = 12'hfff;
rom[64898] = 12'hfff;
rom[64899] = 12'hfff;
rom[64900] = 12'hfff;
rom[64901] = 12'hfff;
rom[64902] = 12'hfff;
rom[64903] = 12'hfff;
rom[64904] = 12'hfff;
rom[64905] = 12'hfff;
rom[64906] = 12'hfff;
rom[64907] = 12'hfff;
rom[64908] = 12'hfff;
rom[64909] = 12'hfff;
rom[64910] = 12'hfff;
rom[64911] = 12'heee;
rom[64912] = 12'heee;
rom[64913] = 12'heee;
rom[64914] = 12'hddd;
rom[64915] = 12'hddd;
rom[64916] = 12'hddd;
rom[64917] = 12'hddd;
rom[64918] = 12'hddd;
rom[64919] = 12'hddd;
rom[64920] = 12'hddd;
rom[64921] = 12'hccc;
rom[64922] = 12'hccc;
rom[64923] = 12'hccc;
rom[64924] = 12'hbbb;
rom[64925] = 12'hbbb;
rom[64926] = 12'haaa;
rom[64927] = 12'haaa;
rom[64928] = 12'h999;
rom[64929] = 12'h999;
rom[64930] = 12'h999;
rom[64931] = 12'h888;
rom[64932] = 12'h888;
rom[64933] = 12'h888;
rom[64934] = 12'h888;
rom[64935] = 12'h888;
rom[64936] = 12'h777;
rom[64937] = 12'h777;
rom[64938] = 12'h666;
rom[64939] = 12'h666;
rom[64940] = 12'h666;
rom[64941] = 12'h666;
rom[64942] = 12'h666;
rom[64943] = 12'h666;
rom[64944] = 12'h666;
rom[64945] = 12'h666;
rom[64946] = 12'h666;
rom[64947] = 12'h666;
rom[64948] = 12'h555;
rom[64949] = 12'h555;
rom[64950] = 12'h555;
rom[64951] = 12'h444;
rom[64952] = 12'h444;
rom[64953] = 12'h333;
rom[64954] = 12'h333;
rom[64955] = 12'h333;
rom[64956] = 12'h333;
rom[64957] = 12'h333;
rom[64958] = 12'h333;
rom[64959] = 12'h333;
rom[64960] = 12'h222;
rom[64961] = 12'h222;
rom[64962] = 12'h222;
rom[64963] = 12'h222;
rom[64964] = 12'h111;
rom[64965] = 12'h111;
rom[64966] = 12'h111;
rom[64967] = 12'h111;
rom[64968] = 12'h111;
rom[64969] = 12'h111;
rom[64970] = 12'h111;
rom[64971] = 12'h111;
rom[64972] = 12'h111;
rom[64973] = 12'h111;
rom[64974] = 12'h111;
rom[64975] = 12'h111;
rom[64976] = 12'h111;
rom[64977] = 12'h111;
rom[64978] = 12'h111;
rom[64979] = 12'h  0;
rom[64980] = 12'h  0;
rom[64981] = 12'h  0;
rom[64982] = 12'h  0;
rom[64983] = 12'h  0;
rom[64984] = 12'h  0;
rom[64985] = 12'h  0;
rom[64986] = 12'h  0;
rom[64987] = 12'h  0;
rom[64988] = 12'h  0;
rom[64989] = 12'h111;
rom[64990] = 12'h  0;
rom[64991] = 12'h  0;
rom[64992] = 12'h  0;
rom[64993] = 12'h  0;
rom[64994] = 12'h  0;
rom[64995] = 12'h  0;
rom[64996] = 12'h  0;
rom[64997] = 12'h  0;
rom[64998] = 12'h  0;
rom[64999] = 12'h  0;
rom[65000] = 12'h  0;
rom[65001] = 12'h  0;
rom[65002] = 12'h  0;
rom[65003] = 12'h  0;
rom[65004] = 12'h  0;
rom[65005] = 12'h  0;
rom[65006] = 12'h  0;
rom[65007] = 12'h  0;
rom[65008] = 12'h  0;
rom[65009] = 12'h111;
rom[65010] = 12'h111;
rom[65011] = 12'h111;
rom[65012] = 12'h111;
rom[65013] = 12'h111;
rom[65014] = 12'h111;
rom[65015] = 12'h111;
rom[65016] = 12'h111;
rom[65017] = 12'h111;
rom[65018] = 12'h  0;
rom[65019] = 12'h  0;
rom[65020] = 12'h  0;
rom[65021] = 12'h  0;
rom[65022] = 12'h  0;
rom[65023] = 12'h  0;
rom[65024] = 12'h  0;
rom[65025] = 12'h  0;
rom[65026] = 12'h  0;
rom[65027] = 12'h  0;
rom[65028] = 12'h  0;
rom[65029] = 12'h  0;
rom[65030] = 12'h  0;
rom[65031] = 12'h  0;
rom[65032] = 12'h  0;
rom[65033] = 12'h  0;
rom[65034] = 12'h  0;
rom[65035] = 12'h  0;
rom[65036] = 12'h  0;
rom[65037] = 12'h  0;
rom[65038] = 12'h  0;
rom[65039] = 12'h  0;
rom[65040] = 12'h  0;
rom[65041] = 12'h  0;
rom[65042] = 12'h  0;
rom[65043] = 12'h  0;
rom[65044] = 12'h  0;
rom[65045] = 12'h  0;
rom[65046] = 12'h  0;
rom[65047] = 12'h  0;
rom[65048] = 12'h  0;
rom[65049] = 12'h  0;
rom[65050] = 12'h  0;
rom[65051] = 12'h  0;
rom[65052] = 12'h  0;
rom[65053] = 12'h  0;
rom[65054] = 12'h  0;
rom[65055] = 12'h  0;
rom[65056] = 12'h  0;
rom[65057] = 12'h  0;
rom[65058] = 12'h  0;
rom[65059] = 12'h  0;
rom[65060] = 12'h  0;
rom[65061] = 12'h  0;
rom[65062] = 12'h  0;
rom[65063] = 12'h  0;
rom[65064] = 12'h  0;
rom[65065] = 12'h  0;
rom[65066] = 12'h  0;
rom[65067] = 12'h  0;
rom[65068] = 12'h  0;
rom[65069] = 12'h  0;
rom[65070] = 12'h  0;
rom[65071] = 12'h  0;
rom[65072] = 12'h111;
rom[65073] = 12'h111;
rom[65074] = 12'h111;
rom[65075] = 12'h222;
rom[65076] = 12'h222;
rom[65077] = 12'h333;
rom[65078] = 12'h444;
rom[65079] = 12'h555;
rom[65080] = 12'h444;
rom[65081] = 12'h444;
rom[65082] = 12'h444;
rom[65083] = 12'h333;
rom[65084] = 12'h222;
rom[65085] = 12'h111;
rom[65086] = 12'h111;
rom[65087] = 12'h111;
rom[65088] = 12'h111;
rom[65089] = 12'h111;
rom[65090] = 12'h111;
rom[65091] = 12'h111;
rom[65092] = 12'h111;
rom[65093] = 12'h111;
rom[65094] = 12'h111;
rom[65095] = 12'h111;
rom[65096] = 12'h222;
rom[65097] = 12'h222;
rom[65098] = 12'h333;
rom[65099] = 12'h444;
rom[65100] = 12'h444;
rom[65101] = 12'h444;
rom[65102] = 12'h444;
rom[65103] = 12'h333;
rom[65104] = 12'h444;
rom[65105] = 12'h444;
rom[65106] = 12'h444;
rom[65107] = 12'h444;
rom[65108] = 12'h444;
rom[65109] = 12'h444;
rom[65110] = 12'h555;
rom[65111] = 12'h555;
rom[65112] = 12'h666;
rom[65113] = 12'h666;
rom[65114] = 12'h777;
rom[65115] = 12'h777;
rom[65116] = 12'h888;
rom[65117] = 12'h888;
rom[65118] = 12'h888;
rom[65119] = 12'h888;
rom[65120] = 12'h888;
rom[65121] = 12'h888;
rom[65122] = 12'h888;
rom[65123] = 12'h888;
rom[65124] = 12'h888;
rom[65125] = 12'h888;
rom[65126] = 12'h999;
rom[65127] = 12'h999;
rom[65128] = 12'h999;
rom[65129] = 12'h999;
rom[65130] = 12'h999;
rom[65131] = 12'h999;
rom[65132] = 12'haaa;
rom[65133] = 12'haaa;
rom[65134] = 12'haaa;
rom[65135] = 12'haaa;
rom[65136] = 12'hbbb;
rom[65137] = 12'hbbb;
rom[65138] = 12'hbbb;
rom[65139] = 12'hbbb;
rom[65140] = 12'hccc;
rom[65141] = 12'hccc;
rom[65142] = 12'hccc;
rom[65143] = 12'hddd;
rom[65144] = 12'heee;
rom[65145] = 12'heee;
rom[65146] = 12'hfff;
rom[65147] = 12'hfff;
rom[65148] = 12'hfff;
rom[65149] = 12'hfff;
rom[65150] = 12'hfff;
rom[65151] = 12'hfff;
rom[65152] = 12'heee;
rom[65153] = 12'heee;
rom[65154] = 12'hddd;
rom[65155] = 12'hddd;
rom[65156] = 12'hddd;
rom[65157] = 12'hccc;
rom[65158] = 12'hccc;
rom[65159] = 12'hbbb;
rom[65160] = 12'hbbb;
rom[65161] = 12'hbbb;
rom[65162] = 12'hbbb;
rom[65163] = 12'haaa;
rom[65164] = 12'haaa;
rom[65165] = 12'haaa;
rom[65166] = 12'haaa;
rom[65167] = 12'haaa;
rom[65168] = 12'haaa;
rom[65169] = 12'haaa;
rom[65170] = 12'haaa;
rom[65171] = 12'haaa;
rom[65172] = 12'haaa;
rom[65173] = 12'hbbb;
rom[65174] = 12'hbbb;
rom[65175] = 12'hbbb;
rom[65176] = 12'hccc;
rom[65177] = 12'hccc;
rom[65178] = 12'hbbb;
rom[65179] = 12'haaa;
rom[65180] = 12'haaa;
rom[65181] = 12'h999;
rom[65182] = 12'h888;
rom[65183] = 12'h888;
rom[65184] = 12'h888;
rom[65185] = 12'h777;
rom[65186] = 12'h777;
rom[65187] = 12'h777;
rom[65188] = 12'h777;
rom[65189] = 12'h777;
rom[65190] = 12'h777;
rom[65191] = 12'h666;
rom[65192] = 12'h777;
rom[65193] = 12'h777;
rom[65194] = 12'h666;
rom[65195] = 12'h666;
rom[65196] = 12'h777;
rom[65197] = 12'h777;
rom[65198] = 12'h777;
rom[65199] = 12'h777;
rom[65200] = 12'hfff;
rom[65201] = 12'hfff;
rom[65202] = 12'hfff;
rom[65203] = 12'hfff;
rom[65204] = 12'hfff;
rom[65205] = 12'hfff;
rom[65206] = 12'hfff;
rom[65207] = 12'hfff;
rom[65208] = 12'hfff;
rom[65209] = 12'hfff;
rom[65210] = 12'hfff;
rom[65211] = 12'hfff;
rom[65212] = 12'hfff;
rom[65213] = 12'hfff;
rom[65214] = 12'hfff;
rom[65215] = 12'hfff;
rom[65216] = 12'hfff;
rom[65217] = 12'hfff;
rom[65218] = 12'hfff;
rom[65219] = 12'hfff;
rom[65220] = 12'hfff;
rom[65221] = 12'hfff;
rom[65222] = 12'hfff;
rom[65223] = 12'hfff;
rom[65224] = 12'hfff;
rom[65225] = 12'hfff;
rom[65226] = 12'hfff;
rom[65227] = 12'hfff;
rom[65228] = 12'hfff;
rom[65229] = 12'hfff;
rom[65230] = 12'hfff;
rom[65231] = 12'hfff;
rom[65232] = 12'hfff;
rom[65233] = 12'hfff;
rom[65234] = 12'hfff;
rom[65235] = 12'hfff;
rom[65236] = 12'hfff;
rom[65237] = 12'hfff;
rom[65238] = 12'hfff;
rom[65239] = 12'hfff;
rom[65240] = 12'hfff;
rom[65241] = 12'hfff;
rom[65242] = 12'hfff;
rom[65243] = 12'hfff;
rom[65244] = 12'hfff;
rom[65245] = 12'hfff;
rom[65246] = 12'hfff;
rom[65247] = 12'hfff;
rom[65248] = 12'hfff;
rom[65249] = 12'hfff;
rom[65250] = 12'hfff;
rom[65251] = 12'hfff;
rom[65252] = 12'hfff;
rom[65253] = 12'hfff;
rom[65254] = 12'hfff;
rom[65255] = 12'hfff;
rom[65256] = 12'hfff;
rom[65257] = 12'hfff;
rom[65258] = 12'hfff;
rom[65259] = 12'hfff;
rom[65260] = 12'hfff;
rom[65261] = 12'hfff;
rom[65262] = 12'hfff;
rom[65263] = 12'hfff;
rom[65264] = 12'hfff;
rom[65265] = 12'hfff;
rom[65266] = 12'hfff;
rom[65267] = 12'hfff;
rom[65268] = 12'hfff;
rom[65269] = 12'hfff;
rom[65270] = 12'hfff;
rom[65271] = 12'hfff;
rom[65272] = 12'hfff;
rom[65273] = 12'hfff;
rom[65274] = 12'hfff;
rom[65275] = 12'hfff;
rom[65276] = 12'hfff;
rom[65277] = 12'hfff;
rom[65278] = 12'hfff;
rom[65279] = 12'hfff;
rom[65280] = 12'hfff;
rom[65281] = 12'hfff;
rom[65282] = 12'hfff;
rom[65283] = 12'hfff;
rom[65284] = 12'hfff;
rom[65285] = 12'hfff;
rom[65286] = 12'hfff;
rom[65287] = 12'hfff;
rom[65288] = 12'hfff;
rom[65289] = 12'hfff;
rom[65290] = 12'hfff;
rom[65291] = 12'hfff;
rom[65292] = 12'hfff;
rom[65293] = 12'hfff;
rom[65294] = 12'hfff;
rom[65295] = 12'hfff;
rom[65296] = 12'hfff;
rom[65297] = 12'hfff;
rom[65298] = 12'hfff;
rom[65299] = 12'hfff;
rom[65300] = 12'hfff;
rom[65301] = 12'hfff;
rom[65302] = 12'hfff;
rom[65303] = 12'hfff;
rom[65304] = 12'hfff;
rom[65305] = 12'hfff;
rom[65306] = 12'hfff;
rom[65307] = 12'hfff;
rom[65308] = 12'hfff;
rom[65309] = 12'hfff;
rom[65310] = 12'hfff;
rom[65311] = 12'heee;
rom[65312] = 12'heee;
rom[65313] = 12'heee;
rom[65314] = 12'hddd;
rom[65315] = 12'hddd;
rom[65316] = 12'hddd;
rom[65317] = 12'hddd;
rom[65318] = 12'hccc;
rom[65319] = 12'hccc;
rom[65320] = 12'hccc;
rom[65321] = 12'hccc;
rom[65322] = 12'hccc;
rom[65323] = 12'hccc;
rom[65324] = 12'hccc;
rom[65325] = 12'hbbb;
rom[65326] = 12'hbbb;
rom[65327] = 12'hbbb;
rom[65328] = 12'haaa;
rom[65329] = 12'haaa;
rom[65330] = 12'h999;
rom[65331] = 12'h999;
rom[65332] = 12'h999;
rom[65333] = 12'h999;
rom[65334] = 12'h888;
rom[65335] = 12'h888;
rom[65336] = 12'h777;
rom[65337] = 12'h777;
rom[65338] = 12'h777;
rom[65339] = 12'h666;
rom[65340] = 12'h666;
rom[65341] = 12'h666;
rom[65342] = 12'h666;
rom[65343] = 12'h666;
rom[65344] = 12'h555;
rom[65345] = 12'h666;
rom[65346] = 12'h666;
rom[65347] = 12'h666;
rom[65348] = 12'h666;
rom[65349] = 12'h555;
rom[65350] = 12'h555;
rom[65351] = 12'h444;
rom[65352] = 12'h444;
rom[65353] = 12'h444;
rom[65354] = 12'h444;
rom[65355] = 12'h333;
rom[65356] = 12'h333;
rom[65357] = 12'h333;
rom[65358] = 12'h333;
rom[65359] = 12'h333;
rom[65360] = 12'h333;
rom[65361] = 12'h222;
rom[65362] = 12'h222;
rom[65363] = 12'h222;
rom[65364] = 12'h111;
rom[65365] = 12'h111;
rom[65366] = 12'h111;
rom[65367] = 12'h111;
rom[65368] = 12'h111;
rom[65369] = 12'h111;
rom[65370] = 12'h111;
rom[65371] = 12'h111;
rom[65372] = 12'h111;
rom[65373] = 12'h111;
rom[65374] = 12'h111;
rom[65375] = 12'h111;
rom[65376] = 12'h111;
rom[65377] = 12'h111;
rom[65378] = 12'h111;
rom[65379] = 12'h111;
rom[65380] = 12'h  0;
rom[65381] = 12'h111;
rom[65382] = 12'h111;
rom[65383] = 12'h111;
rom[65384] = 12'h  0;
rom[65385] = 12'h  0;
rom[65386] = 12'h  0;
rom[65387] = 12'h  0;
rom[65388] = 12'h  0;
rom[65389] = 12'h111;
rom[65390] = 12'h  0;
rom[65391] = 12'h  0;
rom[65392] = 12'h  0;
rom[65393] = 12'h  0;
rom[65394] = 12'h  0;
rom[65395] = 12'h  0;
rom[65396] = 12'h  0;
rom[65397] = 12'h  0;
rom[65398] = 12'h  0;
rom[65399] = 12'h  0;
rom[65400] = 12'h  0;
rom[65401] = 12'h  0;
rom[65402] = 12'h  0;
rom[65403] = 12'h  0;
rom[65404] = 12'h  0;
rom[65405] = 12'h  0;
rom[65406] = 12'h  0;
rom[65407] = 12'h  0;
rom[65408] = 12'h111;
rom[65409] = 12'h111;
rom[65410] = 12'h111;
rom[65411] = 12'h111;
rom[65412] = 12'h111;
rom[65413] = 12'h111;
rom[65414] = 12'h111;
rom[65415] = 12'h111;
rom[65416] = 12'h111;
rom[65417] = 12'h  0;
rom[65418] = 12'h  0;
rom[65419] = 12'h  0;
rom[65420] = 12'h  0;
rom[65421] = 12'h  0;
rom[65422] = 12'h  0;
rom[65423] = 12'h  0;
rom[65424] = 12'h  0;
rom[65425] = 12'h  0;
rom[65426] = 12'h  0;
rom[65427] = 12'h  0;
rom[65428] = 12'h  0;
rom[65429] = 12'h  0;
rom[65430] = 12'h  0;
rom[65431] = 12'h  0;
rom[65432] = 12'h  0;
rom[65433] = 12'h  0;
rom[65434] = 12'h  0;
rom[65435] = 12'h  0;
rom[65436] = 12'h  0;
rom[65437] = 12'h  0;
rom[65438] = 12'h  0;
rom[65439] = 12'h  0;
rom[65440] = 12'h  0;
rom[65441] = 12'h  0;
rom[65442] = 12'h  0;
rom[65443] = 12'h  0;
rom[65444] = 12'h  0;
rom[65445] = 12'h  0;
rom[65446] = 12'h  0;
rom[65447] = 12'h  0;
rom[65448] = 12'h  0;
rom[65449] = 12'h  0;
rom[65450] = 12'h  0;
rom[65451] = 12'h  0;
rom[65452] = 12'h  0;
rom[65453] = 12'h  0;
rom[65454] = 12'h  0;
rom[65455] = 12'h  0;
rom[65456] = 12'h  0;
rom[65457] = 12'h  0;
rom[65458] = 12'h  0;
rom[65459] = 12'h  0;
rom[65460] = 12'h  0;
rom[65461] = 12'h  0;
rom[65462] = 12'h  0;
rom[65463] = 12'h  0;
rom[65464] = 12'h  0;
rom[65465] = 12'h  0;
rom[65466] = 12'h  0;
rom[65467] = 12'h  0;
rom[65468] = 12'h  0;
rom[65469] = 12'h  0;
rom[65470] = 12'h  0;
rom[65471] = 12'h  0;
rom[65472] = 12'h  0;
rom[65473] = 12'h111;
rom[65474] = 12'h111;
rom[65475] = 12'h222;
rom[65476] = 12'h333;
rom[65477] = 12'h333;
rom[65478] = 12'h444;
rom[65479] = 12'h555;
rom[65480] = 12'h444;
rom[65481] = 12'h444;
rom[65482] = 12'h444;
rom[65483] = 12'h333;
rom[65484] = 12'h222;
rom[65485] = 12'h111;
rom[65486] = 12'h111;
rom[65487] = 12'h111;
rom[65488] = 12'h111;
rom[65489] = 12'h111;
rom[65490] = 12'h111;
rom[65491] = 12'h111;
rom[65492] = 12'h111;
rom[65493] = 12'h111;
rom[65494] = 12'h111;
rom[65495] = 12'h111;
rom[65496] = 12'h222;
rom[65497] = 12'h222;
rom[65498] = 12'h333;
rom[65499] = 12'h333;
rom[65500] = 12'h444;
rom[65501] = 12'h444;
rom[65502] = 12'h444;
rom[65503] = 12'h333;
rom[65504] = 12'h444;
rom[65505] = 12'h444;
rom[65506] = 12'h444;
rom[65507] = 12'h444;
rom[65508] = 12'h444;
rom[65509] = 12'h444;
rom[65510] = 12'h444;
rom[65511] = 12'h555;
rom[65512] = 12'h555;
rom[65513] = 12'h666;
rom[65514] = 12'h777;
rom[65515] = 12'h777;
rom[65516] = 12'h888;
rom[65517] = 12'h888;
rom[65518] = 12'h888;
rom[65519] = 12'h888;
rom[65520] = 12'h888;
rom[65521] = 12'h888;
rom[65522] = 12'h888;
rom[65523] = 12'h888;
rom[65524] = 12'h888;
rom[65525] = 12'h999;
rom[65526] = 12'h999;
rom[65527] = 12'h999;
rom[65528] = 12'h999;
rom[65529] = 12'h999;
rom[65530] = 12'h999;
rom[65531] = 12'haaa;
rom[65532] = 12'haaa;
rom[65533] = 12'haaa;
rom[65534] = 12'hbbb;
rom[65535] = 12'hbbb;
rom[65536] = 12'hbbb;
rom[65537] = 12'hbbb;
rom[65538] = 12'hbbb;
rom[65539] = 12'hccc;
rom[65540] = 12'hccc;
rom[65541] = 12'hccc;
rom[65542] = 12'hddd;
rom[65543] = 12'hddd;
rom[65544] = 12'heee;
rom[65545] = 12'hfff;
rom[65546] = 12'hfff;
rom[65547] = 12'hfff;
rom[65548] = 12'hfff;
rom[65549] = 12'hfff;
rom[65550] = 12'hfff;
rom[65551] = 12'heee;
rom[65552] = 12'heee;
rom[65553] = 12'heee;
rom[65554] = 12'hddd;
rom[65555] = 12'hddd;
rom[65556] = 12'hccc;
rom[65557] = 12'hccc;
rom[65558] = 12'hccc;
rom[65559] = 12'hbbb;
rom[65560] = 12'hbbb;
rom[65561] = 12'hbbb;
rom[65562] = 12'hbbb;
rom[65563] = 12'haaa;
rom[65564] = 12'haaa;
rom[65565] = 12'haaa;
rom[65566] = 12'haaa;
rom[65567] = 12'haaa;
rom[65568] = 12'haaa;
rom[65569] = 12'haaa;
rom[65570] = 12'h999;
rom[65571] = 12'h999;
rom[65572] = 12'haaa;
rom[65573] = 12'haaa;
rom[65574] = 12'haaa;
rom[65575] = 12'hbbb;
rom[65576] = 12'hccc;
rom[65577] = 12'hccc;
rom[65578] = 12'hbbb;
rom[65579] = 12'hbbb;
rom[65580] = 12'haaa;
rom[65581] = 12'h999;
rom[65582] = 12'h999;
rom[65583] = 12'h888;
rom[65584] = 12'h888;
rom[65585] = 12'h777;
rom[65586] = 12'h777;
rom[65587] = 12'h777;
rom[65588] = 12'h777;
rom[65589] = 12'h777;
rom[65590] = 12'h777;
rom[65591] = 12'h666;
rom[65592] = 12'h777;
rom[65593] = 12'h777;
rom[65594] = 12'h777;
rom[65595] = 12'h777;
rom[65596] = 12'h777;
rom[65597] = 12'h777;
rom[65598] = 12'h777;
rom[65599] = 12'h777;
rom[65600] = 12'hfff;
rom[65601] = 12'hfff;
rom[65602] = 12'hfff;
rom[65603] = 12'hfff;
rom[65604] = 12'hfff;
rom[65605] = 12'hfff;
rom[65606] = 12'hfff;
rom[65607] = 12'hfff;
rom[65608] = 12'hfff;
rom[65609] = 12'hfff;
rom[65610] = 12'hfff;
rom[65611] = 12'hfff;
rom[65612] = 12'hfff;
rom[65613] = 12'hfff;
rom[65614] = 12'hfff;
rom[65615] = 12'hfff;
rom[65616] = 12'hfff;
rom[65617] = 12'hfff;
rom[65618] = 12'hfff;
rom[65619] = 12'hfff;
rom[65620] = 12'hfff;
rom[65621] = 12'hfff;
rom[65622] = 12'hfff;
rom[65623] = 12'hfff;
rom[65624] = 12'hfff;
rom[65625] = 12'hfff;
rom[65626] = 12'hfff;
rom[65627] = 12'hfff;
rom[65628] = 12'hfff;
rom[65629] = 12'hfff;
rom[65630] = 12'hfff;
rom[65631] = 12'hfff;
rom[65632] = 12'hfff;
rom[65633] = 12'hfff;
rom[65634] = 12'hfff;
rom[65635] = 12'hfff;
rom[65636] = 12'hfff;
rom[65637] = 12'hfff;
rom[65638] = 12'hfff;
rom[65639] = 12'hfff;
rom[65640] = 12'hfff;
rom[65641] = 12'hfff;
rom[65642] = 12'hfff;
rom[65643] = 12'hfff;
rom[65644] = 12'hfff;
rom[65645] = 12'hfff;
rom[65646] = 12'hfff;
rom[65647] = 12'hfff;
rom[65648] = 12'hfff;
rom[65649] = 12'hfff;
rom[65650] = 12'hfff;
rom[65651] = 12'hfff;
rom[65652] = 12'hfff;
rom[65653] = 12'hfff;
rom[65654] = 12'hfff;
rom[65655] = 12'hfff;
rom[65656] = 12'hfff;
rom[65657] = 12'hfff;
rom[65658] = 12'hfff;
rom[65659] = 12'hfff;
rom[65660] = 12'hfff;
rom[65661] = 12'hfff;
rom[65662] = 12'hfff;
rom[65663] = 12'hfff;
rom[65664] = 12'hfff;
rom[65665] = 12'hfff;
rom[65666] = 12'hfff;
rom[65667] = 12'hfff;
rom[65668] = 12'hfff;
rom[65669] = 12'hfff;
rom[65670] = 12'hfff;
rom[65671] = 12'hfff;
rom[65672] = 12'hfff;
rom[65673] = 12'hfff;
rom[65674] = 12'hfff;
rom[65675] = 12'hfff;
rom[65676] = 12'hfff;
rom[65677] = 12'hfff;
rom[65678] = 12'hfff;
rom[65679] = 12'hfff;
rom[65680] = 12'hfff;
rom[65681] = 12'hfff;
rom[65682] = 12'hfff;
rom[65683] = 12'hfff;
rom[65684] = 12'hfff;
rom[65685] = 12'hfff;
rom[65686] = 12'hfff;
rom[65687] = 12'hfff;
rom[65688] = 12'hfff;
rom[65689] = 12'hfff;
rom[65690] = 12'hfff;
rom[65691] = 12'hfff;
rom[65692] = 12'hfff;
rom[65693] = 12'hfff;
rom[65694] = 12'hfff;
rom[65695] = 12'hfff;
rom[65696] = 12'hfff;
rom[65697] = 12'hfff;
rom[65698] = 12'hfff;
rom[65699] = 12'hfff;
rom[65700] = 12'hfff;
rom[65701] = 12'hfff;
rom[65702] = 12'hfff;
rom[65703] = 12'hfff;
rom[65704] = 12'hfff;
rom[65705] = 12'hfff;
rom[65706] = 12'hfff;
rom[65707] = 12'hfff;
rom[65708] = 12'hfff;
rom[65709] = 12'hfff;
rom[65710] = 12'hfff;
rom[65711] = 12'heee;
rom[65712] = 12'heee;
rom[65713] = 12'heee;
rom[65714] = 12'hddd;
rom[65715] = 12'hddd;
rom[65716] = 12'hddd;
rom[65717] = 12'hccc;
rom[65718] = 12'hccc;
rom[65719] = 12'hccc;
rom[65720] = 12'hccc;
rom[65721] = 12'hbbb;
rom[65722] = 12'hbbb;
rom[65723] = 12'hbbb;
rom[65724] = 12'hbbb;
rom[65725] = 12'hbbb;
rom[65726] = 12'hbbb;
rom[65727] = 12'hbbb;
rom[65728] = 12'haaa;
rom[65729] = 12'haaa;
rom[65730] = 12'haaa;
rom[65731] = 12'h999;
rom[65732] = 12'h999;
rom[65733] = 12'h999;
rom[65734] = 12'h999;
rom[65735] = 12'h999;
rom[65736] = 12'h888;
rom[65737] = 12'h888;
rom[65738] = 12'h777;
rom[65739] = 12'h777;
rom[65740] = 12'h666;
rom[65741] = 12'h666;
rom[65742] = 12'h555;
rom[65743] = 12'h555;
rom[65744] = 12'h555;
rom[65745] = 12'h555;
rom[65746] = 12'h666;
rom[65747] = 12'h666;
rom[65748] = 12'h666;
rom[65749] = 12'h666;
rom[65750] = 12'h555;
rom[65751] = 12'h555;
rom[65752] = 12'h444;
rom[65753] = 12'h444;
rom[65754] = 12'h444;
rom[65755] = 12'h444;
rom[65756] = 12'h333;
rom[65757] = 12'h333;
rom[65758] = 12'h333;
rom[65759] = 12'h333;
rom[65760] = 12'h333;
rom[65761] = 12'h333;
rom[65762] = 12'h222;
rom[65763] = 12'h222;
rom[65764] = 12'h222;
rom[65765] = 12'h222;
rom[65766] = 12'h222;
rom[65767] = 12'h111;
rom[65768] = 12'h111;
rom[65769] = 12'h111;
rom[65770] = 12'h111;
rom[65771] = 12'h111;
rom[65772] = 12'h111;
rom[65773] = 12'h111;
rom[65774] = 12'h111;
rom[65775] = 12'h111;
rom[65776] = 12'h111;
rom[65777] = 12'h111;
rom[65778] = 12'h111;
rom[65779] = 12'h111;
rom[65780] = 12'h111;
rom[65781] = 12'h111;
rom[65782] = 12'h111;
rom[65783] = 12'h111;
rom[65784] = 12'h111;
rom[65785] = 12'h  0;
rom[65786] = 12'h  0;
rom[65787] = 12'h  0;
rom[65788] = 12'h111;
rom[65789] = 12'h111;
rom[65790] = 12'h  0;
rom[65791] = 12'h  0;
rom[65792] = 12'h  0;
rom[65793] = 12'h  0;
rom[65794] = 12'h  0;
rom[65795] = 12'h  0;
rom[65796] = 12'h  0;
rom[65797] = 12'h  0;
rom[65798] = 12'h  0;
rom[65799] = 12'h  0;
rom[65800] = 12'h  0;
rom[65801] = 12'h  0;
rom[65802] = 12'h  0;
rom[65803] = 12'h  0;
rom[65804] = 12'h  0;
rom[65805] = 12'h  0;
rom[65806] = 12'h  0;
rom[65807] = 12'h  0;
rom[65808] = 12'h111;
rom[65809] = 12'h111;
rom[65810] = 12'h111;
rom[65811] = 12'h111;
rom[65812] = 12'h111;
rom[65813] = 12'h111;
rom[65814] = 12'h111;
rom[65815] = 12'h111;
rom[65816] = 12'h  0;
rom[65817] = 12'h  0;
rom[65818] = 12'h  0;
rom[65819] = 12'h  0;
rom[65820] = 12'h  0;
rom[65821] = 12'h  0;
rom[65822] = 12'h  0;
rom[65823] = 12'h  0;
rom[65824] = 12'h  0;
rom[65825] = 12'h  0;
rom[65826] = 12'h  0;
rom[65827] = 12'h  0;
rom[65828] = 12'h  0;
rom[65829] = 12'h  0;
rom[65830] = 12'h  0;
rom[65831] = 12'h  0;
rom[65832] = 12'h  0;
rom[65833] = 12'h  0;
rom[65834] = 12'h  0;
rom[65835] = 12'h  0;
rom[65836] = 12'h  0;
rom[65837] = 12'h  0;
rom[65838] = 12'h  0;
rom[65839] = 12'h  0;
rom[65840] = 12'h  0;
rom[65841] = 12'h  0;
rom[65842] = 12'h  0;
rom[65843] = 12'h  0;
rom[65844] = 12'h  0;
rom[65845] = 12'h  0;
rom[65846] = 12'h  0;
rom[65847] = 12'h  0;
rom[65848] = 12'h  0;
rom[65849] = 12'h  0;
rom[65850] = 12'h  0;
rom[65851] = 12'h  0;
rom[65852] = 12'h  0;
rom[65853] = 12'h  0;
rom[65854] = 12'h  0;
rom[65855] = 12'h  0;
rom[65856] = 12'h  0;
rom[65857] = 12'h  0;
rom[65858] = 12'h  0;
rom[65859] = 12'h  0;
rom[65860] = 12'h  0;
rom[65861] = 12'h  0;
rom[65862] = 12'h  0;
rom[65863] = 12'h  0;
rom[65864] = 12'h  0;
rom[65865] = 12'h  0;
rom[65866] = 12'h  0;
rom[65867] = 12'h  0;
rom[65868] = 12'h  0;
rom[65869] = 12'h  0;
rom[65870] = 12'h  0;
rom[65871] = 12'h  0;
rom[65872] = 12'h  0;
rom[65873] = 12'h111;
rom[65874] = 12'h111;
rom[65875] = 12'h222;
rom[65876] = 12'h333;
rom[65877] = 12'h444;
rom[65878] = 12'h444;
rom[65879] = 12'h555;
rom[65880] = 12'h444;
rom[65881] = 12'h555;
rom[65882] = 12'h444;
rom[65883] = 12'h333;
rom[65884] = 12'h222;
rom[65885] = 12'h111;
rom[65886] = 12'h111;
rom[65887] = 12'h111;
rom[65888] = 12'h111;
rom[65889] = 12'h111;
rom[65890] = 12'h111;
rom[65891] = 12'h111;
rom[65892] = 12'h111;
rom[65893] = 12'h111;
rom[65894] = 12'h111;
rom[65895] = 12'h111;
rom[65896] = 12'h222;
rom[65897] = 12'h222;
rom[65898] = 12'h333;
rom[65899] = 12'h333;
rom[65900] = 12'h444;
rom[65901] = 12'h444;
rom[65902] = 12'h444;
rom[65903] = 12'h333;
rom[65904] = 12'h444;
rom[65905] = 12'h444;
rom[65906] = 12'h444;
rom[65907] = 12'h444;
rom[65908] = 12'h444;
rom[65909] = 12'h444;
rom[65910] = 12'h444;
rom[65911] = 12'h555;
rom[65912] = 12'h555;
rom[65913] = 12'h666;
rom[65914] = 12'h777;
rom[65915] = 12'h777;
rom[65916] = 12'h888;
rom[65917] = 12'h888;
rom[65918] = 12'h888;
rom[65919] = 12'h888;
rom[65920] = 12'h888;
rom[65921] = 12'h888;
rom[65922] = 12'h888;
rom[65923] = 12'h888;
rom[65924] = 12'h999;
rom[65925] = 12'h999;
rom[65926] = 12'h999;
rom[65927] = 12'h999;
rom[65928] = 12'h999;
rom[65929] = 12'h999;
rom[65930] = 12'haaa;
rom[65931] = 12'haaa;
rom[65932] = 12'haaa;
rom[65933] = 12'haaa;
rom[65934] = 12'hbbb;
rom[65935] = 12'hbbb;
rom[65936] = 12'hbbb;
rom[65937] = 12'hbbb;
rom[65938] = 12'hccc;
rom[65939] = 12'hccc;
rom[65940] = 12'hccc;
rom[65941] = 12'hddd;
rom[65942] = 12'hddd;
rom[65943] = 12'heee;
rom[65944] = 12'hfff;
rom[65945] = 12'hfff;
rom[65946] = 12'hfff;
rom[65947] = 12'hfff;
rom[65948] = 12'hfff;
rom[65949] = 12'hfff;
rom[65950] = 12'hfff;
rom[65951] = 12'heee;
rom[65952] = 12'heee;
rom[65953] = 12'hddd;
rom[65954] = 12'hddd;
rom[65955] = 12'hccc;
rom[65956] = 12'hccc;
rom[65957] = 12'hccc;
rom[65958] = 12'hbbb;
rom[65959] = 12'hbbb;
rom[65960] = 12'hbbb;
rom[65961] = 12'hbbb;
rom[65962] = 12'hbbb;
rom[65963] = 12'haaa;
rom[65964] = 12'haaa;
rom[65965] = 12'haaa;
rom[65966] = 12'haaa;
rom[65967] = 12'haaa;
rom[65968] = 12'h999;
rom[65969] = 12'h999;
rom[65970] = 12'h999;
rom[65971] = 12'h999;
rom[65972] = 12'h999;
rom[65973] = 12'h999;
rom[65974] = 12'haaa;
rom[65975] = 12'haaa;
rom[65976] = 12'hbbb;
rom[65977] = 12'hbbb;
rom[65978] = 12'hbbb;
rom[65979] = 12'hccc;
rom[65980] = 12'hbbb;
rom[65981] = 12'haaa;
rom[65982] = 12'h999;
rom[65983] = 12'h888;
rom[65984] = 12'h888;
rom[65985] = 12'h888;
rom[65986] = 12'h777;
rom[65987] = 12'h777;
rom[65988] = 12'h777;
rom[65989] = 12'h777;
rom[65990] = 12'h777;
rom[65991] = 12'h777;
rom[65992] = 12'h777;
rom[65993] = 12'h777;
rom[65994] = 12'h777;
rom[65995] = 12'h777;
rom[65996] = 12'h777;
rom[65997] = 12'h777;
rom[65998] = 12'h777;
rom[65999] = 12'h777;
rom[66000] = 12'hfff;
rom[66001] = 12'hfff;
rom[66002] = 12'hfff;
rom[66003] = 12'hfff;
rom[66004] = 12'hfff;
rom[66005] = 12'hfff;
rom[66006] = 12'hfff;
rom[66007] = 12'hfff;
rom[66008] = 12'hfff;
rom[66009] = 12'hfff;
rom[66010] = 12'hfff;
rom[66011] = 12'hfff;
rom[66012] = 12'hfff;
rom[66013] = 12'hfff;
rom[66014] = 12'hfff;
rom[66015] = 12'hfff;
rom[66016] = 12'hfff;
rom[66017] = 12'hfff;
rom[66018] = 12'hfff;
rom[66019] = 12'hfff;
rom[66020] = 12'hfff;
rom[66021] = 12'hfff;
rom[66022] = 12'hfff;
rom[66023] = 12'hfff;
rom[66024] = 12'hfff;
rom[66025] = 12'hfff;
rom[66026] = 12'hfff;
rom[66027] = 12'hfff;
rom[66028] = 12'hfff;
rom[66029] = 12'hfff;
rom[66030] = 12'hfff;
rom[66031] = 12'hfff;
rom[66032] = 12'hfff;
rom[66033] = 12'hfff;
rom[66034] = 12'hfff;
rom[66035] = 12'hfff;
rom[66036] = 12'hfff;
rom[66037] = 12'hfff;
rom[66038] = 12'hfff;
rom[66039] = 12'hfff;
rom[66040] = 12'hfff;
rom[66041] = 12'hfff;
rom[66042] = 12'hfff;
rom[66043] = 12'hfff;
rom[66044] = 12'hfff;
rom[66045] = 12'hfff;
rom[66046] = 12'hfff;
rom[66047] = 12'hfff;
rom[66048] = 12'hfff;
rom[66049] = 12'hfff;
rom[66050] = 12'hfff;
rom[66051] = 12'hfff;
rom[66052] = 12'hfff;
rom[66053] = 12'hfff;
rom[66054] = 12'hfff;
rom[66055] = 12'hfff;
rom[66056] = 12'hfff;
rom[66057] = 12'hfff;
rom[66058] = 12'hfff;
rom[66059] = 12'hfff;
rom[66060] = 12'hfff;
rom[66061] = 12'hfff;
rom[66062] = 12'hfff;
rom[66063] = 12'hfff;
rom[66064] = 12'hfff;
rom[66065] = 12'hfff;
rom[66066] = 12'hfff;
rom[66067] = 12'hfff;
rom[66068] = 12'hfff;
rom[66069] = 12'hfff;
rom[66070] = 12'hfff;
rom[66071] = 12'hfff;
rom[66072] = 12'hfff;
rom[66073] = 12'hfff;
rom[66074] = 12'hfff;
rom[66075] = 12'hfff;
rom[66076] = 12'hfff;
rom[66077] = 12'hfff;
rom[66078] = 12'hfff;
rom[66079] = 12'hfff;
rom[66080] = 12'hfff;
rom[66081] = 12'hfff;
rom[66082] = 12'hfff;
rom[66083] = 12'hfff;
rom[66084] = 12'hfff;
rom[66085] = 12'hfff;
rom[66086] = 12'hfff;
rom[66087] = 12'hfff;
rom[66088] = 12'hfff;
rom[66089] = 12'hfff;
rom[66090] = 12'hfff;
rom[66091] = 12'hfff;
rom[66092] = 12'hfff;
rom[66093] = 12'hfff;
rom[66094] = 12'hfff;
rom[66095] = 12'hfff;
rom[66096] = 12'hfff;
rom[66097] = 12'hfff;
rom[66098] = 12'hfff;
rom[66099] = 12'hfff;
rom[66100] = 12'hfff;
rom[66101] = 12'hfff;
rom[66102] = 12'hfff;
rom[66103] = 12'hfff;
rom[66104] = 12'hfff;
rom[66105] = 12'hfff;
rom[66106] = 12'hfff;
rom[66107] = 12'hfff;
rom[66108] = 12'hfff;
rom[66109] = 12'hfff;
rom[66110] = 12'hfff;
rom[66111] = 12'heee;
rom[66112] = 12'heee;
rom[66113] = 12'heee;
rom[66114] = 12'hddd;
rom[66115] = 12'hddd;
rom[66116] = 12'hddd;
rom[66117] = 12'hccc;
rom[66118] = 12'hccc;
rom[66119] = 12'hccc;
rom[66120] = 12'hbbb;
rom[66121] = 12'hbbb;
rom[66122] = 12'haaa;
rom[66123] = 12'haaa;
rom[66124] = 12'haaa;
rom[66125] = 12'haaa;
rom[66126] = 12'haaa;
rom[66127] = 12'haaa;
rom[66128] = 12'haaa;
rom[66129] = 12'h999;
rom[66130] = 12'h999;
rom[66131] = 12'h999;
rom[66132] = 12'h999;
rom[66133] = 12'h999;
rom[66134] = 12'h999;
rom[66135] = 12'h999;
rom[66136] = 12'h999;
rom[66137] = 12'h999;
rom[66138] = 12'h888;
rom[66139] = 12'h777;
rom[66140] = 12'h666;
rom[66141] = 12'h666;
rom[66142] = 12'h666;
rom[66143] = 12'h555;
rom[66144] = 12'h555;
rom[66145] = 12'h555;
rom[66146] = 12'h555;
rom[66147] = 12'h666;
rom[66148] = 12'h666;
rom[66149] = 12'h666;
rom[66150] = 12'h555;
rom[66151] = 12'h555;
rom[66152] = 12'h444;
rom[66153] = 12'h444;
rom[66154] = 12'h444;
rom[66155] = 12'h444;
rom[66156] = 12'h333;
rom[66157] = 12'h333;
rom[66158] = 12'h333;
rom[66159] = 12'h333;
rom[66160] = 12'h333;
rom[66161] = 12'h333;
rom[66162] = 12'h222;
rom[66163] = 12'h222;
rom[66164] = 12'h222;
rom[66165] = 12'h222;
rom[66166] = 12'h222;
rom[66167] = 12'h222;
rom[66168] = 12'h111;
rom[66169] = 12'h111;
rom[66170] = 12'h111;
rom[66171] = 12'h111;
rom[66172] = 12'h111;
rom[66173] = 12'h111;
rom[66174] = 12'h111;
rom[66175] = 12'h111;
rom[66176] = 12'h111;
rom[66177] = 12'h111;
rom[66178] = 12'h111;
rom[66179] = 12'h111;
rom[66180] = 12'h111;
rom[66181] = 12'h111;
rom[66182] = 12'h111;
rom[66183] = 12'h111;
rom[66184] = 12'h111;
rom[66185] = 12'h111;
rom[66186] = 12'h111;
rom[66187] = 12'h111;
rom[66188] = 12'h111;
rom[66189] = 12'h111;
rom[66190] = 12'h  0;
rom[66191] = 12'h  0;
rom[66192] = 12'h  0;
rom[66193] = 12'h  0;
rom[66194] = 12'h  0;
rom[66195] = 12'h  0;
rom[66196] = 12'h  0;
rom[66197] = 12'h  0;
rom[66198] = 12'h  0;
rom[66199] = 12'h  0;
rom[66200] = 12'h  0;
rom[66201] = 12'h  0;
rom[66202] = 12'h  0;
rom[66203] = 12'h  0;
rom[66204] = 12'h  0;
rom[66205] = 12'h  0;
rom[66206] = 12'h  0;
rom[66207] = 12'h111;
rom[66208] = 12'h111;
rom[66209] = 12'h111;
rom[66210] = 12'h111;
rom[66211] = 12'h111;
rom[66212] = 12'h111;
rom[66213] = 12'h111;
rom[66214] = 12'h111;
rom[66215] = 12'h111;
rom[66216] = 12'h  0;
rom[66217] = 12'h  0;
rom[66218] = 12'h111;
rom[66219] = 12'h111;
rom[66220] = 12'h111;
rom[66221] = 12'h  0;
rom[66222] = 12'h  0;
rom[66223] = 12'h  0;
rom[66224] = 12'h  0;
rom[66225] = 12'h  0;
rom[66226] = 12'h  0;
rom[66227] = 12'h  0;
rom[66228] = 12'h  0;
rom[66229] = 12'h  0;
rom[66230] = 12'h  0;
rom[66231] = 12'h  0;
rom[66232] = 12'h  0;
rom[66233] = 12'h  0;
rom[66234] = 12'h  0;
rom[66235] = 12'h  0;
rom[66236] = 12'h  0;
rom[66237] = 12'h  0;
rom[66238] = 12'h  0;
rom[66239] = 12'h  0;
rom[66240] = 12'h  0;
rom[66241] = 12'h  0;
rom[66242] = 12'h  0;
rom[66243] = 12'h  0;
rom[66244] = 12'h  0;
rom[66245] = 12'h  0;
rom[66246] = 12'h  0;
rom[66247] = 12'h  0;
rom[66248] = 12'h  0;
rom[66249] = 12'h  0;
rom[66250] = 12'h  0;
rom[66251] = 12'h  0;
rom[66252] = 12'h  0;
rom[66253] = 12'h  0;
rom[66254] = 12'h  0;
rom[66255] = 12'h  0;
rom[66256] = 12'h  0;
rom[66257] = 12'h  0;
rom[66258] = 12'h  0;
rom[66259] = 12'h  0;
rom[66260] = 12'h  0;
rom[66261] = 12'h  0;
rom[66262] = 12'h  0;
rom[66263] = 12'h  0;
rom[66264] = 12'h  0;
rom[66265] = 12'h  0;
rom[66266] = 12'h  0;
rom[66267] = 12'h  0;
rom[66268] = 12'h  0;
rom[66269] = 12'h  0;
rom[66270] = 12'h  0;
rom[66271] = 12'h  0;
rom[66272] = 12'h  0;
rom[66273] = 12'h111;
rom[66274] = 12'h111;
rom[66275] = 12'h222;
rom[66276] = 12'h333;
rom[66277] = 12'h444;
rom[66278] = 12'h444;
rom[66279] = 12'h555;
rom[66280] = 12'h555;
rom[66281] = 12'h555;
rom[66282] = 12'h444;
rom[66283] = 12'h333;
rom[66284] = 12'h111;
rom[66285] = 12'h111;
rom[66286] = 12'h111;
rom[66287] = 12'h111;
rom[66288] = 12'h111;
rom[66289] = 12'h111;
rom[66290] = 12'h111;
rom[66291] = 12'h111;
rom[66292] = 12'h111;
rom[66293] = 12'h111;
rom[66294] = 12'h111;
rom[66295] = 12'h111;
rom[66296] = 12'h111;
rom[66297] = 12'h222;
rom[66298] = 12'h222;
rom[66299] = 12'h333;
rom[66300] = 12'h333;
rom[66301] = 12'h333;
rom[66302] = 12'h333;
rom[66303] = 12'h333;
rom[66304] = 12'h333;
rom[66305] = 12'h444;
rom[66306] = 12'h444;
rom[66307] = 12'h444;
rom[66308] = 12'h444;
rom[66309] = 12'h444;
rom[66310] = 12'h555;
rom[66311] = 12'h555;
rom[66312] = 12'h555;
rom[66313] = 12'h666;
rom[66314] = 12'h777;
rom[66315] = 12'h777;
rom[66316] = 12'h888;
rom[66317] = 12'h888;
rom[66318] = 12'h888;
rom[66319] = 12'h999;
rom[66320] = 12'h888;
rom[66321] = 12'h888;
rom[66322] = 12'h888;
rom[66323] = 12'h999;
rom[66324] = 12'h999;
rom[66325] = 12'h999;
rom[66326] = 12'h999;
rom[66327] = 12'h999;
rom[66328] = 12'h999;
rom[66329] = 12'haaa;
rom[66330] = 12'haaa;
rom[66331] = 12'haaa;
rom[66332] = 12'haaa;
rom[66333] = 12'hbbb;
rom[66334] = 12'hbbb;
rom[66335] = 12'hbbb;
rom[66336] = 12'hbbb;
rom[66337] = 12'hccc;
rom[66338] = 12'hccc;
rom[66339] = 12'hccc;
rom[66340] = 12'hddd;
rom[66341] = 12'hddd;
rom[66342] = 12'heee;
rom[66343] = 12'heee;
rom[66344] = 12'hfff;
rom[66345] = 12'hfff;
rom[66346] = 12'hfff;
rom[66347] = 12'hfff;
rom[66348] = 12'hfff;
rom[66349] = 12'hfff;
rom[66350] = 12'heee;
rom[66351] = 12'heee;
rom[66352] = 12'hddd;
rom[66353] = 12'hddd;
rom[66354] = 12'hccc;
rom[66355] = 12'hccc;
rom[66356] = 12'hccc;
rom[66357] = 12'hccc;
rom[66358] = 12'hbbb;
rom[66359] = 12'hbbb;
rom[66360] = 12'hbbb;
rom[66361] = 12'hbbb;
rom[66362] = 12'haaa;
rom[66363] = 12'haaa;
rom[66364] = 12'haaa;
rom[66365] = 12'haaa;
rom[66366] = 12'haaa;
rom[66367] = 12'haaa;
rom[66368] = 12'h999;
rom[66369] = 12'h999;
rom[66370] = 12'h999;
rom[66371] = 12'h999;
rom[66372] = 12'h999;
rom[66373] = 12'h999;
rom[66374] = 12'h999;
rom[66375] = 12'h999;
rom[66376] = 12'haaa;
rom[66377] = 12'haaa;
rom[66378] = 12'hbbb;
rom[66379] = 12'hccc;
rom[66380] = 12'hccc;
rom[66381] = 12'hbbb;
rom[66382] = 12'haaa;
rom[66383] = 12'h999;
rom[66384] = 12'h888;
rom[66385] = 12'h888;
rom[66386] = 12'h777;
rom[66387] = 12'h777;
rom[66388] = 12'h777;
rom[66389] = 12'h777;
rom[66390] = 12'h777;
rom[66391] = 12'h777;
rom[66392] = 12'h777;
rom[66393] = 12'h777;
rom[66394] = 12'h777;
rom[66395] = 12'h777;
rom[66396] = 12'h666;
rom[66397] = 12'h666;
rom[66398] = 12'h777;
rom[66399] = 12'h777;
rom[66400] = 12'hfff;
rom[66401] = 12'hfff;
rom[66402] = 12'hfff;
rom[66403] = 12'hfff;
rom[66404] = 12'hfff;
rom[66405] = 12'hfff;
rom[66406] = 12'hfff;
rom[66407] = 12'hfff;
rom[66408] = 12'hfff;
rom[66409] = 12'hfff;
rom[66410] = 12'hfff;
rom[66411] = 12'hfff;
rom[66412] = 12'hfff;
rom[66413] = 12'hfff;
rom[66414] = 12'hfff;
rom[66415] = 12'hfff;
rom[66416] = 12'hfff;
rom[66417] = 12'hfff;
rom[66418] = 12'hfff;
rom[66419] = 12'hfff;
rom[66420] = 12'hfff;
rom[66421] = 12'hfff;
rom[66422] = 12'hfff;
rom[66423] = 12'hfff;
rom[66424] = 12'hfff;
rom[66425] = 12'hfff;
rom[66426] = 12'hfff;
rom[66427] = 12'hfff;
rom[66428] = 12'hfff;
rom[66429] = 12'hfff;
rom[66430] = 12'hfff;
rom[66431] = 12'hfff;
rom[66432] = 12'hfff;
rom[66433] = 12'hfff;
rom[66434] = 12'hfff;
rom[66435] = 12'hfff;
rom[66436] = 12'hfff;
rom[66437] = 12'hfff;
rom[66438] = 12'hfff;
rom[66439] = 12'hfff;
rom[66440] = 12'hfff;
rom[66441] = 12'hfff;
rom[66442] = 12'hfff;
rom[66443] = 12'hfff;
rom[66444] = 12'hfff;
rom[66445] = 12'hfff;
rom[66446] = 12'hfff;
rom[66447] = 12'hfff;
rom[66448] = 12'hfff;
rom[66449] = 12'hfff;
rom[66450] = 12'hfff;
rom[66451] = 12'hfff;
rom[66452] = 12'hfff;
rom[66453] = 12'hfff;
rom[66454] = 12'hfff;
rom[66455] = 12'hfff;
rom[66456] = 12'hfff;
rom[66457] = 12'hfff;
rom[66458] = 12'hfff;
rom[66459] = 12'hfff;
rom[66460] = 12'hfff;
rom[66461] = 12'hfff;
rom[66462] = 12'hfff;
rom[66463] = 12'hfff;
rom[66464] = 12'hfff;
rom[66465] = 12'hfff;
rom[66466] = 12'hfff;
rom[66467] = 12'hfff;
rom[66468] = 12'hfff;
rom[66469] = 12'hfff;
rom[66470] = 12'hfff;
rom[66471] = 12'hfff;
rom[66472] = 12'hfff;
rom[66473] = 12'hfff;
rom[66474] = 12'hfff;
rom[66475] = 12'hfff;
rom[66476] = 12'hfff;
rom[66477] = 12'hfff;
rom[66478] = 12'hfff;
rom[66479] = 12'hfff;
rom[66480] = 12'hfff;
rom[66481] = 12'hfff;
rom[66482] = 12'hfff;
rom[66483] = 12'hfff;
rom[66484] = 12'hfff;
rom[66485] = 12'hfff;
rom[66486] = 12'hfff;
rom[66487] = 12'hfff;
rom[66488] = 12'hfff;
rom[66489] = 12'hfff;
rom[66490] = 12'hfff;
rom[66491] = 12'hfff;
rom[66492] = 12'hfff;
rom[66493] = 12'hfff;
rom[66494] = 12'hfff;
rom[66495] = 12'hfff;
rom[66496] = 12'hfff;
rom[66497] = 12'hfff;
rom[66498] = 12'hfff;
rom[66499] = 12'hfff;
rom[66500] = 12'hfff;
rom[66501] = 12'hfff;
rom[66502] = 12'hfff;
rom[66503] = 12'hfff;
rom[66504] = 12'hfff;
rom[66505] = 12'hfff;
rom[66506] = 12'hfff;
rom[66507] = 12'hfff;
rom[66508] = 12'hfff;
rom[66509] = 12'hfff;
rom[66510] = 12'hfff;
rom[66511] = 12'heee;
rom[66512] = 12'heee;
rom[66513] = 12'heee;
rom[66514] = 12'hddd;
rom[66515] = 12'hddd;
rom[66516] = 12'hccc;
rom[66517] = 12'hccc;
rom[66518] = 12'hccc;
rom[66519] = 12'hccc;
rom[66520] = 12'hbbb;
rom[66521] = 12'hbbb;
rom[66522] = 12'haaa;
rom[66523] = 12'haaa;
rom[66524] = 12'haaa;
rom[66525] = 12'h999;
rom[66526] = 12'h999;
rom[66527] = 12'h999;
rom[66528] = 12'h888;
rom[66529] = 12'h888;
rom[66530] = 12'h888;
rom[66531] = 12'h888;
rom[66532] = 12'h888;
rom[66533] = 12'h888;
rom[66534] = 12'h888;
rom[66535] = 12'h888;
rom[66536] = 12'h999;
rom[66537] = 12'h999;
rom[66538] = 12'h888;
rom[66539] = 12'h888;
rom[66540] = 12'h888;
rom[66541] = 12'h777;
rom[66542] = 12'h777;
rom[66543] = 12'h777;
rom[66544] = 12'h666;
rom[66545] = 12'h666;
rom[66546] = 12'h555;
rom[66547] = 12'h555;
rom[66548] = 12'h555;
rom[66549] = 12'h555;
rom[66550] = 12'h555;
rom[66551] = 12'h555;
rom[66552] = 12'h555;
rom[66553] = 12'h444;
rom[66554] = 12'h444;
rom[66555] = 12'h444;
rom[66556] = 12'h444;
rom[66557] = 12'h333;
rom[66558] = 12'h333;
rom[66559] = 12'h333;
rom[66560] = 12'h333;
rom[66561] = 12'h333;
rom[66562] = 12'h333;
rom[66563] = 12'h222;
rom[66564] = 12'h222;
rom[66565] = 12'h222;
rom[66566] = 12'h222;
rom[66567] = 12'h222;
rom[66568] = 12'h222;
rom[66569] = 12'h222;
rom[66570] = 12'h111;
rom[66571] = 12'h111;
rom[66572] = 12'h111;
rom[66573] = 12'h111;
rom[66574] = 12'h111;
rom[66575] = 12'h111;
rom[66576] = 12'h111;
rom[66577] = 12'h111;
rom[66578] = 12'h111;
rom[66579] = 12'h111;
rom[66580] = 12'h111;
rom[66581] = 12'h111;
rom[66582] = 12'h111;
rom[66583] = 12'h111;
rom[66584] = 12'h111;
rom[66585] = 12'h111;
rom[66586] = 12'h111;
rom[66587] = 12'h111;
rom[66588] = 12'h111;
rom[66589] = 12'h111;
rom[66590] = 12'h111;
rom[66591] = 12'h  0;
rom[66592] = 12'h  0;
rom[66593] = 12'h  0;
rom[66594] = 12'h  0;
rom[66595] = 12'h  0;
rom[66596] = 12'h  0;
rom[66597] = 12'h  0;
rom[66598] = 12'h  0;
rom[66599] = 12'h  0;
rom[66600] = 12'h  0;
rom[66601] = 12'h  0;
rom[66602] = 12'h  0;
rom[66603] = 12'h  0;
rom[66604] = 12'h  0;
rom[66605] = 12'h  0;
rom[66606] = 12'h  0;
rom[66607] = 12'h111;
rom[66608] = 12'h111;
rom[66609] = 12'h111;
rom[66610] = 12'h111;
rom[66611] = 12'h111;
rom[66612] = 12'h111;
rom[66613] = 12'h111;
rom[66614] = 12'h111;
rom[66615] = 12'h111;
rom[66616] = 12'h  0;
rom[66617] = 12'h  0;
rom[66618] = 12'h111;
rom[66619] = 12'h111;
rom[66620] = 12'h111;
rom[66621] = 12'h  0;
rom[66622] = 12'h  0;
rom[66623] = 12'h  0;
rom[66624] = 12'h  0;
rom[66625] = 12'h  0;
rom[66626] = 12'h  0;
rom[66627] = 12'h  0;
rom[66628] = 12'h  0;
rom[66629] = 12'h  0;
rom[66630] = 12'h  0;
rom[66631] = 12'h  0;
rom[66632] = 12'h  0;
rom[66633] = 12'h  0;
rom[66634] = 12'h  0;
rom[66635] = 12'h  0;
rom[66636] = 12'h  0;
rom[66637] = 12'h  0;
rom[66638] = 12'h  0;
rom[66639] = 12'h  0;
rom[66640] = 12'h  0;
rom[66641] = 12'h  0;
rom[66642] = 12'h  0;
rom[66643] = 12'h  0;
rom[66644] = 12'h  0;
rom[66645] = 12'h  0;
rom[66646] = 12'h  0;
rom[66647] = 12'h  0;
rom[66648] = 12'h  0;
rom[66649] = 12'h  0;
rom[66650] = 12'h  0;
rom[66651] = 12'h  0;
rom[66652] = 12'h  0;
rom[66653] = 12'h  0;
rom[66654] = 12'h  0;
rom[66655] = 12'h  0;
rom[66656] = 12'h  0;
rom[66657] = 12'h  0;
rom[66658] = 12'h  0;
rom[66659] = 12'h  0;
rom[66660] = 12'h  0;
rom[66661] = 12'h  0;
rom[66662] = 12'h  0;
rom[66663] = 12'h  0;
rom[66664] = 12'h  0;
rom[66665] = 12'h  0;
rom[66666] = 12'h  0;
rom[66667] = 12'h  0;
rom[66668] = 12'h  0;
rom[66669] = 12'h  0;
rom[66670] = 12'h  0;
rom[66671] = 12'h  0;
rom[66672] = 12'h111;
rom[66673] = 12'h111;
rom[66674] = 12'h222;
rom[66675] = 12'h222;
rom[66676] = 12'h333;
rom[66677] = 12'h444;
rom[66678] = 12'h444;
rom[66679] = 12'h555;
rom[66680] = 12'h555;
rom[66681] = 12'h555;
rom[66682] = 12'h444;
rom[66683] = 12'h222;
rom[66684] = 12'h111;
rom[66685] = 12'h111;
rom[66686] = 12'h111;
rom[66687] = 12'h111;
rom[66688] = 12'h111;
rom[66689] = 12'h111;
rom[66690] = 12'h111;
rom[66691] = 12'h111;
rom[66692] = 12'h111;
rom[66693] = 12'h111;
rom[66694] = 12'h111;
rom[66695] = 12'h111;
rom[66696] = 12'h111;
rom[66697] = 12'h111;
rom[66698] = 12'h222;
rom[66699] = 12'h333;
rom[66700] = 12'h333;
rom[66701] = 12'h333;
rom[66702] = 12'h333;
rom[66703] = 12'h333;
rom[66704] = 12'h333;
rom[66705] = 12'h333;
rom[66706] = 12'h444;
rom[66707] = 12'h444;
rom[66708] = 12'h444;
rom[66709] = 12'h444;
rom[66710] = 12'h555;
rom[66711] = 12'h555;
rom[66712] = 12'h555;
rom[66713] = 12'h666;
rom[66714] = 12'h777;
rom[66715] = 12'h777;
rom[66716] = 12'h888;
rom[66717] = 12'h888;
rom[66718] = 12'h888;
rom[66719] = 12'h999;
rom[66720] = 12'h999;
rom[66721] = 12'h999;
rom[66722] = 12'h999;
rom[66723] = 12'h999;
rom[66724] = 12'h999;
rom[66725] = 12'h999;
rom[66726] = 12'h999;
rom[66727] = 12'h999;
rom[66728] = 12'haaa;
rom[66729] = 12'haaa;
rom[66730] = 12'haaa;
rom[66731] = 12'haaa;
rom[66732] = 12'hbbb;
rom[66733] = 12'hbbb;
rom[66734] = 12'hbbb;
rom[66735] = 12'hbbb;
rom[66736] = 12'hccc;
rom[66737] = 12'hccc;
rom[66738] = 12'hccc;
rom[66739] = 12'hddd;
rom[66740] = 12'hddd;
rom[66741] = 12'heee;
rom[66742] = 12'hfff;
rom[66743] = 12'hfff;
rom[66744] = 12'hfff;
rom[66745] = 12'hfff;
rom[66746] = 12'hfff;
rom[66747] = 12'hfff;
rom[66748] = 12'hfff;
rom[66749] = 12'hfff;
rom[66750] = 12'heee;
rom[66751] = 12'heee;
rom[66752] = 12'hddd;
rom[66753] = 12'hddd;
rom[66754] = 12'hccc;
rom[66755] = 12'hccc;
rom[66756] = 12'hbbb;
rom[66757] = 12'hbbb;
rom[66758] = 12'hbbb;
rom[66759] = 12'haaa;
rom[66760] = 12'haaa;
rom[66761] = 12'haaa;
rom[66762] = 12'haaa;
rom[66763] = 12'haaa;
rom[66764] = 12'h999;
rom[66765] = 12'h999;
rom[66766] = 12'h999;
rom[66767] = 12'h999;
rom[66768] = 12'h999;
rom[66769] = 12'h999;
rom[66770] = 12'h999;
rom[66771] = 12'h999;
rom[66772] = 12'h999;
rom[66773] = 12'h999;
rom[66774] = 12'h999;
rom[66775] = 12'h999;
rom[66776] = 12'h999;
rom[66777] = 12'haaa;
rom[66778] = 12'haaa;
rom[66779] = 12'hbbb;
rom[66780] = 12'hbbb;
rom[66781] = 12'hbbb;
rom[66782] = 12'hbbb;
rom[66783] = 12'haaa;
rom[66784] = 12'h999;
rom[66785] = 12'h888;
rom[66786] = 12'h888;
rom[66787] = 12'h777;
rom[66788] = 12'h777;
rom[66789] = 12'h777;
rom[66790] = 12'h777;
rom[66791] = 12'h777;
rom[66792] = 12'h777;
rom[66793] = 12'h777;
rom[66794] = 12'h777;
rom[66795] = 12'h666;
rom[66796] = 12'h666;
rom[66797] = 12'h666;
rom[66798] = 12'h666;
rom[66799] = 12'h666;
rom[66800] = 12'hfff;
rom[66801] = 12'hfff;
rom[66802] = 12'hfff;
rom[66803] = 12'hfff;
rom[66804] = 12'hfff;
rom[66805] = 12'hfff;
rom[66806] = 12'hfff;
rom[66807] = 12'hfff;
rom[66808] = 12'hfff;
rom[66809] = 12'hfff;
rom[66810] = 12'hfff;
rom[66811] = 12'hfff;
rom[66812] = 12'hfff;
rom[66813] = 12'hfff;
rom[66814] = 12'hfff;
rom[66815] = 12'hfff;
rom[66816] = 12'hfff;
rom[66817] = 12'hfff;
rom[66818] = 12'hfff;
rom[66819] = 12'hfff;
rom[66820] = 12'hfff;
rom[66821] = 12'hfff;
rom[66822] = 12'hfff;
rom[66823] = 12'hfff;
rom[66824] = 12'hfff;
rom[66825] = 12'hfff;
rom[66826] = 12'hfff;
rom[66827] = 12'hfff;
rom[66828] = 12'hfff;
rom[66829] = 12'hfff;
rom[66830] = 12'hfff;
rom[66831] = 12'hfff;
rom[66832] = 12'hfff;
rom[66833] = 12'hfff;
rom[66834] = 12'hfff;
rom[66835] = 12'hfff;
rom[66836] = 12'hfff;
rom[66837] = 12'hfff;
rom[66838] = 12'hfff;
rom[66839] = 12'hfff;
rom[66840] = 12'hfff;
rom[66841] = 12'hfff;
rom[66842] = 12'hfff;
rom[66843] = 12'hfff;
rom[66844] = 12'hfff;
rom[66845] = 12'hfff;
rom[66846] = 12'hfff;
rom[66847] = 12'hfff;
rom[66848] = 12'hfff;
rom[66849] = 12'hfff;
rom[66850] = 12'hfff;
rom[66851] = 12'hfff;
rom[66852] = 12'hfff;
rom[66853] = 12'hfff;
rom[66854] = 12'hfff;
rom[66855] = 12'hfff;
rom[66856] = 12'hfff;
rom[66857] = 12'hfff;
rom[66858] = 12'hfff;
rom[66859] = 12'hfff;
rom[66860] = 12'hfff;
rom[66861] = 12'hfff;
rom[66862] = 12'hfff;
rom[66863] = 12'hfff;
rom[66864] = 12'hfff;
rom[66865] = 12'hfff;
rom[66866] = 12'hfff;
rom[66867] = 12'hfff;
rom[66868] = 12'hfff;
rom[66869] = 12'hfff;
rom[66870] = 12'hfff;
rom[66871] = 12'hfff;
rom[66872] = 12'hfff;
rom[66873] = 12'hfff;
rom[66874] = 12'hfff;
rom[66875] = 12'hfff;
rom[66876] = 12'hfff;
rom[66877] = 12'hfff;
rom[66878] = 12'hfff;
rom[66879] = 12'hfff;
rom[66880] = 12'hfff;
rom[66881] = 12'hfff;
rom[66882] = 12'hfff;
rom[66883] = 12'hfff;
rom[66884] = 12'hfff;
rom[66885] = 12'hfff;
rom[66886] = 12'hfff;
rom[66887] = 12'hfff;
rom[66888] = 12'hfff;
rom[66889] = 12'hfff;
rom[66890] = 12'hfff;
rom[66891] = 12'hfff;
rom[66892] = 12'hfff;
rom[66893] = 12'hfff;
rom[66894] = 12'hfff;
rom[66895] = 12'hfff;
rom[66896] = 12'hfff;
rom[66897] = 12'hfff;
rom[66898] = 12'hfff;
rom[66899] = 12'hfff;
rom[66900] = 12'hfff;
rom[66901] = 12'hfff;
rom[66902] = 12'hfff;
rom[66903] = 12'hfff;
rom[66904] = 12'hfff;
rom[66905] = 12'hfff;
rom[66906] = 12'hfff;
rom[66907] = 12'hfff;
rom[66908] = 12'hfff;
rom[66909] = 12'hfff;
rom[66910] = 12'hfff;
rom[66911] = 12'heee;
rom[66912] = 12'heee;
rom[66913] = 12'heee;
rom[66914] = 12'hddd;
rom[66915] = 12'hddd;
rom[66916] = 12'hccc;
rom[66917] = 12'hccc;
rom[66918] = 12'hbbb;
rom[66919] = 12'hbbb;
rom[66920] = 12'hbbb;
rom[66921] = 12'hbbb;
rom[66922] = 12'hbbb;
rom[66923] = 12'haaa;
rom[66924] = 12'haaa;
rom[66925] = 12'h999;
rom[66926] = 12'h999;
rom[66927] = 12'h888;
rom[66928] = 12'h888;
rom[66929] = 12'h888;
rom[66930] = 12'h888;
rom[66931] = 12'h777;
rom[66932] = 12'h777;
rom[66933] = 12'h777;
rom[66934] = 12'h777;
rom[66935] = 12'h777;
rom[66936] = 12'h777;
rom[66937] = 12'h888;
rom[66938] = 12'h888;
rom[66939] = 12'h999;
rom[66940] = 12'h999;
rom[66941] = 12'h888;
rom[66942] = 12'h888;
rom[66943] = 12'h777;
rom[66944] = 12'h777;
rom[66945] = 12'h777;
rom[66946] = 12'h666;
rom[66947] = 12'h555;
rom[66948] = 12'h555;
rom[66949] = 12'h555;
rom[66950] = 12'h666;
rom[66951] = 12'h666;
rom[66952] = 12'h555;
rom[66953] = 12'h555;
rom[66954] = 12'h444;
rom[66955] = 12'h444;
rom[66956] = 12'h444;
rom[66957] = 12'h444;
rom[66958] = 12'h444;
rom[66959] = 12'h333;
rom[66960] = 12'h333;
rom[66961] = 12'h333;
rom[66962] = 12'h333;
rom[66963] = 12'h222;
rom[66964] = 12'h222;
rom[66965] = 12'h222;
rom[66966] = 12'h222;
rom[66967] = 12'h222;
rom[66968] = 12'h222;
rom[66969] = 12'h222;
rom[66970] = 12'h111;
rom[66971] = 12'h111;
rom[66972] = 12'h111;
rom[66973] = 12'h111;
rom[66974] = 12'h111;
rom[66975] = 12'h111;
rom[66976] = 12'h111;
rom[66977] = 12'h111;
rom[66978] = 12'h111;
rom[66979] = 12'h111;
rom[66980] = 12'h111;
rom[66981] = 12'h111;
rom[66982] = 12'h111;
rom[66983] = 12'h111;
rom[66984] = 12'h111;
rom[66985] = 12'h111;
rom[66986] = 12'h111;
rom[66987] = 12'h111;
rom[66988] = 12'h111;
rom[66989] = 12'h111;
rom[66990] = 12'h111;
rom[66991] = 12'h111;
rom[66992] = 12'h  0;
rom[66993] = 12'h  0;
rom[66994] = 12'h  0;
rom[66995] = 12'h  0;
rom[66996] = 12'h  0;
rom[66997] = 12'h  0;
rom[66998] = 12'h  0;
rom[66999] = 12'h  0;
rom[67000] = 12'h  0;
rom[67001] = 12'h  0;
rom[67002] = 12'h  0;
rom[67003] = 12'h  0;
rom[67004] = 12'h  0;
rom[67005] = 12'h  0;
rom[67006] = 12'h111;
rom[67007] = 12'h111;
rom[67008] = 12'h111;
rom[67009] = 12'h111;
rom[67010] = 12'h111;
rom[67011] = 12'h111;
rom[67012] = 12'h111;
rom[67013] = 12'h111;
rom[67014] = 12'h111;
rom[67015] = 12'h  0;
rom[67016] = 12'h  0;
rom[67017] = 12'h  0;
rom[67018] = 12'h111;
rom[67019] = 12'h111;
rom[67020] = 12'h111;
rom[67021] = 12'h  0;
rom[67022] = 12'h  0;
rom[67023] = 12'h  0;
rom[67024] = 12'h  0;
rom[67025] = 12'h  0;
rom[67026] = 12'h  0;
rom[67027] = 12'h  0;
rom[67028] = 12'h  0;
rom[67029] = 12'h  0;
rom[67030] = 12'h  0;
rom[67031] = 12'h  0;
rom[67032] = 12'h  0;
rom[67033] = 12'h  0;
rom[67034] = 12'h  0;
rom[67035] = 12'h  0;
rom[67036] = 12'h  0;
rom[67037] = 12'h  0;
rom[67038] = 12'h  0;
rom[67039] = 12'h  0;
rom[67040] = 12'h  0;
rom[67041] = 12'h  0;
rom[67042] = 12'h  0;
rom[67043] = 12'h  0;
rom[67044] = 12'h  0;
rom[67045] = 12'h  0;
rom[67046] = 12'h  0;
rom[67047] = 12'h  0;
rom[67048] = 12'h  0;
rom[67049] = 12'h  0;
rom[67050] = 12'h  0;
rom[67051] = 12'h  0;
rom[67052] = 12'h  0;
rom[67053] = 12'h  0;
rom[67054] = 12'h  0;
rom[67055] = 12'h  0;
rom[67056] = 12'h  0;
rom[67057] = 12'h  0;
rom[67058] = 12'h  0;
rom[67059] = 12'h  0;
rom[67060] = 12'h  0;
rom[67061] = 12'h  0;
rom[67062] = 12'h  0;
rom[67063] = 12'h  0;
rom[67064] = 12'h  0;
rom[67065] = 12'h  0;
rom[67066] = 12'h  0;
rom[67067] = 12'h  0;
rom[67068] = 12'h  0;
rom[67069] = 12'h  0;
rom[67070] = 12'h111;
rom[67071] = 12'h  0;
rom[67072] = 12'h111;
rom[67073] = 12'h111;
rom[67074] = 12'h222;
rom[67075] = 12'h222;
rom[67076] = 12'h333;
rom[67077] = 12'h444;
rom[67078] = 12'h444;
rom[67079] = 12'h444;
rom[67080] = 12'h555;
rom[67081] = 12'h555;
rom[67082] = 12'h444;
rom[67083] = 12'h222;
rom[67084] = 12'h111;
rom[67085] = 12'h111;
rom[67086] = 12'h111;
rom[67087] = 12'h111;
rom[67088] = 12'h111;
rom[67089] = 12'h111;
rom[67090] = 12'h111;
rom[67091] = 12'h111;
rom[67092] = 12'h111;
rom[67093] = 12'h111;
rom[67094] = 12'h111;
rom[67095] = 12'h111;
rom[67096] = 12'h111;
rom[67097] = 12'h111;
rom[67098] = 12'h222;
rom[67099] = 12'h333;
rom[67100] = 12'h333;
rom[67101] = 12'h333;
rom[67102] = 12'h333;
rom[67103] = 12'h333;
rom[67104] = 12'h333;
rom[67105] = 12'h333;
rom[67106] = 12'h444;
rom[67107] = 12'h444;
rom[67108] = 12'h444;
rom[67109] = 12'h555;
rom[67110] = 12'h555;
rom[67111] = 12'h555;
rom[67112] = 12'h555;
rom[67113] = 12'h666;
rom[67114] = 12'h777;
rom[67115] = 12'h777;
rom[67116] = 12'h888;
rom[67117] = 12'h888;
rom[67118] = 12'h999;
rom[67119] = 12'h999;
rom[67120] = 12'h999;
rom[67121] = 12'h999;
rom[67122] = 12'h999;
rom[67123] = 12'h999;
rom[67124] = 12'h999;
rom[67125] = 12'h999;
rom[67126] = 12'h999;
rom[67127] = 12'haaa;
rom[67128] = 12'haaa;
rom[67129] = 12'haaa;
rom[67130] = 12'haaa;
rom[67131] = 12'haaa;
rom[67132] = 12'hbbb;
rom[67133] = 12'hbbb;
rom[67134] = 12'hbbb;
rom[67135] = 12'hccc;
rom[67136] = 12'hccc;
rom[67137] = 12'hccc;
rom[67138] = 12'hddd;
rom[67139] = 12'hddd;
rom[67140] = 12'heee;
rom[67141] = 12'heee;
rom[67142] = 12'hfff;
rom[67143] = 12'hfff;
rom[67144] = 12'hfff;
rom[67145] = 12'hfff;
rom[67146] = 12'hfff;
rom[67147] = 12'hfff;
rom[67148] = 12'hfff;
rom[67149] = 12'heee;
rom[67150] = 12'heee;
rom[67151] = 12'hddd;
rom[67152] = 12'hddd;
rom[67153] = 12'hccc;
rom[67154] = 12'hccc;
rom[67155] = 12'hbbb;
rom[67156] = 12'hbbb;
rom[67157] = 12'hbbb;
rom[67158] = 12'haaa;
rom[67159] = 12'haaa;
rom[67160] = 12'haaa;
rom[67161] = 12'haaa;
rom[67162] = 12'haaa;
rom[67163] = 12'h999;
rom[67164] = 12'h999;
rom[67165] = 12'h999;
rom[67166] = 12'h999;
rom[67167] = 12'h999;
rom[67168] = 12'h999;
rom[67169] = 12'h999;
rom[67170] = 12'h999;
rom[67171] = 12'h999;
rom[67172] = 12'h999;
rom[67173] = 12'h999;
rom[67174] = 12'h888;
rom[67175] = 12'h888;
rom[67176] = 12'h888;
rom[67177] = 12'h999;
rom[67178] = 12'haaa;
rom[67179] = 12'hbbb;
rom[67180] = 12'hbbb;
rom[67181] = 12'hbbb;
rom[67182] = 12'hbbb;
rom[67183] = 12'hbbb;
rom[67184] = 12'haaa;
rom[67185] = 12'h999;
rom[67186] = 12'h888;
rom[67187] = 12'h777;
rom[67188] = 12'h777;
rom[67189] = 12'h777;
rom[67190] = 12'h777;
rom[67191] = 12'h777;
rom[67192] = 12'h777;
rom[67193] = 12'h777;
rom[67194] = 12'h666;
rom[67195] = 12'h666;
rom[67196] = 12'h666;
rom[67197] = 12'h666;
rom[67198] = 12'h666;
rom[67199] = 12'h666;
rom[67200] = 12'hfff;
rom[67201] = 12'hfff;
rom[67202] = 12'hfff;
rom[67203] = 12'hfff;
rom[67204] = 12'hfff;
rom[67205] = 12'hfff;
rom[67206] = 12'hfff;
rom[67207] = 12'hfff;
rom[67208] = 12'hfff;
rom[67209] = 12'hfff;
rom[67210] = 12'hfff;
rom[67211] = 12'hfff;
rom[67212] = 12'hfff;
rom[67213] = 12'hfff;
rom[67214] = 12'hfff;
rom[67215] = 12'hfff;
rom[67216] = 12'hfff;
rom[67217] = 12'hfff;
rom[67218] = 12'hfff;
rom[67219] = 12'hfff;
rom[67220] = 12'hfff;
rom[67221] = 12'hfff;
rom[67222] = 12'hfff;
rom[67223] = 12'hfff;
rom[67224] = 12'hfff;
rom[67225] = 12'hfff;
rom[67226] = 12'hfff;
rom[67227] = 12'hfff;
rom[67228] = 12'hfff;
rom[67229] = 12'hfff;
rom[67230] = 12'hfff;
rom[67231] = 12'hfff;
rom[67232] = 12'hfff;
rom[67233] = 12'hfff;
rom[67234] = 12'hfff;
rom[67235] = 12'hfff;
rom[67236] = 12'hfff;
rom[67237] = 12'hfff;
rom[67238] = 12'hfff;
rom[67239] = 12'hfff;
rom[67240] = 12'hfff;
rom[67241] = 12'hfff;
rom[67242] = 12'hfff;
rom[67243] = 12'hfff;
rom[67244] = 12'hfff;
rom[67245] = 12'hfff;
rom[67246] = 12'hfff;
rom[67247] = 12'hfff;
rom[67248] = 12'hfff;
rom[67249] = 12'hfff;
rom[67250] = 12'hfff;
rom[67251] = 12'hfff;
rom[67252] = 12'hfff;
rom[67253] = 12'hfff;
rom[67254] = 12'hfff;
rom[67255] = 12'hfff;
rom[67256] = 12'hfff;
rom[67257] = 12'hfff;
rom[67258] = 12'hfff;
rom[67259] = 12'hfff;
rom[67260] = 12'hfff;
rom[67261] = 12'hfff;
rom[67262] = 12'hfff;
rom[67263] = 12'hfff;
rom[67264] = 12'hfff;
rom[67265] = 12'hfff;
rom[67266] = 12'hfff;
rom[67267] = 12'hfff;
rom[67268] = 12'hfff;
rom[67269] = 12'hfff;
rom[67270] = 12'hfff;
rom[67271] = 12'hfff;
rom[67272] = 12'hfff;
rom[67273] = 12'hfff;
rom[67274] = 12'hfff;
rom[67275] = 12'hfff;
rom[67276] = 12'hfff;
rom[67277] = 12'hfff;
rom[67278] = 12'hfff;
rom[67279] = 12'hfff;
rom[67280] = 12'hfff;
rom[67281] = 12'hfff;
rom[67282] = 12'hfff;
rom[67283] = 12'hfff;
rom[67284] = 12'hfff;
rom[67285] = 12'hfff;
rom[67286] = 12'hfff;
rom[67287] = 12'hfff;
rom[67288] = 12'hfff;
rom[67289] = 12'hfff;
rom[67290] = 12'hfff;
rom[67291] = 12'hfff;
rom[67292] = 12'hfff;
rom[67293] = 12'hfff;
rom[67294] = 12'hfff;
rom[67295] = 12'hfff;
rom[67296] = 12'hfff;
rom[67297] = 12'hfff;
rom[67298] = 12'hfff;
rom[67299] = 12'hfff;
rom[67300] = 12'hfff;
rom[67301] = 12'hfff;
rom[67302] = 12'hfff;
rom[67303] = 12'hfff;
rom[67304] = 12'hfff;
rom[67305] = 12'hfff;
rom[67306] = 12'hfff;
rom[67307] = 12'hfff;
rom[67308] = 12'hfff;
rom[67309] = 12'hfff;
rom[67310] = 12'heee;
rom[67311] = 12'heee;
rom[67312] = 12'heee;
rom[67313] = 12'hddd;
rom[67314] = 12'hddd;
rom[67315] = 12'hccc;
rom[67316] = 12'hccc;
rom[67317] = 12'hbbb;
rom[67318] = 12'hbbb;
rom[67319] = 12'hbbb;
rom[67320] = 12'hbbb;
rom[67321] = 12'haaa;
rom[67322] = 12'haaa;
rom[67323] = 12'haaa;
rom[67324] = 12'h999;
rom[67325] = 12'h999;
rom[67326] = 12'h999;
rom[67327] = 12'h999;
rom[67328] = 12'h888;
rom[67329] = 12'h888;
rom[67330] = 12'h777;
rom[67331] = 12'h777;
rom[67332] = 12'h777;
rom[67333] = 12'h777;
rom[67334] = 12'h777;
rom[67335] = 12'h777;
rom[67336] = 12'h777;
rom[67337] = 12'h777;
rom[67338] = 12'h777;
rom[67339] = 12'h777;
rom[67340] = 12'h777;
rom[67341] = 12'h777;
rom[67342] = 12'h777;
rom[67343] = 12'h777;
rom[67344] = 12'h777;
rom[67345] = 12'h777;
rom[67346] = 12'h777;
rom[67347] = 12'h777;
rom[67348] = 12'h777;
rom[67349] = 12'h666;
rom[67350] = 12'h666;
rom[67351] = 12'h666;
rom[67352] = 12'h555;
rom[67353] = 12'h555;
rom[67354] = 12'h555;
rom[67355] = 12'h555;
rom[67356] = 12'h444;
rom[67357] = 12'h444;
rom[67358] = 12'h444;
rom[67359] = 12'h444;
rom[67360] = 12'h444;
rom[67361] = 12'h333;
rom[67362] = 12'h333;
rom[67363] = 12'h333;
rom[67364] = 12'h333;
rom[67365] = 12'h333;
rom[67366] = 12'h222;
rom[67367] = 12'h222;
rom[67368] = 12'h222;
rom[67369] = 12'h222;
rom[67370] = 12'h222;
rom[67371] = 12'h222;
rom[67372] = 12'h222;
rom[67373] = 12'h222;
rom[67374] = 12'h111;
rom[67375] = 12'h111;
rom[67376] = 12'h111;
rom[67377] = 12'h111;
rom[67378] = 12'h111;
rom[67379] = 12'h111;
rom[67380] = 12'h111;
rom[67381] = 12'h111;
rom[67382] = 12'h111;
rom[67383] = 12'h111;
rom[67384] = 12'h111;
rom[67385] = 12'h111;
rom[67386] = 12'h111;
rom[67387] = 12'h111;
rom[67388] = 12'h111;
rom[67389] = 12'h111;
rom[67390] = 12'h111;
rom[67391] = 12'h111;
rom[67392] = 12'h  0;
rom[67393] = 12'h  0;
rom[67394] = 12'h  0;
rom[67395] = 12'h  0;
rom[67396] = 12'h  0;
rom[67397] = 12'h  0;
rom[67398] = 12'h  0;
rom[67399] = 12'h  0;
rom[67400] = 12'h  0;
rom[67401] = 12'h  0;
rom[67402] = 12'h  0;
rom[67403] = 12'h  0;
rom[67404] = 12'h  0;
rom[67405] = 12'h111;
rom[67406] = 12'h111;
rom[67407] = 12'h  0;
rom[67408] = 12'h111;
rom[67409] = 12'h111;
rom[67410] = 12'h111;
rom[67411] = 12'h111;
rom[67412] = 12'h111;
rom[67413] = 12'h111;
rom[67414] = 12'h111;
rom[67415] = 12'h  0;
rom[67416] = 12'h  0;
rom[67417] = 12'h  0;
rom[67418] = 12'h111;
rom[67419] = 12'h111;
rom[67420] = 12'h  0;
rom[67421] = 12'h  0;
rom[67422] = 12'h  0;
rom[67423] = 12'h  0;
rom[67424] = 12'h  0;
rom[67425] = 12'h  0;
rom[67426] = 12'h  0;
rom[67427] = 12'h  0;
rom[67428] = 12'h  0;
rom[67429] = 12'h  0;
rom[67430] = 12'h  0;
rom[67431] = 12'h  0;
rom[67432] = 12'h  0;
rom[67433] = 12'h  0;
rom[67434] = 12'h  0;
rom[67435] = 12'h  0;
rom[67436] = 12'h  0;
rom[67437] = 12'h  0;
rom[67438] = 12'h  0;
rom[67439] = 12'h  0;
rom[67440] = 12'h  0;
rom[67441] = 12'h  0;
rom[67442] = 12'h  0;
rom[67443] = 12'h  0;
rom[67444] = 12'h  0;
rom[67445] = 12'h  0;
rom[67446] = 12'h  0;
rom[67447] = 12'h  0;
rom[67448] = 12'h  0;
rom[67449] = 12'h  0;
rom[67450] = 12'h  0;
rom[67451] = 12'h  0;
rom[67452] = 12'h  0;
rom[67453] = 12'h  0;
rom[67454] = 12'h  0;
rom[67455] = 12'h  0;
rom[67456] = 12'h  0;
rom[67457] = 12'h  0;
rom[67458] = 12'h  0;
rom[67459] = 12'h  0;
rom[67460] = 12'h  0;
rom[67461] = 12'h  0;
rom[67462] = 12'h  0;
rom[67463] = 12'h  0;
rom[67464] = 12'h  0;
rom[67465] = 12'h  0;
rom[67466] = 12'h  0;
rom[67467] = 12'h  0;
rom[67468] = 12'h  0;
rom[67469] = 12'h  0;
rom[67470] = 12'h  0;
rom[67471] = 12'h  0;
rom[67472] = 12'h111;
rom[67473] = 12'h111;
rom[67474] = 12'h222;
rom[67475] = 12'h333;
rom[67476] = 12'h333;
rom[67477] = 12'h444;
rom[67478] = 12'h444;
rom[67479] = 12'h555;
rom[67480] = 12'h555;
rom[67481] = 12'h555;
rom[67482] = 12'h444;
rom[67483] = 12'h222;
rom[67484] = 12'h111;
rom[67485] = 12'h111;
rom[67486] = 12'h111;
rom[67487] = 12'h  0;
rom[67488] = 12'h111;
rom[67489] = 12'h111;
rom[67490] = 12'h111;
rom[67491] = 12'h111;
rom[67492] = 12'h111;
rom[67493] = 12'h111;
rom[67494] = 12'h111;
rom[67495] = 12'h111;
rom[67496] = 12'h111;
rom[67497] = 12'h111;
rom[67498] = 12'h111;
rom[67499] = 12'h222;
rom[67500] = 12'h333;
rom[67501] = 12'h333;
rom[67502] = 12'h333;
rom[67503] = 12'h333;
rom[67504] = 12'h333;
rom[67505] = 12'h333;
rom[67506] = 12'h444;
rom[67507] = 12'h444;
rom[67508] = 12'h555;
rom[67509] = 12'h555;
rom[67510] = 12'h555;
rom[67511] = 12'h444;
rom[67512] = 12'h555;
rom[67513] = 12'h666;
rom[67514] = 12'h777;
rom[67515] = 12'h888;
rom[67516] = 12'h888;
rom[67517] = 12'h999;
rom[67518] = 12'h999;
rom[67519] = 12'h999;
rom[67520] = 12'h999;
rom[67521] = 12'h999;
rom[67522] = 12'h999;
rom[67523] = 12'h999;
rom[67524] = 12'h999;
rom[67525] = 12'h999;
rom[67526] = 12'haaa;
rom[67527] = 12'haaa;
rom[67528] = 12'haaa;
rom[67529] = 12'haaa;
rom[67530] = 12'haaa;
rom[67531] = 12'hbbb;
rom[67532] = 12'hbbb;
rom[67533] = 12'hccc;
rom[67534] = 12'hccc;
rom[67535] = 12'hccc;
rom[67536] = 12'hccc;
rom[67537] = 12'hddd;
rom[67538] = 12'hddd;
rom[67539] = 12'heee;
rom[67540] = 12'heee;
rom[67541] = 12'hfff;
rom[67542] = 12'hfff;
rom[67543] = 12'hfff;
rom[67544] = 12'hfff;
rom[67545] = 12'hfff;
rom[67546] = 12'hfff;
rom[67547] = 12'hfff;
rom[67548] = 12'hfff;
rom[67549] = 12'heee;
rom[67550] = 12'hddd;
rom[67551] = 12'hddd;
rom[67552] = 12'hccc;
rom[67553] = 12'hccc;
rom[67554] = 12'hbbb;
rom[67555] = 12'hbbb;
rom[67556] = 12'haaa;
rom[67557] = 12'haaa;
rom[67558] = 12'haaa;
rom[67559] = 12'h999;
rom[67560] = 12'h999;
rom[67561] = 12'h999;
rom[67562] = 12'h999;
rom[67563] = 12'h999;
rom[67564] = 12'h999;
rom[67565] = 12'h888;
rom[67566] = 12'h888;
rom[67567] = 12'h888;
rom[67568] = 12'h888;
rom[67569] = 12'h888;
rom[67570] = 12'h888;
rom[67571] = 12'h888;
rom[67572] = 12'h888;
rom[67573] = 12'h888;
rom[67574] = 12'h888;
rom[67575] = 12'h888;
rom[67576] = 12'h888;
rom[67577] = 12'h888;
rom[67578] = 12'h999;
rom[67579] = 12'h999;
rom[67580] = 12'haaa;
rom[67581] = 12'hbbb;
rom[67582] = 12'hbbb;
rom[67583] = 12'hbbb;
rom[67584] = 12'hbbb;
rom[67585] = 12'haaa;
rom[67586] = 12'h999;
rom[67587] = 12'h888;
rom[67588] = 12'h777;
rom[67589] = 12'h777;
rom[67590] = 12'h777;
rom[67591] = 12'h666;
rom[67592] = 12'h777;
rom[67593] = 12'h666;
rom[67594] = 12'h666;
rom[67595] = 12'h666;
rom[67596] = 12'h666;
rom[67597] = 12'h666;
rom[67598] = 12'h666;
rom[67599] = 12'h666;
rom[67600] = 12'hfff;
rom[67601] = 12'hfff;
rom[67602] = 12'hfff;
rom[67603] = 12'hfff;
rom[67604] = 12'hfff;
rom[67605] = 12'hfff;
rom[67606] = 12'hfff;
rom[67607] = 12'hfff;
rom[67608] = 12'hfff;
rom[67609] = 12'hfff;
rom[67610] = 12'hfff;
rom[67611] = 12'hfff;
rom[67612] = 12'hfff;
rom[67613] = 12'hfff;
rom[67614] = 12'hfff;
rom[67615] = 12'hfff;
rom[67616] = 12'hfff;
rom[67617] = 12'hfff;
rom[67618] = 12'hfff;
rom[67619] = 12'hfff;
rom[67620] = 12'hfff;
rom[67621] = 12'hfff;
rom[67622] = 12'hfff;
rom[67623] = 12'hfff;
rom[67624] = 12'hfff;
rom[67625] = 12'hfff;
rom[67626] = 12'hfff;
rom[67627] = 12'hfff;
rom[67628] = 12'hfff;
rom[67629] = 12'hfff;
rom[67630] = 12'hfff;
rom[67631] = 12'hfff;
rom[67632] = 12'hfff;
rom[67633] = 12'hfff;
rom[67634] = 12'hfff;
rom[67635] = 12'hfff;
rom[67636] = 12'hfff;
rom[67637] = 12'hfff;
rom[67638] = 12'hfff;
rom[67639] = 12'hfff;
rom[67640] = 12'hfff;
rom[67641] = 12'hfff;
rom[67642] = 12'hfff;
rom[67643] = 12'hfff;
rom[67644] = 12'hfff;
rom[67645] = 12'hfff;
rom[67646] = 12'hfff;
rom[67647] = 12'hfff;
rom[67648] = 12'hfff;
rom[67649] = 12'hfff;
rom[67650] = 12'hfff;
rom[67651] = 12'hfff;
rom[67652] = 12'hfff;
rom[67653] = 12'hfff;
rom[67654] = 12'hfff;
rom[67655] = 12'hfff;
rom[67656] = 12'hfff;
rom[67657] = 12'hfff;
rom[67658] = 12'hfff;
rom[67659] = 12'hfff;
rom[67660] = 12'hfff;
rom[67661] = 12'hfff;
rom[67662] = 12'hfff;
rom[67663] = 12'hfff;
rom[67664] = 12'hfff;
rom[67665] = 12'hfff;
rom[67666] = 12'hfff;
rom[67667] = 12'hfff;
rom[67668] = 12'hfff;
rom[67669] = 12'hfff;
rom[67670] = 12'hfff;
rom[67671] = 12'hfff;
rom[67672] = 12'hfff;
rom[67673] = 12'hfff;
rom[67674] = 12'hfff;
rom[67675] = 12'hfff;
rom[67676] = 12'hfff;
rom[67677] = 12'hfff;
rom[67678] = 12'hfff;
rom[67679] = 12'hfff;
rom[67680] = 12'hfff;
rom[67681] = 12'hfff;
rom[67682] = 12'hfff;
rom[67683] = 12'hfff;
rom[67684] = 12'hfff;
rom[67685] = 12'hfff;
rom[67686] = 12'hfff;
rom[67687] = 12'hfff;
rom[67688] = 12'hfff;
rom[67689] = 12'hfff;
rom[67690] = 12'hfff;
rom[67691] = 12'hfff;
rom[67692] = 12'hfff;
rom[67693] = 12'hfff;
rom[67694] = 12'hfff;
rom[67695] = 12'hfff;
rom[67696] = 12'hfff;
rom[67697] = 12'hfff;
rom[67698] = 12'hfff;
rom[67699] = 12'hfff;
rom[67700] = 12'hfff;
rom[67701] = 12'hfff;
rom[67702] = 12'hfff;
rom[67703] = 12'hfff;
rom[67704] = 12'hfff;
rom[67705] = 12'hfff;
rom[67706] = 12'hfff;
rom[67707] = 12'hfff;
rom[67708] = 12'hfff;
rom[67709] = 12'hfff;
rom[67710] = 12'heee;
rom[67711] = 12'heee;
rom[67712] = 12'heee;
rom[67713] = 12'hddd;
rom[67714] = 12'hddd;
rom[67715] = 12'hccc;
rom[67716] = 12'hccc;
rom[67717] = 12'hbbb;
rom[67718] = 12'hbbb;
rom[67719] = 12'hbbb;
rom[67720] = 12'haaa;
rom[67721] = 12'haaa;
rom[67722] = 12'h999;
rom[67723] = 12'h999;
rom[67724] = 12'h999;
rom[67725] = 12'h888;
rom[67726] = 12'h888;
rom[67727] = 12'h888;
rom[67728] = 12'h888;
rom[67729] = 12'h888;
rom[67730] = 12'h777;
rom[67731] = 12'h777;
rom[67732] = 12'h777;
rom[67733] = 12'h777;
rom[67734] = 12'h777;
rom[67735] = 12'h777;
rom[67736] = 12'h666;
rom[67737] = 12'h666;
rom[67738] = 12'h666;
rom[67739] = 12'h666;
rom[67740] = 12'h666;
rom[67741] = 12'h666;
rom[67742] = 12'h666;
rom[67743] = 12'h666;
rom[67744] = 12'h777;
rom[67745] = 12'h777;
rom[67746] = 12'h777;
rom[67747] = 12'h777;
rom[67748] = 12'h777;
rom[67749] = 12'h666;
rom[67750] = 12'h666;
rom[67751] = 12'h666;
rom[67752] = 12'h666;
rom[67753] = 12'h666;
rom[67754] = 12'h666;
rom[67755] = 12'h555;
rom[67756] = 12'h555;
rom[67757] = 12'h444;
rom[67758] = 12'h444;
rom[67759] = 12'h444;
rom[67760] = 12'h444;
rom[67761] = 12'h444;
rom[67762] = 12'h333;
rom[67763] = 12'h333;
rom[67764] = 12'h333;
rom[67765] = 12'h333;
rom[67766] = 12'h222;
rom[67767] = 12'h222;
rom[67768] = 12'h222;
rom[67769] = 12'h222;
rom[67770] = 12'h222;
rom[67771] = 12'h222;
rom[67772] = 12'h222;
rom[67773] = 12'h222;
rom[67774] = 12'h222;
rom[67775] = 12'h111;
rom[67776] = 12'h111;
rom[67777] = 12'h111;
rom[67778] = 12'h111;
rom[67779] = 12'h111;
rom[67780] = 12'h111;
rom[67781] = 12'h111;
rom[67782] = 12'h111;
rom[67783] = 12'h111;
rom[67784] = 12'h111;
rom[67785] = 12'h111;
rom[67786] = 12'h111;
rom[67787] = 12'h111;
rom[67788] = 12'h111;
rom[67789] = 12'h111;
rom[67790] = 12'h111;
rom[67791] = 12'h111;
rom[67792] = 12'h111;
rom[67793] = 12'h111;
rom[67794] = 12'h111;
rom[67795] = 12'h  0;
rom[67796] = 12'h  0;
rom[67797] = 12'h  0;
rom[67798] = 12'h  0;
rom[67799] = 12'h  0;
rom[67800] = 12'h  0;
rom[67801] = 12'h  0;
rom[67802] = 12'h  0;
rom[67803] = 12'h  0;
rom[67804] = 12'h111;
rom[67805] = 12'h111;
rom[67806] = 12'h111;
rom[67807] = 12'h  0;
rom[67808] = 12'h111;
rom[67809] = 12'h111;
rom[67810] = 12'h111;
rom[67811] = 12'h111;
rom[67812] = 12'h111;
rom[67813] = 12'h111;
rom[67814] = 12'h111;
rom[67815] = 12'h  0;
rom[67816] = 12'h  0;
rom[67817] = 12'h111;
rom[67818] = 12'h111;
rom[67819] = 12'h111;
rom[67820] = 12'h  0;
rom[67821] = 12'h  0;
rom[67822] = 12'h  0;
rom[67823] = 12'h  0;
rom[67824] = 12'h  0;
rom[67825] = 12'h  0;
rom[67826] = 12'h  0;
rom[67827] = 12'h  0;
rom[67828] = 12'h  0;
rom[67829] = 12'h  0;
rom[67830] = 12'h  0;
rom[67831] = 12'h  0;
rom[67832] = 12'h  0;
rom[67833] = 12'h  0;
rom[67834] = 12'h  0;
rom[67835] = 12'h  0;
rom[67836] = 12'h  0;
rom[67837] = 12'h  0;
rom[67838] = 12'h  0;
rom[67839] = 12'h  0;
rom[67840] = 12'h  0;
rom[67841] = 12'h  0;
rom[67842] = 12'h  0;
rom[67843] = 12'h  0;
rom[67844] = 12'h  0;
rom[67845] = 12'h  0;
rom[67846] = 12'h  0;
rom[67847] = 12'h  0;
rom[67848] = 12'h  0;
rom[67849] = 12'h  0;
rom[67850] = 12'h  0;
rom[67851] = 12'h  0;
rom[67852] = 12'h  0;
rom[67853] = 12'h  0;
rom[67854] = 12'h  0;
rom[67855] = 12'h  0;
rom[67856] = 12'h  0;
rom[67857] = 12'h  0;
rom[67858] = 12'h  0;
rom[67859] = 12'h  0;
rom[67860] = 12'h  0;
rom[67861] = 12'h  0;
rom[67862] = 12'h  0;
rom[67863] = 12'h  0;
rom[67864] = 12'h  0;
rom[67865] = 12'h  0;
rom[67866] = 12'h  0;
rom[67867] = 12'h  0;
rom[67868] = 12'h  0;
rom[67869] = 12'h  0;
rom[67870] = 12'h  0;
rom[67871] = 12'h111;
rom[67872] = 12'h111;
rom[67873] = 12'h111;
rom[67874] = 12'h222;
rom[67875] = 12'h333;
rom[67876] = 12'h333;
rom[67877] = 12'h444;
rom[67878] = 12'h444;
rom[67879] = 12'h555;
rom[67880] = 12'h555;
rom[67881] = 12'h555;
rom[67882] = 12'h444;
rom[67883] = 12'h222;
rom[67884] = 12'h111;
rom[67885] = 12'h111;
rom[67886] = 12'h111;
rom[67887] = 12'h111;
rom[67888] = 12'h111;
rom[67889] = 12'h111;
rom[67890] = 12'h111;
rom[67891] = 12'h111;
rom[67892] = 12'h111;
rom[67893] = 12'h111;
rom[67894] = 12'h111;
rom[67895] = 12'h111;
rom[67896] = 12'h111;
rom[67897] = 12'h111;
rom[67898] = 12'h111;
rom[67899] = 12'h222;
rom[67900] = 12'h333;
rom[67901] = 12'h333;
rom[67902] = 12'h333;
rom[67903] = 12'h333;
rom[67904] = 12'h333;
rom[67905] = 12'h333;
rom[67906] = 12'h333;
rom[67907] = 12'h444;
rom[67908] = 12'h555;
rom[67909] = 12'h555;
rom[67910] = 12'h555;
rom[67911] = 12'h555;
rom[67912] = 12'h555;
rom[67913] = 12'h666;
rom[67914] = 12'h777;
rom[67915] = 12'h777;
rom[67916] = 12'h888;
rom[67917] = 12'h999;
rom[67918] = 12'h999;
rom[67919] = 12'h999;
rom[67920] = 12'h999;
rom[67921] = 12'h999;
rom[67922] = 12'h999;
rom[67923] = 12'h999;
rom[67924] = 12'haaa;
rom[67925] = 12'haaa;
rom[67926] = 12'haaa;
rom[67927] = 12'haaa;
rom[67928] = 12'haaa;
rom[67929] = 12'haaa;
rom[67930] = 12'hbbb;
rom[67931] = 12'hbbb;
rom[67932] = 12'hbbb;
rom[67933] = 12'hccc;
rom[67934] = 12'hccc;
rom[67935] = 12'hccc;
rom[67936] = 12'hccc;
rom[67937] = 12'hddd;
rom[67938] = 12'heee;
rom[67939] = 12'heee;
rom[67940] = 12'hfff;
rom[67941] = 12'hfff;
rom[67942] = 12'hfff;
rom[67943] = 12'hfff;
rom[67944] = 12'hfff;
rom[67945] = 12'hfff;
rom[67946] = 12'hfff;
rom[67947] = 12'hfff;
rom[67948] = 12'heee;
rom[67949] = 12'heee;
rom[67950] = 12'hddd;
rom[67951] = 12'hccc;
rom[67952] = 12'hbbb;
rom[67953] = 12'hbbb;
rom[67954] = 12'hbbb;
rom[67955] = 12'haaa;
rom[67956] = 12'haaa;
rom[67957] = 12'haaa;
rom[67958] = 12'h999;
rom[67959] = 12'h999;
rom[67960] = 12'h999;
rom[67961] = 12'h999;
rom[67962] = 12'h999;
rom[67963] = 12'h999;
rom[67964] = 12'h888;
rom[67965] = 12'h888;
rom[67966] = 12'h888;
rom[67967] = 12'h888;
rom[67968] = 12'h777;
rom[67969] = 12'h777;
rom[67970] = 12'h777;
rom[67971] = 12'h777;
rom[67972] = 12'h777;
rom[67973] = 12'h777;
rom[67974] = 12'h888;
rom[67975] = 12'h888;
rom[67976] = 12'h888;
rom[67977] = 12'h888;
rom[67978] = 12'h888;
rom[67979] = 12'h999;
rom[67980] = 12'h999;
rom[67981] = 12'haaa;
rom[67982] = 12'haaa;
rom[67983] = 12'hbbb;
rom[67984] = 12'hbbb;
rom[67985] = 12'hbbb;
rom[67986] = 12'haaa;
rom[67987] = 12'h999;
rom[67988] = 12'h888;
rom[67989] = 12'h777;
rom[67990] = 12'h777;
rom[67991] = 12'h666;
rom[67992] = 12'h666;
rom[67993] = 12'h666;
rom[67994] = 12'h666;
rom[67995] = 12'h666;
rom[67996] = 12'h666;
rom[67997] = 12'h666;
rom[67998] = 12'h666;
rom[67999] = 12'h666;
rom[68000] = 12'hfff;
rom[68001] = 12'hfff;
rom[68002] = 12'hfff;
rom[68003] = 12'hfff;
rom[68004] = 12'hfff;
rom[68005] = 12'hfff;
rom[68006] = 12'hfff;
rom[68007] = 12'hfff;
rom[68008] = 12'hfff;
rom[68009] = 12'hfff;
rom[68010] = 12'hfff;
rom[68011] = 12'hfff;
rom[68012] = 12'hfff;
rom[68013] = 12'hfff;
rom[68014] = 12'hfff;
rom[68015] = 12'hfff;
rom[68016] = 12'hfff;
rom[68017] = 12'hfff;
rom[68018] = 12'hfff;
rom[68019] = 12'hfff;
rom[68020] = 12'hfff;
rom[68021] = 12'hfff;
rom[68022] = 12'hfff;
rom[68023] = 12'hfff;
rom[68024] = 12'hfff;
rom[68025] = 12'hfff;
rom[68026] = 12'hfff;
rom[68027] = 12'hfff;
rom[68028] = 12'hfff;
rom[68029] = 12'hfff;
rom[68030] = 12'hfff;
rom[68031] = 12'hfff;
rom[68032] = 12'hfff;
rom[68033] = 12'hfff;
rom[68034] = 12'hfff;
rom[68035] = 12'hfff;
rom[68036] = 12'hfff;
rom[68037] = 12'hfff;
rom[68038] = 12'hfff;
rom[68039] = 12'hfff;
rom[68040] = 12'hfff;
rom[68041] = 12'hfff;
rom[68042] = 12'hfff;
rom[68043] = 12'hfff;
rom[68044] = 12'hfff;
rom[68045] = 12'hfff;
rom[68046] = 12'hfff;
rom[68047] = 12'hfff;
rom[68048] = 12'hfff;
rom[68049] = 12'hfff;
rom[68050] = 12'hfff;
rom[68051] = 12'hfff;
rom[68052] = 12'hfff;
rom[68053] = 12'hfff;
rom[68054] = 12'hfff;
rom[68055] = 12'hfff;
rom[68056] = 12'hfff;
rom[68057] = 12'hfff;
rom[68058] = 12'hfff;
rom[68059] = 12'hfff;
rom[68060] = 12'hfff;
rom[68061] = 12'hfff;
rom[68062] = 12'hfff;
rom[68063] = 12'hfff;
rom[68064] = 12'hfff;
rom[68065] = 12'hfff;
rom[68066] = 12'hfff;
rom[68067] = 12'hfff;
rom[68068] = 12'hfff;
rom[68069] = 12'hfff;
rom[68070] = 12'hfff;
rom[68071] = 12'hfff;
rom[68072] = 12'hfff;
rom[68073] = 12'hfff;
rom[68074] = 12'hfff;
rom[68075] = 12'hfff;
rom[68076] = 12'hfff;
rom[68077] = 12'hfff;
rom[68078] = 12'hfff;
rom[68079] = 12'hfff;
rom[68080] = 12'hfff;
rom[68081] = 12'hfff;
rom[68082] = 12'hfff;
rom[68083] = 12'hfff;
rom[68084] = 12'hfff;
rom[68085] = 12'hfff;
rom[68086] = 12'hfff;
rom[68087] = 12'hfff;
rom[68088] = 12'hfff;
rom[68089] = 12'hfff;
rom[68090] = 12'hfff;
rom[68091] = 12'hfff;
rom[68092] = 12'hfff;
rom[68093] = 12'hfff;
rom[68094] = 12'hfff;
rom[68095] = 12'hfff;
rom[68096] = 12'hfff;
rom[68097] = 12'hfff;
rom[68098] = 12'hfff;
rom[68099] = 12'hfff;
rom[68100] = 12'hfff;
rom[68101] = 12'hfff;
rom[68102] = 12'hfff;
rom[68103] = 12'hfff;
rom[68104] = 12'hfff;
rom[68105] = 12'hfff;
rom[68106] = 12'hfff;
rom[68107] = 12'hfff;
rom[68108] = 12'hfff;
rom[68109] = 12'hfff;
rom[68110] = 12'heee;
rom[68111] = 12'heee;
rom[68112] = 12'hddd;
rom[68113] = 12'hddd;
rom[68114] = 12'hddd;
rom[68115] = 12'hccc;
rom[68116] = 12'hccc;
rom[68117] = 12'hbbb;
rom[68118] = 12'hbbb;
rom[68119] = 12'haaa;
rom[68120] = 12'haaa;
rom[68121] = 12'h999;
rom[68122] = 12'h999;
rom[68123] = 12'h999;
rom[68124] = 12'h999;
rom[68125] = 12'h888;
rom[68126] = 12'h888;
rom[68127] = 12'h888;
rom[68128] = 12'h888;
rom[68129] = 12'h888;
rom[68130] = 12'h777;
rom[68131] = 12'h777;
rom[68132] = 12'h777;
rom[68133] = 12'h777;
rom[68134] = 12'h666;
rom[68135] = 12'h666;
rom[68136] = 12'h666;
rom[68137] = 12'h666;
rom[68138] = 12'h666;
rom[68139] = 12'h555;
rom[68140] = 12'h555;
rom[68141] = 12'h555;
rom[68142] = 12'h555;
rom[68143] = 12'h555;
rom[68144] = 12'h666;
rom[68145] = 12'h666;
rom[68146] = 12'h666;
rom[68147] = 12'h666;
rom[68148] = 12'h666;
rom[68149] = 12'h666;
rom[68150] = 12'h666;
rom[68151] = 12'h666;
rom[68152] = 12'h666;
rom[68153] = 12'h666;
rom[68154] = 12'h666;
rom[68155] = 12'h666;
rom[68156] = 12'h555;
rom[68157] = 12'h555;
rom[68158] = 12'h555;
rom[68159] = 12'h555;
rom[68160] = 12'h444;
rom[68161] = 12'h444;
rom[68162] = 12'h444;
rom[68163] = 12'h333;
rom[68164] = 12'h333;
rom[68165] = 12'h333;
rom[68166] = 12'h333;
rom[68167] = 12'h222;
rom[68168] = 12'h222;
rom[68169] = 12'h222;
rom[68170] = 12'h222;
rom[68171] = 12'h222;
rom[68172] = 12'h222;
rom[68173] = 12'h222;
rom[68174] = 12'h222;
rom[68175] = 12'h222;
rom[68176] = 12'h222;
rom[68177] = 12'h222;
rom[68178] = 12'h111;
rom[68179] = 12'h111;
rom[68180] = 12'h111;
rom[68181] = 12'h111;
rom[68182] = 12'h111;
rom[68183] = 12'h111;
rom[68184] = 12'h111;
rom[68185] = 12'h111;
rom[68186] = 12'h111;
rom[68187] = 12'h111;
rom[68188] = 12'h111;
rom[68189] = 12'h111;
rom[68190] = 12'h111;
rom[68191] = 12'h111;
rom[68192] = 12'h111;
rom[68193] = 12'h111;
rom[68194] = 12'h111;
rom[68195] = 12'h111;
rom[68196] = 12'h111;
rom[68197] = 12'h  0;
rom[68198] = 12'h111;
rom[68199] = 12'h111;
rom[68200] = 12'h  0;
rom[68201] = 12'h111;
rom[68202] = 12'h  0;
rom[68203] = 12'h111;
rom[68204] = 12'h111;
rom[68205] = 12'h111;
rom[68206] = 12'h111;
rom[68207] = 12'h111;
rom[68208] = 12'h111;
rom[68209] = 12'h111;
rom[68210] = 12'h111;
rom[68211] = 12'h111;
rom[68212] = 12'h111;
rom[68213] = 12'h111;
rom[68214] = 12'h111;
rom[68215] = 12'h111;
rom[68216] = 12'h111;
rom[68217] = 12'h111;
rom[68218] = 12'h111;
rom[68219] = 12'h111;
rom[68220] = 12'h  0;
rom[68221] = 12'h  0;
rom[68222] = 12'h  0;
rom[68223] = 12'h  0;
rom[68224] = 12'h  0;
rom[68225] = 12'h  0;
rom[68226] = 12'h  0;
rom[68227] = 12'h  0;
rom[68228] = 12'h  0;
rom[68229] = 12'h  0;
rom[68230] = 12'h  0;
rom[68231] = 12'h  0;
rom[68232] = 12'h  0;
rom[68233] = 12'h  0;
rom[68234] = 12'h  0;
rom[68235] = 12'h  0;
rom[68236] = 12'h  0;
rom[68237] = 12'h  0;
rom[68238] = 12'h  0;
rom[68239] = 12'h  0;
rom[68240] = 12'h  0;
rom[68241] = 12'h  0;
rom[68242] = 12'h  0;
rom[68243] = 12'h  0;
rom[68244] = 12'h  0;
rom[68245] = 12'h  0;
rom[68246] = 12'h  0;
rom[68247] = 12'h  0;
rom[68248] = 12'h  0;
rom[68249] = 12'h  0;
rom[68250] = 12'h  0;
rom[68251] = 12'h  0;
rom[68252] = 12'h  0;
rom[68253] = 12'h  0;
rom[68254] = 12'h  0;
rom[68255] = 12'h  0;
rom[68256] = 12'h  0;
rom[68257] = 12'h  0;
rom[68258] = 12'h  0;
rom[68259] = 12'h  0;
rom[68260] = 12'h  0;
rom[68261] = 12'h  0;
rom[68262] = 12'h  0;
rom[68263] = 12'h  0;
rom[68264] = 12'h  0;
rom[68265] = 12'h  0;
rom[68266] = 12'h  0;
rom[68267] = 12'h  0;
rom[68268] = 12'h  0;
rom[68269] = 12'h  0;
rom[68270] = 12'h111;
rom[68271] = 12'h111;
rom[68272] = 12'h111;
rom[68273] = 12'h222;
rom[68274] = 12'h222;
rom[68275] = 12'h333;
rom[68276] = 12'h333;
rom[68277] = 12'h333;
rom[68278] = 12'h444;
rom[68279] = 12'h555;
rom[68280] = 12'h555;
rom[68281] = 12'h555;
rom[68282] = 12'h333;
rom[68283] = 12'h222;
rom[68284] = 12'h111;
rom[68285] = 12'h111;
rom[68286] = 12'h111;
rom[68287] = 12'h111;
rom[68288] = 12'h111;
rom[68289] = 12'h111;
rom[68290] = 12'h111;
rom[68291] = 12'h111;
rom[68292] = 12'h111;
rom[68293] = 12'h111;
rom[68294] = 12'h111;
rom[68295] = 12'h111;
rom[68296] = 12'h111;
rom[68297] = 12'h111;
rom[68298] = 12'h111;
rom[68299] = 12'h222;
rom[68300] = 12'h333;
rom[68301] = 12'h333;
rom[68302] = 12'h333;
rom[68303] = 12'h333;
rom[68304] = 12'h333;
rom[68305] = 12'h333;
rom[68306] = 12'h333;
rom[68307] = 12'h444;
rom[68308] = 12'h444;
rom[68309] = 12'h555;
rom[68310] = 12'h555;
rom[68311] = 12'h555;
rom[68312] = 12'h555;
rom[68313] = 12'h666;
rom[68314] = 12'h777;
rom[68315] = 12'h777;
rom[68316] = 12'h888;
rom[68317] = 12'h999;
rom[68318] = 12'h999;
rom[68319] = 12'h999;
rom[68320] = 12'h999;
rom[68321] = 12'h999;
rom[68322] = 12'h999;
rom[68323] = 12'haaa;
rom[68324] = 12'haaa;
rom[68325] = 12'haaa;
rom[68326] = 12'haaa;
rom[68327] = 12'haaa;
rom[68328] = 12'haaa;
rom[68329] = 12'hbbb;
rom[68330] = 12'hbbb;
rom[68331] = 12'hbbb;
rom[68332] = 12'hccc;
rom[68333] = 12'hccc;
rom[68334] = 12'hccc;
rom[68335] = 12'hccc;
rom[68336] = 12'hddd;
rom[68337] = 12'hddd;
rom[68338] = 12'heee;
rom[68339] = 12'hfff;
rom[68340] = 12'hfff;
rom[68341] = 12'hfff;
rom[68342] = 12'hfff;
rom[68343] = 12'hfff;
rom[68344] = 12'hfff;
rom[68345] = 12'hfff;
rom[68346] = 12'hfff;
rom[68347] = 12'heee;
rom[68348] = 12'heee;
rom[68349] = 12'hddd;
rom[68350] = 12'hccc;
rom[68351] = 12'hccc;
rom[68352] = 12'hbbb;
rom[68353] = 12'hbbb;
rom[68354] = 12'haaa;
rom[68355] = 12'haaa;
rom[68356] = 12'h999;
rom[68357] = 12'h999;
rom[68358] = 12'h999;
rom[68359] = 12'h888;
rom[68360] = 12'h888;
rom[68361] = 12'h888;
rom[68362] = 12'h888;
rom[68363] = 12'h888;
rom[68364] = 12'h888;
rom[68365] = 12'h888;
rom[68366] = 12'h777;
rom[68367] = 12'h777;
rom[68368] = 12'h777;
rom[68369] = 12'h777;
rom[68370] = 12'h777;
rom[68371] = 12'h777;
rom[68372] = 12'h777;
rom[68373] = 12'h777;
rom[68374] = 12'h777;
rom[68375] = 12'h777;
rom[68376] = 12'h777;
rom[68377] = 12'h777;
rom[68378] = 12'h777;
rom[68379] = 12'h888;
rom[68380] = 12'h888;
rom[68381] = 12'h999;
rom[68382] = 12'haaa;
rom[68383] = 12'haaa;
rom[68384] = 12'hbbb;
rom[68385] = 12'hbbb;
rom[68386] = 12'hbbb;
rom[68387] = 12'haaa;
rom[68388] = 12'h999;
rom[68389] = 12'h888;
rom[68390] = 12'h777;
rom[68391] = 12'h666;
rom[68392] = 12'h666;
rom[68393] = 12'h666;
rom[68394] = 12'h666;
rom[68395] = 12'h666;
rom[68396] = 12'h666;
rom[68397] = 12'h666;
rom[68398] = 12'h666;
rom[68399] = 12'h666;
rom[68400] = 12'hfff;
rom[68401] = 12'hfff;
rom[68402] = 12'hfff;
rom[68403] = 12'hfff;
rom[68404] = 12'hfff;
rom[68405] = 12'hfff;
rom[68406] = 12'hfff;
rom[68407] = 12'hfff;
rom[68408] = 12'hfff;
rom[68409] = 12'hfff;
rom[68410] = 12'hfff;
rom[68411] = 12'hfff;
rom[68412] = 12'hfff;
rom[68413] = 12'hfff;
rom[68414] = 12'hfff;
rom[68415] = 12'hfff;
rom[68416] = 12'hfff;
rom[68417] = 12'hfff;
rom[68418] = 12'hfff;
rom[68419] = 12'hfff;
rom[68420] = 12'hfff;
rom[68421] = 12'hfff;
rom[68422] = 12'hfff;
rom[68423] = 12'hfff;
rom[68424] = 12'hfff;
rom[68425] = 12'hfff;
rom[68426] = 12'hfff;
rom[68427] = 12'hfff;
rom[68428] = 12'hfff;
rom[68429] = 12'hfff;
rom[68430] = 12'hfff;
rom[68431] = 12'hfff;
rom[68432] = 12'hfff;
rom[68433] = 12'hfff;
rom[68434] = 12'hfff;
rom[68435] = 12'hfff;
rom[68436] = 12'hfff;
rom[68437] = 12'hfff;
rom[68438] = 12'hfff;
rom[68439] = 12'hfff;
rom[68440] = 12'hfff;
rom[68441] = 12'hfff;
rom[68442] = 12'hfff;
rom[68443] = 12'hfff;
rom[68444] = 12'hfff;
rom[68445] = 12'hfff;
rom[68446] = 12'hfff;
rom[68447] = 12'hfff;
rom[68448] = 12'hfff;
rom[68449] = 12'hfff;
rom[68450] = 12'hfff;
rom[68451] = 12'hfff;
rom[68452] = 12'hfff;
rom[68453] = 12'hfff;
rom[68454] = 12'hfff;
rom[68455] = 12'hfff;
rom[68456] = 12'hfff;
rom[68457] = 12'hfff;
rom[68458] = 12'hfff;
rom[68459] = 12'hfff;
rom[68460] = 12'hfff;
rom[68461] = 12'hfff;
rom[68462] = 12'hfff;
rom[68463] = 12'hfff;
rom[68464] = 12'hfff;
rom[68465] = 12'hfff;
rom[68466] = 12'hfff;
rom[68467] = 12'hfff;
rom[68468] = 12'hfff;
rom[68469] = 12'hfff;
rom[68470] = 12'hfff;
rom[68471] = 12'hfff;
rom[68472] = 12'hfff;
rom[68473] = 12'hfff;
rom[68474] = 12'hfff;
rom[68475] = 12'hfff;
rom[68476] = 12'hfff;
rom[68477] = 12'hfff;
rom[68478] = 12'hfff;
rom[68479] = 12'hfff;
rom[68480] = 12'hfff;
rom[68481] = 12'hfff;
rom[68482] = 12'hfff;
rom[68483] = 12'hfff;
rom[68484] = 12'hfff;
rom[68485] = 12'hfff;
rom[68486] = 12'hfff;
rom[68487] = 12'hfff;
rom[68488] = 12'hfff;
rom[68489] = 12'hfff;
rom[68490] = 12'hfff;
rom[68491] = 12'hfff;
rom[68492] = 12'hfff;
rom[68493] = 12'hfff;
rom[68494] = 12'hfff;
rom[68495] = 12'hfff;
rom[68496] = 12'hfff;
rom[68497] = 12'hfff;
rom[68498] = 12'hfff;
rom[68499] = 12'hfff;
rom[68500] = 12'hfff;
rom[68501] = 12'hfff;
rom[68502] = 12'hfff;
rom[68503] = 12'hfff;
rom[68504] = 12'hfff;
rom[68505] = 12'hfff;
rom[68506] = 12'hfff;
rom[68507] = 12'hfff;
rom[68508] = 12'hfff;
rom[68509] = 12'hfff;
rom[68510] = 12'heee;
rom[68511] = 12'heee;
rom[68512] = 12'hddd;
rom[68513] = 12'hddd;
rom[68514] = 12'hccc;
rom[68515] = 12'hccc;
rom[68516] = 12'hbbb;
rom[68517] = 12'hbbb;
rom[68518] = 12'haaa;
rom[68519] = 12'haaa;
rom[68520] = 12'haaa;
rom[68521] = 12'h999;
rom[68522] = 12'h999;
rom[68523] = 12'h999;
rom[68524] = 12'h999;
rom[68525] = 12'h888;
rom[68526] = 12'h888;
rom[68527] = 12'h888;
rom[68528] = 12'h888;
rom[68529] = 12'h777;
rom[68530] = 12'h777;
rom[68531] = 12'h777;
rom[68532] = 12'h777;
rom[68533] = 12'h666;
rom[68534] = 12'h666;
rom[68535] = 12'h666;
rom[68536] = 12'h666;
rom[68537] = 12'h555;
rom[68538] = 12'h555;
rom[68539] = 12'h555;
rom[68540] = 12'h555;
rom[68541] = 12'h555;
rom[68542] = 12'h555;
rom[68543] = 12'h555;
rom[68544] = 12'h555;
rom[68545] = 12'h555;
rom[68546] = 12'h555;
rom[68547] = 12'h555;
rom[68548] = 12'h666;
rom[68549] = 12'h666;
rom[68550] = 12'h666;
rom[68551] = 12'h666;
rom[68552] = 12'h666;
rom[68553] = 12'h666;
rom[68554] = 12'h666;
rom[68555] = 12'h666;
rom[68556] = 12'h666;
rom[68557] = 12'h666;
rom[68558] = 12'h666;
rom[68559] = 12'h666;
rom[68560] = 12'h555;
rom[68561] = 12'h444;
rom[68562] = 12'h444;
rom[68563] = 12'h444;
rom[68564] = 12'h444;
rom[68565] = 12'h333;
rom[68566] = 12'h333;
rom[68567] = 12'h333;
rom[68568] = 12'h333;
rom[68569] = 12'h222;
rom[68570] = 12'h222;
rom[68571] = 12'h222;
rom[68572] = 12'h222;
rom[68573] = 12'h222;
rom[68574] = 12'h222;
rom[68575] = 12'h222;
rom[68576] = 12'h222;
rom[68577] = 12'h222;
rom[68578] = 12'h222;
rom[68579] = 12'h222;
rom[68580] = 12'h222;
rom[68581] = 12'h222;
rom[68582] = 12'h111;
rom[68583] = 12'h111;
rom[68584] = 12'h111;
rom[68585] = 12'h111;
rom[68586] = 12'h111;
rom[68587] = 12'h111;
rom[68588] = 12'h111;
rom[68589] = 12'h111;
rom[68590] = 12'h111;
rom[68591] = 12'h111;
rom[68592] = 12'h111;
rom[68593] = 12'h111;
rom[68594] = 12'h111;
rom[68595] = 12'h111;
rom[68596] = 12'h111;
rom[68597] = 12'h111;
rom[68598] = 12'h111;
rom[68599] = 12'h111;
rom[68600] = 12'h111;
rom[68601] = 12'h111;
rom[68602] = 12'h111;
rom[68603] = 12'h111;
rom[68604] = 12'h111;
rom[68605] = 12'h111;
rom[68606] = 12'h111;
rom[68607] = 12'h111;
rom[68608] = 12'h222;
rom[68609] = 12'h111;
rom[68610] = 12'h111;
rom[68611] = 12'h111;
rom[68612] = 12'h111;
rom[68613] = 12'h111;
rom[68614] = 12'h111;
rom[68615] = 12'h111;
rom[68616] = 12'h111;
rom[68617] = 12'h111;
rom[68618] = 12'h111;
rom[68619] = 12'h  0;
rom[68620] = 12'h  0;
rom[68621] = 12'h  0;
rom[68622] = 12'h  0;
rom[68623] = 12'h  0;
rom[68624] = 12'h  0;
rom[68625] = 12'h  0;
rom[68626] = 12'h  0;
rom[68627] = 12'h  0;
rom[68628] = 12'h  0;
rom[68629] = 12'h  0;
rom[68630] = 12'h  0;
rom[68631] = 12'h  0;
rom[68632] = 12'h  0;
rom[68633] = 12'h  0;
rom[68634] = 12'h  0;
rom[68635] = 12'h  0;
rom[68636] = 12'h  0;
rom[68637] = 12'h  0;
rom[68638] = 12'h  0;
rom[68639] = 12'h  0;
rom[68640] = 12'h  0;
rom[68641] = 12'h  0;
rom[68642] = 12'h  0;
rom[68643] = 12'h  0;
rom[68644] = 12'h  0;
rom[68645] = 12'h  0;
rom[68646] = 12'h  0;
rom[68647] = 12'h  0;
rom[68648] = 12'h  0;
rom[68649] = 12'h  0;
rom[68650] = 12'h  0;
rom[68651] = 12'h  0;
rom[68652] = 12'h  0;
rom[68653] = 12'h  0;
rom[68654] = 12'h  0;
rom[68655] = 12'h  0;
rom[68656] = 12'h  0;
rom[68657] = 12'h  0;
rom[68658] = 12'h  0;
rom[68659] = 12'h  0;
rom[68660] = 12'h  0;
rom[68661] = 12'h  0;
rom[68662] = 12'h  0;
rom[68663] = 12'h  0;
rom[68664] = 12'h  0;
rom[68665] = 12'h  0;
rom[68666] = 12'h  0;
rom[68667] = 12'h  0;
rom[68668] = 12'h  0;
rom[68669] = 12'h  0;
rom[68670] = 12'h111;
rom[68671] = 12'h111;
rom[68672] = 12'h111;
rom[68673] = 12'h222;
rom[68674] = 12'h222;
rom[68675] = 12'h333;
rom[68676] = 12'h333;
rom[68677] = 12'h333;
rom[68678] = 12'h444;
rom[68679] = 12'h555;
rom[68680] = 12'h666;
rom[68681] = 12'h555;
rom[68682] = 12'h333;
rom[68683] = 12'h111;
rom[68684] = 12'h111;
rom[68685] = 12'h111;
rom[68686] = 12'h111;
rom[68687] = 12'h111;
rom[68688] = 12'h111;
rom[68689] = 12'h111;
rom[68690] = 12'h111;
rom[68691] = 12'h111;
rom[68692] = 12'h111;
rom[68693] = 12'h111;
rom[68694] = 12'h111;
rom[68695] = 12'h111;
rom[68696] = 12'h111;
rom[68697] = 12'h111;
rom[68698] = 12'h111;
rom[68699] = 12'h222;
rom[68700] = 12'h333;
rom[68701] = 12'h333;
rom[68702] = 12'h333;
rom[68703] = 12'h333;
rom[68704] = 12'h333;
rom[68705] = 12'h333;
rom[68706] = 12'h333;
rom[68707] = 12'h444;
rom[68708] = 12'h444;
rom[68709] = 12'h555;
rom[68710] = 12'h555;
rom[68711] = 12'h555;
rom[68712] = 12'h555;
rom[68713] = 12'h666;
rom[68714] = 12'h777;
rom[68715] = 12'h777;
rom[68716] = 12'h888;
rom[68717] = 12'h999;
rom[68718] = 12'h999;
rom[68719] = 12'haaa;
rom[68720] = 12'haaa;
rom[68721] = 12'haaa;
rom[68722] = 12'haaa;
rom[68723] = 12'haaa;
rom[68724] = 12'haaa;
rom[68725] = 12'haaa;
rom[68726] = 12'haaa;
rom[68727] = 12'hbbb;
rom[68728] = 12'hbbb;
rom[68729] = 12'hbbb;
rom[68730] = 12'hbbb;
rom[68731] = 12'hbbb;
rom[68732] = 12'hccc;
rom[68733] = 12'hccc;
rom[68734] = 12'hddd;
rom[68735] = 12'hddd;
rom[68736] = 12'hddd;
rom[68737] = 12'heee;
rom[68738] = 12'hfff;
rom[68739] = 12'hfff;
rom[68740] = 12'hfff;
rom[68741] = 12'hfff;
rom[68742] = 12'hfff;
rom[68743] = 12'hfff;
rom[68744] = 12'hfff;
rom[68745] = 12'hfff;
rom[68746] = 12'heee;
rom[68747] = 12'heee;
rom[68748] = 12'hddd;
rom[68749] = 12'hccc;
rom[68750] = 12'hccc;
rom[68751] = 12'hbbb;
rom[68752] = 12'haaa;
rom[68753] = 12'haaa;
rom[68754] = 12'haaa;
rom[68755] = 12'h999;
rom[68756] = 12'h999;
rom[68757] = 12'h999;
rom[68758] = 12'h888;
rom[68759] = 12'h888;
rom[68760] = 12'h888;
rom[68761] = 12'h888;
rom[68762] = 12'h888;
rom[68763] = 12'h888;
rom[68764] = 12'h888;
rom[68765] = 12'h888;
rom[68766] = 12'h777;
rom[68767] = 12'h777;
rom[68768] = 12'h777;
rom[68769] = 12'h777;
rom[68770] = 12'h777;
rom[68771] = 12'h777;
rom[68772] = 12'h777;
rom[68773] = 12'h777;
rom[68774] = 12'h777;
rom[68775] = 12'h777;
rom[68776] = 12'h777;
rom[68777] = 12'h777;
rom[68778] = 12'h777;
rom[68779] = 12'h777;
rom[68780] = 12'h888;
rom[68781] = 12'h888;
rom[68782] = 12'h999;
rom[68783] = 12'h999;
rom[68784] = 12'haaa;
rom[68785] = 12'hbbb;
rom[68786] = 12'hbbb;
rom[68787] = 12'hbbb;
rom[68788] = 12'haaa;
rom[68789] = 12'h999;
rom[68790] = 12'h888;
rom[68791] = 12'h777;
rom[68792] = 12'h666;
rom[68793] = 12'h666;
rom[68794] = 12'h666;
rom[68795] = 12'h666;
rom[68796] = 12'h666;
rom[68797] = 12'h666;
rom[68798] = 12'h666;
rom[68799] = 12'h555;
rom[68800] = 12'hfff;
rom[68801] = 12'hfff;
rom[68802] = 12'hfff;
rom[68803] = 12'hfff;
rom[68804] = 12'hfff;
rom[68805] = 12'hfff;
rom[68806] = 12'hfff;
rom[68807] = 12'hfff;
rom[68808] = 12'hfff;
rom[68809] = 12'hfff;
rom[68810] = 12'hfff;
rom[68811] = 12'hfff;
rom[68812] = 12'hfff;
rom[68813] = 12'hfff;
rom[68814] = 12'hfff;
rom[68815] = 12'hfff;
rom[68816] = 12'hfff;
rom[68817] = 12'hfff;
rom[68818] = 12'hfff;
rom[68819] = 12'hfff;
rom[68820] = 12'hfff;
rom[68821] = 12'hfff;
rom[68822] = 12'hfff;
rom[68823] = 12'hfff;
rom[68824] = 12'hfff;
rom[68825] = 12'hfff;
rom[68826] = 12'hfff;
rom[68827] = 12'hfff;
rom[68828] = 12'hfff;
rom[68829] = 12'hfff;
rom[68830] = 12'hfff;
rom[68831] = 12'hfff;
rom[68832] = 12'hfff;
rom[68833] = 12'hfff;
rom[68834] = 12'hfff;
rom[68835] = 12'hfff;
rom[68836] = 12'hfff;
rom[68837] = 12'hfff;
rom[68838] = 12'hfff;
rom[68839] = 12'hfff;
rom[68840] = 12'hfff;
rom[68841] = 12'hfff;
rom[68842] = 12'hfff;
rom[68843] = 12'hfff;
rom[68844] = 12'hfff;
rom[68845] = 12'hfff;
rom[68846] = 12'hfff;
rom[68847] = 12'hfff;
rom[68848] = 12'hfff;
rom[68849] = 12'hfff;
rom[68850] = 12'hfff;
rom[68851] = 12'hfff;
rom[68852] = 12'hfff;
rom[68853] = 12'hfff;
rom[68854] = 12'hfff;
rom[68855] = 12'hfff;
rom[68856] = 12'hfff;
rom[68857] = 12'hfff;
rom[68858] = 12'hfff;
rom[68859] = 12'hfff;
rom[68860] = 12'hfff;
rom[68861] = 12'hfff;
rom[68862] = 12'hfff;
rom[68863] = 12'hfff;
rom[68864] = 12'hfff;
rom[68865] = 12'hfff;
rom[68866] = 12'hfff;
rom[68867] = 12'hfff;
rom[68868] = 12'hfff;
rom[68869] = 12'hfff;
rom[68870] = 12'hfff;
rom[68871] = 12'hfff;
rom[68872] = 12'hfff;
rom[68873] = 12'hfff;
rom[68874] = 12'hfff;
rom[68875] = 12'hfff;
rom[68876] = 12'hfff;
rom[68877] = 12'hfff;
rom[68878] = 12'hfff;
rom[68879] = 12'hfff;
rom[68880] = 12'hfff;
rom[68881] = 12'hfff;
rom[68882] = 12'hfff;
rom[68883] = 12'hfff;
rom[68884] = 12'hfff;
rom[68885] = 12'hfff;
rom[68886] = 12'hfff;
rom[68887] = 12'hfff;
rom[68888] = 12'hfff;
rom[68889] = 12'hfff;
rom[68890] = 12'hfff;
rom[68891] = 12'hfff;
rom[68892] = 12'hfff;
rom[68893] = 12'hfff;
rom[68894] = 12'hfff;
rom[68895] = 12'hfff;
rom[68896] = 12'hfff;
rom[68897] = 12'hfff;
rom[68898] = 12'hfff;
rom[68899] = 12'hfff;
rom[68900] = 12'hfff;
rom[68901] = 12'hfff;
rom[68902] = 12'hfff;
rom[68903] = 12'hfff;
rom[68904] = 12'hfff;
rom[68905] = 12'hfff;
rom[68906] = 12'hfff;
rom[68907] = 12'hfff;
rom[68908] = 12'hfff;
rom[68909] = 12'hfff;
rom[68910] = 12'heee;
rom[68911] = 12'heee;
rom[68912] = 12'hddd;
rom[68913] = 12'hddd;
rom[68914] = 12'hccc;
rom[68915] = 12'hbbb;
rom[68916] = 12'hbbb;
rom[68917] = 12'haaa;
rom[68918] = 12'haaa;
rom[68919] = 12'haaa;
rom[68920] = 12'h999;
rom[68921] = 12'h999;
rom[68922] = 12'h999;
rom[68923] = 12'h888;
rom[68924] = 12'h888;
rom[68925] = 12'h888;
rom[68926] = 12'h888;
rom[68927] = 12'h888;
rom[68928] = 12'h888;
rom[68929] = 12'h777;
rom[68930] = 12'h777;
rom[68931] = 12'h777;
rom[68932] = 12'h777;
rom[68933] = 12'h666;
rom[68934] = 12'h666;
rom[68935] = 12'h666;
rom[68936] = 12'h666;
rom[68937] = 12'h666;
rom[68938] = 12'h555;
rom[68939] = 12'h555;
rom[68940] = 12'h555;
rom[68941] = 12'h555;
rom[68942] = 12'h555;
rom[68943] = 12'h555;
rom[68944] = 12'h555;
rom[68945] = 12'h555;
rom[68946] = 12'h555;
rom[68947] = 12'h555;
rom[68948] = 12'h555;
rom[68949] = 12'h555;
rom[68950] = 12'h555;
rom[68951] = 12'h666;
rom[68952] = 12'h555;
rom[68953] = 12'h555;
rom[68954] = 12'h666;
rom[68955] = 12'h666;
rom[68956] = 12'h666;
rom[68957] = 12'h666;
rom[68958] = 12'h666;
rom[68959] = 12'h666;
rom[68960] = 12'h555;
rom[68961] = 12'h555;
rom[68962] = 12'h555;
rom[68963] = 12'h444;
rom[68964] = 12'h444;
rom[68965] = 12'h444;
rom[68966] = 12'h444;
rom[68967] = 12'h444;
rom[68968] = 12'h333;
rom[68969] = 12'h333;
rom[68970] = 12'h333;
rom[68971] = 12'h333;
rom[68972] = 12'h333;
rom[68973] = 12'h333;
rom[68974] = 12'h333;
rom[68975] = 12'h222;
rom[68976] = 12'h222;
rom[68977] = 12'h222;
rom[68978] = 12'h222;
rom[68979] = 12'h222;
rom[68980] = 12'h222;
rom[68981] = 12'h222;
rom[68982] = 12'h222;
rom[68983] = 12'h222;
rom[68984] = 12'h222;
rom[68985] = 12'h222;
rom[68986] = 12'h111;
rom[68987] = 12'h111;
rom[68988] = 12'h222;
rom[68989] = 12'h222;
rom[68990] = 12'h222;
rom[68991] = 12'h222;
rom[68992] = 12'h111;
rom[68993] = 12'h111;
rom[68994] = 12'h111;
rom[68995] = 12'h111;
rom[68996] = 12'h111;
rom[68997] = 12'h111;
rom[68998] = 12'h111;
rom[68999] = 12'h111;
rom[69000] = 12'h111;
rom[69001] = 12'h111;
rom[69002] = 12'h111;
rom[69003] = 12'h111;
rom[69004] = 12'h111;
rom[69005] = 12'h111;
rom[69006] = 12'h111;
rom[69007] = 12'h111;
rom[69008] = 12'h222;
rom[69009] = 12'h111;
rom[69010] = 12'h111;
rom[69011] = 12'h111;
rom[69012] = 12'h111;
rom[69013] = 12'h111;
rom[69014] = 12'h111;
rom[69015] = 12'h111;
rom[69016] = 12'h111;
rom[69017] = 12'h111;
rom[69018] = 12'h111;
rom[69019] = 12'h  0;
rom[69020] = 12'h  0;
rom[69021] = 12'h  0;
rom[69022] = 12'h  0;
rom[69023] = 12'h  0;
rom[69024] = 12'h  0;
rom[69025] = 12'h  0;
rom[69026] = 12'h  0;
rom[69027] = 12'h  0;
rom[69028] = 12'h  0;
rom[69029] = 12'h  0;
rom[69030] = 12'h  0;
rom[69031] = 12'h  0;
rom[69032] = 12'h  0;
rom[69033] = 12'h  0;
rom[69034] = 12'h  0;
rom[69035] = 12'h  0;
rom[69036] = 12'h  0;
rom[69037] = 12'h  0;
rom[69038] = 12'h  0;
rom[69039] = 12'h  0;
rom[69040] = 12'h  0;
rom[69041] = 12'h  0;
rom[69042] = 12'h  0;
rom[69043] = 12'h  0;
rom[69044] = 12'h  0;
rom[69045] = 12'h  0;
rom[69046] = 12'h  0;
rom[69047] = 12'h  0;
rom[69048] = 12'h  0;
rom[69049] = 12'h  0;
rom[69050] = 12'h  0;
rom[69051] = 12'h  0;
rom[69052] = 12'h  0;
rom[69053] = 12'h  0;
rom[69054] = 12'h  0;
rom[69055] = 12'h  0;
rom[69056] = 12'h  0;
rom[69057] = 12'h  0;
rom[69058] = 12'h  0;
rom[69059] = 12'h  0;
rom[69060] = 12'h  0;
rom[69061] = 12'h  0;
rom[69062] = 12'h  0;
rom[69063] = 12'h  0;
rom[69064] = 12'h  0;
rom[69065] = 12'h  0;
rom[69066] = 12'h  0;
rom[69067] = 12'h  0;
rom[69068] = 12'h  0;
rom[69069] = 12'h  0;
rom[69070] = 12'h111;
rom[69071] = 12'h111;
rom[69072] = 12'h222;
rom[69073] = 12'h222;
rom[69074] = 12'h222;
rom[69075] = 12'h222;
rom[69076] = 12'h333;
rom[69077] = 12'h333;
rom[69078] = 12'h444;
rom[69079] = 12'h555;
rom[69080] = 12'h666;
rom[69081] = 12'h555;
rom[69082] = 12'h333;
rom[69083] = 12'h111;
rom[69084] = 12'h111;
rom[69085] = 12'h111;
rom[69086] = 12'h111;
rom[69087] = 12'h111;
rom[69088] = 12'h111;
rom[69089] = 12'h111;
rom[69090] = 12'h111;
rom[69091] = 12'h111;
rom[69092] = 12'h111;
rom[69093] = 12'h111;
rom[69094] = 12'h111;
rom[69095] = 12'h111;
rom[69096] = 12'h111;
rom[69097] = 12'h111;
rom[69098] = 12'h111;
rom[69099] = 12'h222;
rom[69100] = 12'h222;
rom[69101] = 12'h333;
rom[69102] = 12'h333;
rom[69103] = 12'h333;
rom[69104] = 12'h333;
rom[69105] = 12'h333;
rom[69106] = 12'h333;
rom[69107] = 12'h444;
rom[69108] = 12'h444;
rom[69109] = 12'h555;
rom[69110] = 12'h555;
rom[69111] = 12'h666;
rom[69112] = 12'h666;
rom[69113] = 12'h666;
rom[69114] = 12'h777;
rom[69115] = 12'h888;
rom[69116] = 12'h888;
rom[69117] = 12'h999;
rom[69118] = 12'haaa;
rom[69119] = 12'haaa;
rom[69120] = 12'haaa;
rom[69121] = 12'haaa;
rom[69122] = 12'haaa;
rom[69123] = 12'haaa;
rom[69124] = 12'haaa;
rom[69125] = 12'haaa;
rom[69126] = 12'hbbb;
rom[69127] = 12'hbbb;
rom[69128] = 12'hbbb;
rom[69129] = 12'hbbb;
rom[69130] = 12'hbbb;
rom[69131] = 12'hccc;
rom[69132] = 12'hccc;
rom[69133] = 12'hddd;
rom[69134] = 12'hddd;
rom[69135] = 12'hddd;
rom[69136] = 12'heee;
rom[69137] = 12'hfff;
rom[69138] = 12'hfff;
rom[69139] = 12'hfff;
rom[69140] = 12'hfff;
rom[69141] = 12'hfff;
rom[69142] = 12'hfff;
rom[69143] = 12'hfff;
rom[69144] = 12'hfff;
rom[69145] = 12'hfff;
rom[69146] = 12'heee;
rom[69147] = 12'hddd;
rom[69148] = 12'hddd;
rom[69149] = 12'hccc;
rom[69150] = 12'hbbb;
rom[69151] = 12'hbbb;
rom[69152] = 12'haaa;
rom[69153] = 12'haaa;
rom[69154] = 12'h999;
rom[69155] = 12'h999;
rom[69156] = 12'h999;
rom[69157] = 12'h999;
rom[69158] = 12'h888;
rom[69159] = 12'h888;
rom[69160] = 12'h888;
rom[69161] = 12'h888;
rom[69162] = 12'h888;
rom[69163] = 12'h888;
rom[69164] = 12'h888;
rom[69165] = 12'h777;
rom[69166] = 12'h777;
rom[69167] = 12'h777;
rom[69168] = 12'h777;
rom[69169] = 12'h777;
rom[69170] = 12'h777;
rom[69171] = 12'h777;
rom[69172] = 12'h777;
rom[69173] = 12'h777;
rom[69174] = 12'h777;
rom[69175] = 12'h777;
rom[69176] = 12'h666;
rom[69177] = 12'h777;
rom[69178] = 12'h777;
rom[69179] = 12'h777;
rom[69180] = 12'h777;
rom[69181] = 12'h888;
rom[69182] = 12'h888;
rom[69183] = 12'h888;
rom[69184] = 12'h999;
rom[69185] = 12'haaa;
rom[69186] = 12'haaa;
rom[69187] = 12'hbbb;
rom[69188] = 12'hbbb;
rom[69189] = 12'haaa;
rom[69190] = 12'h999;
rom[69191] = 12'h888;
rom[69192] = 12'h777;
rom[69193] = 12'h777;
rom[69194] = 12'h666;
rom[69195] = 12'h666;
rom[69196] = 12'h666;
rom[69197] = 12'h666;
rom[69198] = 12'h555;
rom[69199] = 12'h555;
rom[69200] = 12'hfff;
rom[69201] = 12'hfff;
rom[69202] = 12'hfff;
rom[69203] = 12'hfff;
rom[69204] = 12'hfff;
rom[69205] = 12'hfff;
rom[69206] = 12'hfff;
rom[69207] = 12'hfff;
rom[69208] = 12'hfff;
rom[69209] = 12'hfff;
rom[69210] = 12'hfff;
rom[69211] = 12'hfff;
rom[69212] = 12'hfff;
rom[69213] = 12'hfff;
rom[69214] = 12'hfff;
rom[69215] = 12'hfff;
rom[69216] = 12'hfff;
rom[69217] = 12'hfff;
rom[69218] = 12'hfff;
rom[69219] = 12'hfff;
rom[69220] = 12'hfff;
rom[69221] = 12'hfff;
rom[69222] = 12'hfff;
rom[69223] = 12'hfff;
rom[69224] = 12'hfff;
rom[69225] = 12'hfff;
rom[69226] = 12'hfff;
rom[69227] = 12'hfff;
rom[69228] = 12'hfff;
rom[69229] = 12'hfff;
rom[69230] = 12'hfff;
rom[69231] = 12'hfff;
rom[69232] = 12'hfff;
rom[69233] = 12'hfff;
rom[69234] = 12'hfff;
rom[69235] = 12'hfff;
rom[69236] = 12'hfff;
rom[69237] = 12'hfff;
rom[69238] = 12'hfff;
rom[69239] = 12'hfff;
rom[69240] = 12'hfff;
rom[69241] = 12'hfff;
rom[69242] = 12'hfff;
rom[69243] = 12'hfff;
rom[69244] = 12'hfff;
rom[69245] = 12'hfff;
rom[69246] = 12'hfff;
rom[69247] = 12'hfff;
rom[69248] = 12'hfff;
rom[69249] = 12'hfff;
rom[69250] = 12'hfff;
rom[69251] = 12'hfff;
rom[69252] = 12'hfff;
rom[69253] = 12'hfff;
rom[69254] = 12'hfff;
rom[69255] = 12'hfff;
rom[69256] = 12'hfff;
rom[69257] = 12'hfff;
rom[69258] = 12'hfff;
rom[69259] = 12'hfff;
rom[69260] = 12'hfff;
rom[69261] = 12'hfff;
rom[69262] = 12'hfff;
rom[69263] = 12'hfff;
rom[69264] = 12'hfff;
rom[69265] = 12'hfff;
rom[69266] = 12'hfff;
rom[69267] = 12'hfff;
rom[69268] = 12'hfff;
rom[69269] = 12'hfff;
rom[69270] = 12'hfff;
rom[69271] = 12'hfff;
rom[69272] = 12'hfff;
rom[69273] = 12'hfff;
rom[69274] = 12'hfff;
rom[69275] = 12'hfff;
rom[69276] = 12'hfff;
rom[69277] = 12'hfff;
rom[69278] = 12'hfff;
rom[69279] = 12'hfff;
rom[69280] = 12'hfff;
rom[69281] = 12'hfff;
rom[69282] = 12'hfff;
rom[69283] = 12'hfff;
rom[69284] = 12'hfff;
rom[69285] = 12'hfff;
rom[69286] = 12'hfff;
rom[69287] = 12'hfff;
rom[69288] = 12'hfff;
rom[69289] = 12'hfff;
rom[69290] = 12'hfff;
rom[69291] = 12'hfff;
rom[69292] = 12'hfff;
rom[69293] = 12'hfff;
rom[69294] = 12'hfff;
rom[69295] = 12'hfff;
rom[69296] = 12'hfff;
rom[69297] = 12'hfff;
rom[69298] = 12'hfff;
rom[69299] = 12'hfff;
rom[69300] = 12'hfff;
rom[69301] = 12'hfff;
rom[69302] = 12'hfff;
rom[69303] = 12'hfff;
rom[69304] = 12'hfff;
rom[69305] = 12'hfff;
rom[69306] = 12'hfff;
rom[69307] = 12'hfff;
rom[69308] = 12'hfff;
rom[69309] = 12'hfff;
rom[69310] = 12'heee;
rom[69311] = 12'heee;
rom[69312] = 12'hddd;
rom[69313] = 12'hccc;
rom[69314] = 12'hccc;
rom[69315] = 12'hbbb;
rom[69316] = 12'hbbb;
rom[69317] = 12'haaa;
rom[69318] = 12'haaa;
rom[69319] = 12'haaa;
rom[69320] = 12'h999;
rom[69321] = 12'h999;
rom[69322] = 12'h999;
rom[69323] = 12'h888;
rom[69324] = 12'h888;
rom[69325] = 12'h888;
rom[69326] = 12'h888;
rom[69327] = 12'h777;
rom[69328] = 12'h888;
rom[69329] = 12'h777;
rom[69330] = 12'h777;
rom[69331] = 12'h777;
rom[69332] = 12'h777;
rom[69333] = 12'h666;
rom[69334] = 12'h666;
rom[69335] = 12'h666;
rom[69336] = 12'h666;
rom[69337] = 12'h555;
rom[69338] = 12'h555;
rom[69339] = 12'h555;
rom[69340] = 12'h555;
rom[69341] = 12'h555;
rom[69342] = 12'h555;
rom[69343] = 12'h555;
rom[69344] = 12'h555;
rom[69345] = 12'h555;
rom[69346] = 12'h555;
rom[69347] = 12'h555;
rom[69348] = 12'h555;
rom[69349] = 12'h555;
rom[69350] = 12'h555;
rom[69351] = 12'h555;
rom[69352] = 12'h555;
rom[69353] = 12'h555;
rom[69354] = 12'h555;
rom[69355] = 12'h555;
rom[69356] = 12'h555;
rom[69357] = 12'h555;
rom[69358] = 12'h555;
rom[69359] = 12'h555;
rom[69360] = 12'h666;
rom[69361] = 12'h555;
rom[69362] = 12'h555;
rom[69363] = 12'h555;
rom[69364] = 12'h555;
rom[69365] = 12'h555;
rom[69366] = 12'h555;
rom[69367] = 12'h444;
rom[69368] = 12'h444;
rom[69369] = 12'h444;
rom[69370] = 12'h444;
rom[69371] = 12'h333;
rom[69372] = 12'h333;
rom[69373] = 12'h333;
rom[69374] = 12'h333;
rom[69375] = 12'h333;
rom[69376] = 12'h333;
rom[69377] = 12'h333;
rom[69378] = 12'h333;
rom[69379] = 12'h333;
rom[69380] = 12'h333;
rom[69381] = 12'h222;
rom[69382] = 12'h222;
rom[69383] = 12'h222;
rom[69384] = 12'h222;
rom[69385] = 12'h222;
rom[69386] = 12'h222;
rom[69387] = 12'h222;
rom[69388] = 12'h222;
rom[69389] = 12'h222;
rom[69390] = 12'h222;
rom[69391] = 12'h222;
rom[69392] = 12'h222;
rom[69393] = 12'h222;
rom[69394] = 12'h111;
rom[69395] = 12'h111;
rom[69396] = 12'h111;
rom[69397] = 12'h111;
rom[69398] = 12'h111;
rom[69399] = 12'h111;
rom[69400] = 12'h111;
rom[69401] = 12'h111;
rom[69402] = 12'h111;
rom[69403] = 12'h111;
rom[69404] = 12'h222;
rom[69405] = 12'h111;
rom[69406] = 12'h111;
rom[69407] = 12'h111;
rom[69408] = 12'h222;
rom[69409] = 12'h111;
rom[69410] = 12'h111;
rom[69411] = 12'h111;
rom[69412] = 12'h111;
rom[69413] = 12'h111;
rom[69414] = 12'h111;
rom[69415] = 12'h111;
rom[69416] = 12'h111;
rom[69417] = 12'h111;
rom[69418] = 12'h  0;
rom[69419] = 12'h  0;
rom[69420] = 12'h  0;
rom[69421] = 12'h  0;
rom[69422] = 12'h  0;
rom[69423] = 12'h  0;
rom[69424] = 12'h  0;
rom[69425] = 12'h  0;
rom[69426] = 12'h  0;
rom[69427] = 12'h  0;
rom[69428] = 12'h  0;
rom[69429] = 12'h  0;
rom[69430] = 12'h  0;
rom[69431] = 12'h  0;
rom[69432] = 12'h  0;
rom[69433] = 12'h  0;
rom[69434] = 12'h  0;
rom[69435] = 12'h  0;
rom[69436] = 12'h  0;
rom[69437] = 12'h  0;
rom[69438] = 12'h  0;
rom[69439] = 12'h  0;
rom[69440] = 12'h  0;
rom[69441] = 12'h  0;
rom[69442] = 12'h  0;
rom[69443] = 12'h  0;
rom[69444] = 12'h  0;
rom[69445] = 12'h  0;
rom[69446] = 12'h  0;
rom[69447] = 12'h  0;
rom[69448] = 12'h  0;
rom[69449] = 12'h  0;
rom[69450] = 12'h  0;
rom[69451] = 12'h  0;
rom[69452] = 12'h  0;
rom[69453] = 12'h  0;
rom[69454] = 12'h  0;
rom[69455] = 12'h  0;
rom[69456] = 12'h  0;
rom[69457] = 12'h  0;
rom[69458] = 12'h  0;
rom[69459] = 12'h  0;
rom[69460] = 12'h  0;
rom[69461] = 12'h  0;
rom[69462] = 12'h  0;
rom[69463] = 12'h  0;
rom[69464] = 12'h  0;
rom[69465] = 12'h  0;
rom[69466] = 12'h  0;
rom[69467] = 12'h  0;
rom[69468] = 12'h  0;
rom[69469] = 12'h  0;
rom[69470] = 12'h111;
rom[69471] = 12'h111;
rom[69472] = 12'h222;
rom[69473] = 12'h222;
rom[69474] = 12'h222;
rom[69475] = 12'h222;
rom[69476] = 12'h333;
rom[69477] = 12'h333;
rom[69478] = 12'h444;
rom[69479] = 12'h555;
rom[69480] = 12'h666;
rom[69481] = 12'h555;
rom[69482] = 12'h333;
rom[69483] = 12'h111;
rom[69484] = 12'h111;
rom[69485] = 12'h111;
rom[69486] = 12'h111;
rom[69487] = 12'h111;
rom[69488] = 12'h111;
rom[69489] = 12'h  0;
rom[69490] = 12'h  0;
rom[69491] = 12'h  0;
rom[69492] = 12'h  0;
rom[69493] = 12'h111;
rom[69494] = 12'h111;
rom[69495] = 12'h111;
rom[69496] = 12'h111;
rom[69497] = 12'h111;
rom[69498] = 12'h111;
rom[69499] = 12'h222;
rom[69500] = 12'h222;
rom[69501] = 12'h333;
rom[69502] = 12'h333;
rom[69503] = 12'h333;
rom[69504] = 12'h333;
rom[69505] = 12'h333;
rom[69506] = 12'h444;
rom[69507] = 12'h444;
rom[69508] = 12'h444;
rom[69509] = 12'h555;
rom[69510] = 12'h555;
rom[69511] = 12'h666;
rom[69512] = 12'h666;
rom[69513] = 12'h666;
rom[69514] = 12'h777;
rom[69515] = 12'h888;
rom[69516] = 12'h999;
rom[69517] = 12'h999;
rom[69518] = 12'haaa;
rom[69519] = 12'haaa;
rom[69520] = 12'haaa;
rom[69521] = 12'haaa;
rom[69522] = 12'haaa;
rom[69523] = 12'haaa;
rom[69524] = 12'haaa;
rom[69525] = 12'hbbb;
rom[69526] = 12'hbbb;
rom[69527] = 12'hbbb;
rom[69528] = 12'hbbb;
rom[69529] = 12'hccc;
rom[69530] = 12'hccc;
rom[69531] = 12'hccc;
rom[69532] = 12'hddd;
rom[69533] = 12'hddd;
rom[69534] = 12'heee;
rom[69535] = 12'heee;
rom[69536] = 12'heee;
rom[69537] = 12'hfff;
rom[69538] = 12'hfff;
rom[69539] = 12'hfff;
rom[69540] = 12'hfff;
rom[69541] = 12'hfff;
rom[69542] = 12'hfff;
rom[69543] = 12'hfff;
rom[69544] = 12'hfff;
rom[69545] = 12'heee;
rom[69546] = 12'hddd;
rom[69547] = 12'hddd;
rom[69548] = 12'hccc;
rom[69549] = 12'hbbb;
rom[69550] = 12'hbbb;
rom[69551] = 12'haaa;
rom[69552] = 12'haaa;
rom[69553] = 12'haaa;
rom[69554] = 12'h999;
rom[69555] = 12'h999;
rom[69556] = 12'h999;
rom[69557] = 12'h888;
rom[69558] = 12'h888;
rom[69559] = 12'h888;
rom[69560] = 12'h888;
rom[69561] = 12'h888;
rom[69562] = 12'h888;
rom[69563] = 12'h777;
rom[69564] = 12'h777;
rom[69565] = 12'h777;
rom[69566] = 12'h777;
rom[69567] = 12'h777;
rom[69568] = 12'h777;
rom[69569] = 12'h777;
rom[69570] = 12'h777;
rom[69571] = 12'h777;
rom[69572] = 12'h777;
rom[69573] = 12'h777;
rom[69574] = 12'h777;
rom[69575] = 12'h777;
rom[69576] = 12'h666;
rom[69577] = 12'h777;
rom[69578] = 12'h777;
rom[69579] = 12'h777;
rom[69580] = 12'h777;
rom[69581] = 12'h777;
rom[69582] = 12'h777;
rom[69583] = 12'h777;
rom[69584] = 12'h888;
rom[69585] = 12'h999;
rom[69586] = 12'haaa;
rom[69587] = 12'haaa;
rom[69588] = 12'hbbb;
rom[69589] = 12'haaa;
rom[69590] = 12'haaa;
rom[69591] = 12'h999;
rom[69592] = 12'h888;
rom[69593] = 12'h777;
rom[69594] = 12'h777;
rom[69595] = 12'h666;
rom[69596] = 12'h666;
rom[69597] = 12'h555;
rom[69598] = 12'h555;
rom[69599] = 12'h555;
rom[69600] = 12'hfff;
rom[69601] = 12'hfff;
rom[69602] = 12'hfff;
rom[69603] = 12'hfff;
rom[69604] = 12'hfff;
rom[69605] = 12'hfff;
rom[69606] = 12'hfff;
rom[69607] = 12'hfff;
rom[69608] = 12'hfff;
rom[69609] = 12'hfff;
rom[69610] = 12'hfff;
rom[69611] = 12'hfff;
rom[69612] = 12'hfff;
rom[69613] = 12'hfff;
rom[69614] = 12'hfff;
rom[69615] = 12'hfff;
rom[69616] = 12'hfff;
rom[69617] = 12'hfff;
rom[69618] = 12'hfff;
rom[69619] = 12'hfff;
rom[69620] = 12'hfff;
rom[69621] = 12'hfff;
rom[69622] = 12'hfff;
rom[69623] = 12'hfff;
rom[69624] = 12'hfff;
rom[69625] = 12'hfff;
rom[69626] = 12'hfff;
rom[69627] = 12'hfff;
rom[69628] = 12'hfff;
rom[69629] = 12'hfff;
rom[69630] = 12'hfff;
rom[69631] = 12'hfff;
rom[69632] = 12'hfff;
rom[69633] = 12'hfff;
rom[69634] = 12'hfff;
rom[69635] = 12'hfff;
rom[69636] = 12'hfff;
rom[69637] = 12'hfff;
rom[69638] = 12'hfff;
rom[69639] = 12'hfff;
rom[69640] = 12'hfff;
rom[69641] = 12'hfff;
rom[69642] = 12'hfff;
rom[69643] = 12'hfff;
rom[69644] = 12'hfff;
rom[69645] = 12'hfff;
rom[69646] = 12'hfff;
rom[69647] = 12'hfff;
rom[69648] = 12'hfff;
rom[69649] = 12'hfff;
rom[69650] = 12'hfff;
rom[69651] = 12'hfff;
rom[69652] = 12'hfff;
rom[69653] = 12'hfff;
rom[69654] = 12'hfff;
rom[69655] = 12'hfff;
rom[69656] = 12'hfff;
rom[69657] = 12'hfff;
rom[69658] = 12'hfff;
rom[69659] = 12'hfff;
rom[69660] = 12'hfff;
rom[69661] = 12'hfff;
rom[69662] = 12'hfff;
rom[69663] = 12'hfff;
rom[69664] = 12'hfff;
rom[69665] = 12'hfff;
rom[69666] = 12'hfff;
rom[69667] = 12'hfff;
rom[69668] = 12'hfff;
rom[69669] = 12'hfff;
rom[69670] = 12'hfff;
rom[69671] = 12'hfff;
rom[69672] = 12'hfff;
rom[69673] = 12'hfff;
rom[69674] = 12'hfff;
rom[69675] = 12'hfff;
rom[69676] = 12'hfff;
rom[69677] = 12'hfff;
rom[69678] = 12'hfff;
rom[69679] = 12'hfff;
rom[69680] = 12'hfff;
rom[69681] = 12'hfff;
rom[69682] = 12'hfff;
rom[69683] = 12'hfff;
rom[69684] = 12'hfff;
rom[69685] = 12'hfff;
rom[69686] = 12'hfff;
rom[69687] = 12'hfff;
rom[69688] = 12'hfff;
rom[69689] = 12'hfff;
rom[69690] = 12'hfff;
rom[69691] = 12'hfff;
rom[69692] = 12'hfff;
rom[69693] = 12'hfff;
rom[69694] = 12'hfff;
rom[69695] = 12'hfff;
rom[69696] = 12'hfff;
rom[69697] = 12'hfff;
rom[69698] = 12'hfff;
rom[69699] = 12'hfff;
rom[69700] = 12'hfff;
rom[69701] = 12'hfff;
rom[69702] = 12'hfff;
rom[69703] = 12'hfff;
rom[69704] = 12'hfff;
rom[69705] = 12'hfff;
rom[69706] = 12'hfff;
rom[69707] = 12'hfff;
rom[69708] = 12'hfff;
rom[69709] = 12'hfff;
rom[69710] = 12'heee;
rom[69711] = 12'heee;
rom[69712] = 12'hddd;
rom[69713] = 12'hccc;
rom[69714] = 12'hccc;
rom[69715] = 12'hbbb;
rom[69716] = 12'haaa;
rom[69717] = 12'haaa;
rom[69718] = 12'haaa;
rom[69719] = 12'h999;
rom[69720] = 12'h999;
rom[69721] = 12'h999;
rom[69722] = 12'h888;
rom[69723] = 12'h888;
rom[69724] = 12'h888;
rom[69725] = 12'h888;
rom[69726] = 12'h888;
rom[69727] = 12'h777;
rom[69728] = 12'h777;
rom[69729] = 12'h777;
rom[69730] = 12'h777;
rom[69731] = 12'h777;
rom[69732] = 12'h777;
rom[69733] = 12'h666;
rom[69734] = 12'h666;
rom[69735] = 12'h666;
rom[69736] = 12'h555;
rom[69737] = 12'h555;
rom[69738] = 12'h555;
rom[69739] = 12'h555;
rom[69740] = 12'h555;
rom[69741] = 12'h555;
rom[69742] = 12'h555;
rom[69743] = 12'h555;
rom[69744] = 12'h555;
rom[69745] = 12'h555;
rom[69746] = 12'h555;
rom[69747] = 12'h555;
rom[69748] = 12'h555;
rom[69749] = 12'h555;
rom[69750] = 12'h555;
rom[69751] = 12'h555;
rom[69752] = 12'h555;
rom[69753] = 12'h555;
rom[69754] = 12'h555;
rom[69755] = 12'h555;
rom[69756] = 12'h555;
rom[69757] = 12'h555;
rom[69758] = 12'h555;
rom[69759] = 12'h555;
rom[69760] = 12'h555;
rom[69761] = 12'h555;
rom[69762] = 12'h555;
rom[69763] = 12'h555;
rom[69764] = 12'h555;
rom[69765] = 12'h555;
rom[69766] = 12'h555;
rom[69767] = 12'h555;
rom[69768] = 12'h555;
rom[69769] = 12'h444;
rom[69770] = 12'h444;
rom[69771] = 12'h444;
rom[69772] = 12'h444;
rom[69773] = 12'h444;
rom[69774] = 12'h333;
rom[69775] = 12'h333;
rom[69776] = 12'h333;
rom[69777] = 12'h333;
rom[69778] = 12'h333;
rom[69779] = 12'h333;
rom[69780] = 12'h333;
rom[69781] = 12'h333;
rom[69782] = 12'h333;
rom[69783] = 12'h333;
rom[69784] = 12'h222;
rom[69785] = 12'h222;
rom[69786] = 12'h222;
rom[69787] = 12'h222;
rom[69788] = 12'h222;
rom[69789] = 12'h222;
rom[69790] = 12'h222;
rom[69791] = 12'h222;
rom[69792] = 12'h222;
rom[69793] = 12'h222;
rom[69794] = 12'h222;
rom[69795] = 12'h111;
rom[69796] = 12'h111;
rom[69797] = 12'h111;
rom[69798] = 12'h111;
rom[69799] = 12'h111;
rom[69800] = 12'h111;
rom[69801] = 12'h111;
rom[69802] = 12'h111;
rom[69803] = 12'h111;
rom[69804] = 12'h222;
rom[69805] = 12'h222;
rom[69806] = 12'h111;
rom[69807] = 12'h111;
rom[69808] = 12'h111;
rom[69809] = 12'h111;
rom[69810] = 12'h111;
rom[69811] = 12'h111;
rom[69812] = 12'h111;
rom[69813] = 12'h222;
rom[69814] = 12'h111;
rom[69815] = 12'h111;
rom[69816] = 12'h111;
rom[69817] = 12'h  0;
rom[69818] = 12'h  0;
rom[69819] = 12'h  0;
rom[69820] = 12'h  0;
rom[69821] = 12'h  0;
rom[69822] = 12'h  0;
rom[69823] = 12'h  0;
rom[69824] = 12'h  0;
rom[69825] = 12'h  0;
rom[69826] = 12'h  0;
rom[69827] = 12'h  0;
rom[69828] = 12'h  0;
rom[69829] = 12'h  0;
rom[69830] = 12'h  0;
rom[69831] = 12'h  0;
rom[69832] = 12'h  0;
rom[69833] = 12'h  0;
rom[69834] = 12'h  0;
rom[69835] = 12'h  0;
rom[69836] = 12'h  0;
rom[69837] = 12'h  0;
rom[69838] = 12'h  0;
rom[69839] = 12'h  0;
rom[69840] = 12'h  0;
rom[69841] = 12'h  0;
rom[69842] = 12'h  0;
rom[69843] = 12'h  0;
rom[69844] = 12'h  0;
rom[69845] = 12'h  0;
rom[69846] = 12'h  0;
rom[69847] = 12'h  0;
rom[69848] = 12'h  0;
rom[69849] = 12'h  0;
rom[69850] = 12'h  0;
rom[69851] = 12'h  0;
rom[69852] = 12'h  0;
rom[69853] = 12'h  0;
rom[69854] = 12'h  0;
rom[69855] = 12'h  0;
rom[69856] = 12'h  0;
rom[69857] = 12'h  0;
rom[69858] = 12'h  0;
rom[69859] = 12'h  0;
rom[69860] = 12'h  0;
rom[69861] = 12'h  0;
rom[69862] = 12'h  0;
rom[69863] = 12'h  0;
rom[69864] = 12'h  0;
rom[69865] = 12'h  0;
rom[69866] = 12'h  0;
rom[69867] = 12'h  0;
rom[69868] = 12'h  0;
rom[69869] = 12'h  0;
rom[69870] = 12'h111;
rom[69871] = 12'h111;
rom[69872] = 12'h111;
rom[69873] = 12'h222;
rom[69874] = 12'h222;
rom[69875] = 12'h222;
rom[69876] = 12'h333;
rom[69877] = 12'h333;
rom[69878] = 12'h444;
rom[69879] = 12'h555;
rom[69880] = 12'h666;
rom[69881] = 12'h555;
rom[69882] = 12'h333;
rom[69883] = 12'h222;
rom[69884] = 12'h111;
rom[69885] = 12'h111;
rom[69886] = 12'h111;
rom[69887] = 12'h  0;
rom[69888] = 12'h  0;
rom[69889] = 12'h  0;
rom[69890] = 12'h  0;
rom[69891] = 12'h  0;
rom[69892] = 12'h  0;
rom[69893] = 12'h  0;
rom[69894] = 12'h111;
rom[69895] = 12'h111;
rom[69896] = 12'h111;
rom[69897] = 12'h111;
rom[69898] = 12'h111;
rom[69899] = 12'h222;
rom[69900] = 12'h222;
rom[69901] = 12'h333;
rom[69902] = 12'h333;
rom[69903] = 12'h333;
rom[69904] = 12'h444;
rom[69905] = 12'h444;
rom[69906] = 12'h444;
rom[69907] = 12'h444;
rom[69908] = 12'h444;
rom[69909] = 12'h555;
rom[69910] = 12'h555;
rom[69911] = 12'h555;
rom[69912] = 12'h666;
rom[69913] = 12'h666;
rom[69914] = 12'h777;
rom[69915] = 12'h888;
rom[69916] = 12'h999;
rom[69917] = 12'h999;
rom[69918] = 12'haaa;
rom[69919] = 12'haaa;
rom[69920] = 12'haaa;
rom[69921] = 12'haaa;
rom[69922] = 12'haaa;
rom[69923] = 12'hbbb;
rom[69924] = 12'hbbb;
rom[69925] = 12'hbbb;
rom[69926] = 12'hbbb;
rom[69927] = 12'hbbb;
rom[69928] = 12'hccc;
rom[69929] = 12'hccc;
rom[69930] = 12'hccc;
rom[69931] = 12'hddd;
rom[69932] = 12'hddd;
rom[69933] = 12'heee;
rom[69934] = 12'heee;
rom[69935] = 12'hfff;
rom[69936] = 12'hfff;
rom[69937] = 12'hfff;
rom[69938] = 12'hfff;
rom[69939] = 12'hfff;
rom[69940] = 12'hfff;
rom[69941] = 12'hfff;
rom[69942] = 12'hfff;
rom[69943] = 12'hfff;
rom[69944] = 12'heee;
rom[69945] = 12'hddd;
rom[69946] = 12'hddd;
rom[69947] = 12'hccc;
rom[69948] = 12'hbbb;
rom[69949] = 12'hbbb;
rom[69950] = 12'haaa;
rom[69951] = 12'haaa;
rom[69952] = 12'h999;
rom[69953] = 12'h999;
rom[69954] = 12'h999;
rom[69955] = 12'h888;
rom[69956] = 12'h888;
rom[69957] = 12'h888;
rom[69958] = 12'h888;
rom[69959] = 12'h888;
rom[69960] = 12'h777;
rom[69961] = 12'h777;
rom[69962] = 12'h777;
rom[69963] = 12'h777;
rom[69964] = 12'h777;
rom[69965] = 12'h777;
rom[69966] = 12'h777;
rom[69967] = 12'h777;
rom[69968] = 12'h777;
rom[69969] = 12'h777;
rom[69970] = 12'h777;
rom[69971] = 12'h777;
rom[69972] = 12'h777;
rom[69973] = 12'h777;
rom[69974] = 12'h777;
rom[69975] = 12'h777;
rom[69976] = 12'h777;
rom[69977] = 12'h777;
rom[69978] = 12'h777;
rom[69979] = 12'h777;
rom[69980] = 12'h777;
rom[69981] = 12'h777;
rom[69982] = 12'h777;
rom[69983] = 12'h777;
rom[69984] = 12'h888;
rom[69985] = 12'h888;
rom[69986] = 12'h999;
rom[69987] = 12'haaa;
rom[69988] = 12'haaa;
rom[69989] = 12'haaa;
rom[69990] = 12'haaa;
rom[69991] = 12'haaa;
rom[69992] = 12'h999;
rom[69993] = 12'h888;
rom[69994] = 12'h888;
rom[69995] = 12'h777;
rom[69996] = 12'h666;
rom[69997] = 12'h666;
rom[69998] = 12'h666;
rom[69999] = 12'h666;
rom[70000] = 12'hfff;
rom[70001] = 12'hfff;
rom[70002] = 12'hfff;
rom[70003] = 12'hfff;
rom[70004] = 12'hfff;
rom[70005] = 12'hfff;
rom[70006] = 12'hfff;
rom[70007] = 12'hfff;
rom[70008] = 12'hfff;
rom[70009] = 12'hfff;
rom[70010] = 12'hfff;
rom[70011] = 12'hfff;
rom[70012] = 12'hfff;
rom[70013] = 12'hfff;
rom[70014] = 12'hfff;
rom[70015] = 12'hfff;
rom[70016] = 12'hfff;
rom[70017] = 12'hfff;
rom[70018] = 12'hfff;
rom[70019] = 12'hfff;
rom[70020] = 12'hfff;
rom[70021] = 12'hfff;
rom[70022] = 12'hfff;
rom[70023] = 12'hfff;
rom[70024] = 12'hfff;
rom[70025] = 12'hfff;
rom[70026] = 12'hfff;
rom[70027] = 12'hfff;
rom[70028] = 12'hfff;
rom[70029] = 12'hfff;
rom[70030] = 12'hfff;
rom[70031] = 12'hfff;
rom[70032] = 12'hfff;
rom[70033] = 12'hfff;
rom[70034] = 12'hfff;
rom[70035] = 12'hfff;
rom[70036] = 12'hfff;
rom[70037] = 12'hfff;
rom[70038] = 12'hfff;
rom[70039] = 12'hfff;
rom[70040] = 12'hfff;
rom[70041] = 12'hfff;
rom[70042] = 12'hfff;
rom[70043] = 12'hfff;
rom[70044] = 12'hfff;
rom[70045] = 12'hfff;
rom[70046] = 12'hfff;
rom[70047] = 12'hfff;
rom[70048] = 12'hfff;
rom[70049] = 12'hfff;
rom[70050] = 12'hfff;
rom[70051] = 12'hfff;
rom[70052] = 12'hfff;
rom[70053] = 12'hfff;
rom[70054] = 12'hfff;
rom[70055] = 12'hfff;
rom[70056] = 12'hfff;
rom[70057] = 12'hfff;
rom[70058] = 12'hfff;
rom[70059] = 12'hfff;
rom[70060] = 12'hfff;
rom[70061] = 12'hfff;
rom[70062] = 12'hfff;
rom[70063] = 12'hfff;
rom[70064] = 12'hfff;
rom[70065] = 12'hfff;
rom[70066] = 12'hfff;
rom[70067] = 12'hfff;
rom[70068] = 12'hfff;
rom[70069] = 12'hfff;
rom[70070] = 12'hfff;
rom[70071] = 12'hfff;
rom[70072] = 12'hfff;
rom[70073] = 12'hfff;
rom[70074] = 12'hfff;
rom[70075] = 12'hfff;
rom[70076] = 12'hfff;
rom[70077] = 12'hfff;
rom[70078] = 12'hfff;
rom[70079] = 12'hfff;
rom[70080] = 12'hfff;
rom[70081] = 12'hfff;
rom[70082] = 12'hfff;
rom[70083] = 12'hfff;
rom[70084] = 12'hfff;
rom[70085] = 12'hfff;
rom[70086] = 12'hfff;
rom[70087] = 12'hfff;
rom[70088] = 12'hfff;
rom[70089] = 12'hfff;
rom[70090] = 12'hfff;
rom[70091] = 12'hfff;
rom[70092] = 12'hfff;
rom[70093] = 12'hfff;
rom[70094] = 12'hfff;
rom[70095] = 12'hfff;
rom[70096] = 12'hfff;
rom[70097] = 12'hfff;
rom[70098] = 12'hfff;
rom[70099] = 12'hfff;
rom[70100] = 12'hfff;
rom[70101] = 12'hfff;
rom[70102] = 12'hfff;
rom[70103] = 12'hfff;
rom[70104] = 12'hfff;
rom[70105] = 12'hfff;
rom[70106] = 12'hfff;
rom[70107] = 12'hfff;
rom[70108] = 12'hfff;
rom[70109] = 12'hfff;
rom[70110] = 12'heee;
rom[70111] = 12'heee;
rom[70112] = 12'hddd;
rom[70113] = 12'hccc;
rom[70114] = 12'hbbb;
rom[70115] = 12'hbbb;
rom[70116] = 12'haaa;
rom[70117] = 12'haaa;
rom[70118] = 12'haaa;
rom[70119] = 12'h999;
rom[70120] = 12'h999;
rom[70121] = 12'h888;
rom[70122] = 12'h888;
rom[70123] = 12'h888;
rom[70124] = 12'h888;
rom[70125] = 12'h888;
rom[70126] = 12'h777;
rom[70127] = 12'h777;
rom[70128] = 12'h777;
rom[70129] = 12'h777;
rom[70130] = 12'h777;
rom[70131] = 12'h777;
rom[70132] = 12'h777;
rom[70133] = 12'h666;
rom[70134] = 12'h666;
rom[70135] = 12'h666;
rom[70136] = 12'h555;
rom[70137] = 12'h555;
rom[70138] = 12'h555;
rom[70139] = 12'h555;
rom[70140] = 12'h555;
rom[70141] = 12'h555;
rom[70142] = 12'h555;
rom[70143] = 12'h555;
rom[70144] = 12'h444;
rom[70145] = 12'h444;
rom[70146] = 12'h444;
rom[70147] = 12'h444;
rom[70148] = 12'h444;
rom[70149] = 12'h444;
rom[70150] = 12'h555;
rom[70151] = 12'h555;
rom[70152] = 12'h555;
rom[70153] = 12'h555;
rom[70154] = 12'h555;
rom[70155] = 12'h555;
rom[70156] = 12'h555;
rom[70157] = 12'h555;
rom[70158] = 12'h555;
rom[70159] = 12'h555;
rom[70160] = 12'h555;
rom[70161] = 12'h555;
rom[70162] = 12'h555;
rom[70163] = 12'h555;
rom[70164] = 12'h555;
rom[70165] = 12'h555;
rom[70166] = 12'h555;
rom[70167] = 12'h555;
rom[70168] = 12'h555;
rom[70169] = 12'h444;
rom[70170] = 12'h444;
rom[70171] = 12'h444;
rom[70172] = 12'h444;
rom[70173] = 12'h333;
rom[70174] = 12'h333;
rom[70175] = 12'h333;
rom[70176] = 12'h333;
rom[70177] = 12'h333;
rom[70178] = 12'h333;
rom[70179] = 12'h333;
rom[70180] = 12'h333;
rom[70181] = 12'h333;
rom[70182] = 12'h333;
rom[70183] = 12'h333;
rom[70184] = 12'h333;
rom[70185] = 12'h333;
rom[70186] = 12'h222;
rom[70187] = 12'h222;
rom[70188] = 12'h222;
rom[70189] = 12'h222;
rom[70190] = 12'h222;
rom[70191] = 12'h222;
rom[70192] = 12'h222;
rom[70193] = 12'h222;
rom[70194] = 12'h222;
rom[70195] = 12'h222;
rom[70196] = 12'h111;
rom[70197] = 12'h111;
rom[70198] = 12'h111;
rom[70199] = 12'h111;
rom[70200] = 12'h111;
rom[70201] = 12'h111;
rom[70202] = 12'h111;
rom[70203] = 12'h222;
rom[70204] = 12'h222;
rom[70205] = 12'h222;
rom[70206] = 12'h111;
rom[70207] = 12'h111;
rom[70208] = 12'h111;
rom[70209] = 12'h111;
rom[70210] = 12'h111;
rom[70211] = 12'h111;
rom[70212] = 12'h222;
rom[70213] = 12'h222;
rom[70214] = 12'h111;
rom[70215] = 12'h111;
rom[70216] = 12'h  0;
rom[70217] = 12'h  0;
rom[70218] = 12'h  0;
rom[70219] = 12'h  0;
rom[70220] = 12'h  0;
rom[70221] = 12'h  0;
rom[70222] = 12'h  0;
rom[70223] = 12'h  0;
rom[70224] = 12'h  0;
rom[70225] = 12'h  0;
rom[70226] = 12'h  0;
rom[70227] = 12'h  0;
rom[70228] = 12'h  0;
rom[70229] = 12'h  0;
rom[70230] = 12'h  0;
rom[70231] = 12'h  0;
rom[70232] = 12'h  0;
rom[70233] = 12'h  0;
rom[70234] = 12'h  0;
rom[70235] = 12'h  0;
rom[70236] = 12'h  0;
rom[70237] = 12'h  0;
rom[70238] = 12'h  0;
rom[70239] = 12'h  0;
rom[70240] = 12'h  0;
rom[70241] = 12'h  0;
rom[70242] = 12'h  0;
rom[70243] = 12'h  0;
rom[70244] = 12'h  0;
rom[70245] = 12'h  0;
rom[70246] = 12'h  0;
rom[70247] = 12'h  0;
rom[70248] = 12'h  0;
rom[70249] = 12'h  0;
rom[70250] = 12'h  0;
rom[70251] = 12'h  0;
rom[70252] = 12'h  0;
rom[70253] = 12'h  0;
rom[70254] = 12'h  0;
rom[70255] = 12'h  0;
rom[70256] = 12'h  0;
rom[70257] = 12'h  0;
rom[70258] = 12'h  0;
rom[70259] = 12'h  0;
rom[70260] = 12'h  0;
rom[70261] = 12'h  0;
rom[70262] = 12'h  0;
rom[70263] = 12'h  0;
rom[70264] = 12'h  0;
rom[70265] = 12'h  0;
rom[70266] = 12'h  0;
rom[70267] = 12'h  0;
rom[70268] = 12'h  0;
rom[70269] = 12'h  0;
rom[70270] = 12'h111;
rom[70271] = 12'h111;
rom[70272] = 12'h111;
rom[70273] = 12'h222;
rom[70274] = 12'h222;
rom[70275] = 12'h222;
rom[70276] = 12'h222;
rom[70277] = 12'h333;
rom[70278] = 12'h444;
rom[70279] = 12'h555;
rom[70280] = 12'h666;
rom[70281] = 12'h555;
rom[70282] = 12'h333;
rom[70283] = 12'h222;
rom[70284] = 12'h111;
rom[70285] = 12'h111;
rom[70286] = 12'h  0;
rom[70287] = 12'h  0;
rom[70288] = 12'h  0;
rom[70289] = 12'h  0;
rom[70290] = 12'h  0;
rom[70291] = 12'h  0;
rom[70292] = 12'h  0;
rom[70293] = 12'h  0;
rom[70294] = 12'h  0;
rom[70295] = 12'h111;
rom[70296] = 12'h111;
rom[70297] = 12'h111;
rom[70298] = 12'h111;
rom[70299] = 12'h111;
rom[70300] = 12'h222;
rom[70301] = 12'h222;
rom[70302] = 12'h333;
rom[70303] = 12'h333;
rom[70304] = 12'h444;
rom[70305] = 12'h444;
rom[70306] = 12'h444;
rom[70307] = 12'h444;
rom[70308] = 12'h444;
rom[70309] = 12'h555;
rom[70310] = 12'h555;
rom[70311] = 12'h555;
rom[70312] = 12'h666;
rom[70313] = 12'h777;
rom[70314] = 12'h777;
rom[70315] = 12'h888;
rom[70316] = 12'h999;
rom[70317] = 12'h999;
rom[70318] = 12'haaa;
rom[70319] = 12'haaa;
rom[70320] = 12'haaa;
rom[70321] = 12'haaa;
rom[70322] = 12'hbbb;
rom[70323] = 12'hbbb;
rom[70324] = 12'hbbb;
rom[70325] = 12'hbbb;
rom[70326] = 12'hccc;
rom[70327] = 12'hccc;
rom[70328] = 12'hccc;
rom[70329] = 12'hccc;
rom[70330] = 12'hccc;
rom[70331] = 12'hddd;
rom[70332] = 12'hddd;
rom[70333] = 12'heee;
rom[70334] = 12'hfff;
rom[70335] = 12'hfff;
rom[70336] = 12'hfff;
rom[70337] = 12'hfff;
rom[70338] = 12'hfff;
rom[70339] = 12'hfff;
rom[70340] = 12'hfff;
rom[70341] = 12'hfff;
rom[70342] = 12'hfff;
rom[70343] = 12'hfff;
rom[70344] = 12'hddd;
rom[70345] = 12'hddd;
rom[70346] = 12'hccc;
rom[70347] = 12'hbbb;
rom[70348] = 12'hbbb;
rom[70349] = 12'haaa;
rom[70350] = 12'haaa;
rom[70351] = 12'h999;
rom[70352] = 12'h999;
rom[70353] = 12'h999;
rom[70354] = 12'h888;
rom[70355] = 12'h888;
rom[70356] = 12'h888;
rom[70357] = 12'h888;
rom[70358] = 12'h888;
rom[70359] = 12'h777;
rom[70360] = 12'h777;
rom[70361] = 12'h777;
rom[70362] = 12'h777;
rom[70363] = 12'h777;
rom[70364] = 12'h666;
rom[70365] = 12'h666;
rom[70366] = 12'h666;
rom[70367] = 12'h666;
rom[70368] = 12'h666;
rom[70369] = 12'h666;
rom[70370] = 12'h666;
rom[70371] = 12'h666;
rom[70372] = 12'h666;
rom[70373] = 12'h777;
rom[70374] = 12'h777;
rom[70375] = 12'h777;
rom[70376] = 12'h777;
rom[70377] = 12'h777;
rom[70378] = 12'h777;
rom[70379] = 12'h777;
rom[70380] = 12'h777;
rom[70381] = 12'h777;
rom[70382] = 12'h777;
rom[70383] = 12'h777;
rom[70384] = 12'h777;
rom[70385] = 12'h888;
rom[70386] = 12'h888;
rom[70387] = 12'h999;
rom[70388] = 12'h999;
rom[70389] = 12'haaa;
rom[70390] = 12'haaa;
rom[70391] = 12'haaa;
rom[70392] = 12'haaa;
rom[70393] = 12'h999;
rom[70394] = 12'h888;
rom[70395] = 12'h888;
rom[70396] = 12'h777;
rom[70397] = 12'h777;
rom[70398] = 12'h777;
rom[70399] = 12'h777;
rom[70400] = 12'hfff;
rom[70401] = 12'hfff;
rom[70402] = 12'hfff;
rom[70403] = 12'hfff;
rom[70404] = 12'hfff;
rom[70405] = 12'hfff;
rom[70406] = 12'hfff;
rom[70407] = 12'hfff;
rom[70408] = 12'hfff;
rom[70409] = 12'hfff;
rom[70410] = 12'hfff;
rom[70411] = 12'hfff;
rom[70412] = 12'hfff;
rom[70413] = 12'hfff;
rom[70414] = 12'hfff;
rom[70415] = 12'hfff;
rom[70416] = 12'hfff;
rom[70417] = 12'hfff;
rom[70418] = 12'hfff;
rom[70419] = 12'hfff;
rom[70420] = 12'hfff;
rom[70421] = 12'hfff;
rom[70422] = 12'hfff;
rom[70423] = 12'hfff;
rom[70424] = 12'hfff;
rom[70425] = 12'hfff;
rom[70426] = 12'hfff;
rom[70427] = 12'hfff;
rom[70428] = 12'hfff;
rom[70429] = 12'hfff;
rom[70430] = 12'hfff;
rom[70431] = 12'hfff;
rom[70432] = 12'hfff;
rom[70433] = 12'hfff;
rom[70434] = 12'hfff;
rom[70435] = 12'hfff;
rom[70436] = 12'hfff;
rom[70437] = 12'hfff;
rom[70438] = 12'hfff;
rom[70439] = 12'hfff;
rom[70440] = 12'hfff;
rom[70441] = 12'hfff;
rom[70442] = 12'hfff;
rom[70443] = 12'hfff;
rom[70444] = 12'hfff;
rom[70445] = 12'hfff;
rom[70446] = 12'hfff;
rom[70447] = 12'hfff;
rom[70448] = 12'hfff;
rom[70449] = 12'hfff;
rom[70450] = 12'hfff;
rom[70451] = 12'hfff;
rom[70452] = 12'hfff;
rom[70453] = 12'hfff;
rom[70454] = 12'hfff;
rom[70455] = 12'hfff;
rom[70456] = 12'hfff;
rom[70457] = 12'hfff;
rom[70458] = 12'hfff;
rom[70459] = 12'hfff;
rom[70460] = 12'hfff;
rom[70461] = 12'hfff;
rom[70462] = 12'hfff;
rom[70463] = 12'hfff;
rom[70464] = 12'hfff;
rom[70465] = 12'hfff;
rom[70466] = 12'hfff;
rom[70467] = 12'hfff;
rom[70468] = 12'hfff;
rom[70469] = 12'hfff;
rom[70470] = 12'hfff;
rom[70471] = 12'hfff;
rom[70472] = 12'hfff;
rom[70473] = 12'hfff;
rom[70474] = 12'hfff;
rom[70475] = 12'hfff;
rom[70476] = 12'hfff;
rom[70477] = 12'hfff;
rom[70478] = 12'hfff;
rom[70479] = 12'hfff;
rom[70480] = 12'hfff;
rom[70481] = 12'hfff;
rom[70482] = 12'hfff;
rom[70483] = 12'hfff;
rom[70484] = 12'hfff;
rom[70485] = 12'hfff;
rom[70486] = 12'hfff;
rom[70487] = 12'hfff;
rom[70488] = 12'hfff;
rom[70489] = 12'hfff;
rom[70490] = 12'hfff;
rom[70491] = 12'hfff;
rom[70492] = 12'hfff;
rom[70493] = 12'hfff;
rom[70494] = 12'hfff;
rom[70495] = 12'hfff;
rom[70496] = 12'hfff;
rom[70497] = 12'hfff;
rom[70498] = 12'hfff;
rom[70499] = 12'hfff;
rom[70500] = 12'hfff;
rom[70501] = 12'hfff;
rom[70502] = 12'hfff;
rom[70503] = 12'hfff;
rom[70504] = 12'hfff;
rom[70505] = 12'hfff;
rom[70506] = 12'hfff;
rom[70507] = 12'hfff;
rom[70508] = 12'hfff;
rom[70509] = 12'hfff;
rom[70510] = 12'heee;
rom[70511] = 12'hddd;
rom[70512] = 12'hddd;
rom[70513] = 12'hccc;
rom[70514] = 12'hccc;
rom[70515] = 12'hbbb;
rom[70516] = 12'hbbb;
rom[70517] = 12'haaa;
rom[70518] = 12'h999;
rom[70519] = 12'h999;
rom[70520] = 12'h888;
rom[70521] = 12'h888;
rom[70522] = 12'h888;
rom[70523] = 12'h888;
rom[70524] = 12'h777;
rom[70525] = 12'h777;
rom[70526] = 12'h777;
rom[70527] = 12'h777;
rom[70528] = 12'h777;
rom[70529] = 12'h777;
rom[70530] = 12'h777;
rom[70531] = 12'h666;
rom[70532] = 12'h666;
rom[70533] = 12'h666;
rom[70534] = 12'h666;
rom[70535] = 12'h666;
rom[70536] = 12'h666;
rom[70537] = 12'h555;
rom[70538] = 12'h555;
rom[70539] = 12'h444;
rom[70540] = 12'h444;
rom[70541] = 12'h444;
rom[70542] = 12'h444;
rom[70543] = 12'h444;
rom[70544] = 12'h444;
rom[70545] = 12'h444;
rom[70546] = 12'h444;
rom[70547] = 12'h444;
rom[70548] = 12'h444;
rom[70549] = 12'h444;
rom[70550] = 12'h444;
rom[70551] = 12'h555;
rom[70552] = 12'h555;
rom[70553] = 12'h555;
rom[70554] = 12'h555;
rom[70555] = 12'h555;
rom[70556] = 12'h555;
rom[70557] = 12'h555;
rom[70558] = 12'h555;
rom[70559] = 12'h555;
rom[70560] = 12'h555;
rom[70561] = 12'h555;
rom[70562] = 12'h555;
rom[70563] = 12'h555;
rom[70564] = 12'h555;
rom[70565] = 12'h555;
rom[70566] = 12'h555;
rom[70567] = 12'h555;
rom[70568] = 12'h555;
rom[70569] = 12'h555;
rom[70570] = 12'h555;
rom[70571] = 12'h444;
rom[70572] = 12'h444;
rom[70573] = 12'h444;
rom[70574] = 12'h333;
rom[70575] = 12'h333;
rom[70576] = 12'h333;
rom[70577] = 12'h333;
rom[70578] = 12'h333;
rom[70579] = 12'h333;
rom[70580] = 12'h333;
rom[70581] = 12'h333;
rom[70582] = 12'h333;
rom[70583] = 12'h333;
rom[70584] = 12'h333;
rom[70585] = 12'h333;
rom[70586] = 12'h333;
rom[70587] = 12'h222;
rom[70588] = 12'h222;
rom[70589] = 12'h222;
rom[70590] = 12'h222;
rom[70591] = 12'h222;
rom[70592] = 12'h222;
rom[70593] = 12'h222;
rom[70594] = 12'h222;
rom[70595] = 12'h222;
rom[70596] = 12'h222;
rom[70597] = 12'h111;
rom[70598] = 12'h111;
rom[70599] = 12'h111;
rom[70600] = 12'h111;
rom[70601] = 12'h222;
rom[70602] = 12'h222;
rom[70603] = 12'h222;
rom[70604] = 12'h222;
rom[70605] = 12'h222;
rom[70606] = 12'h111;
rom[70607] = 12'h111;
rom[70608] = 12'h111;
rom[70609] = 12'h111;
rom[70610] = 12'h111;
rom[70611] = 12'h222;
rom[70612] = 12'h222;
rom[70613] = 12'h222;
rom[70614] = 12'h111;
rom[70615] = 12'h111;
rom[70616] = 12'h  0;
rom[70617] = 12'h  0;
rom[70618] = 12'h  0;
rom[70619] = 12'h  0;
rom[70620] = 12'h  0;
rom[70621] = 12'h  0;
rom[70622] = 12'h  0;
rom[70623] = 12'h  0;
rom[70624] = 12'h  0;
rom[70625] = 12'h  0;
rom[70626] = 12'h  0;
rom[70627] = 12'h  0;
rom[70628] = 12'h  0;
rom[70629] = 12'h  0;
rom[70630] = 12'h  0;
rom[70631] = 12'h  0;
rom[70632] = 12'h  0;
rom[70633] = 12'h  0;
rom[70634] = 12'h  0;
rom[70635] = 12'h  0;
rom[70636] = 12'h  0;
rom[70637] = 12'h  0;
rom[70638] = 12'h  0;
rom[70639] = 12'h  0;
rom[70640] = 12'h  0;
rom[70641] = 12'h  0;
rom[70642] = 12'h  0;
rom[70643] = 12'h  0;
rom[70644] = 12'h  0;
rom[70645] = 12'h  0;
rom[70646] = 12'h  0;
rom[70647] = 12'h  0;
rom[70648] = 12'h  0;
rom[70649] = 12'h  0;
rom[70650] = 12'h  0;
rom[70651] = 12'h  0;
rom[70652] = 12'h  0;
rom[70653] = 12'h  0;
rom[70654] = 12'h  0;
rom[70655] = 12'h  0;
rom[70656] = 12'h  0;
rom[70657] = 12'h  0;
rom[70658] = 12'h  0;
rom[70659] = 12'h  0;
rom[70660] = 12'h  0;
rom[70661] = 12'h  0;
rom[70662] = 12'h  0;
rom[70663] = 12'h  0;
rom[70664] = 12'h  0;
rom[70665] = 12'h  0;
rom[70666] = 12'h  0;
rom[70667] = 12'h  0;
rom[70668] = 12'h  0;
rom[70669] = 12'h  0;
rom[70670] = 12'h111;
rom[70671] = 12'h111;
rom[70672] = 12'h222;
rom[70673] = 12'h222;
rom[70674] = 12'h222;
rom[70675] = 12'h222;
rom[70676] = 12'h333;
rom[70677] = 12'h444;
rom[70678] = 12'h555;
rom[70679] = 12'h555;
rom[70680] = 12'h666;
rom[70681] = 12'h444;
rom[70682] = 12'h222;
rom[70683] = 12'h111;
rom[70684] = 12'h111;
rom[70685] = 12'h111;
rom[70686] = 12'h  0;
rom[70687] = 12'h  0;
rom[70688] = 12'h  0;
rom[70689] = 12'h  0;
rom[70690] = 12'h  0;
rom[70691] = 12'h  0;
rom[70692] = 12'h  0;
rom[70693] = 12'h  0;
rom[70694] = 12'h  0;
rom[70695] = 12'h111;
rom[70696] = 12'h111;
rom[70697] = 12'h111;
rom[70698] = 12'h111;
rom[70699] = 12'h222;
rom[70700] = 12'h222;
rom[70701] = 12'h222;
rom[70702] = 12'h333;
rom[70703] = 12'h333;
rom[70704] = 12'h444;
rom[70705] = 12'h444;
rom[70706] = 12'h444;
rom[70707] = 12'h444;
rom[70708] = 12'h444;
rom[70709] = 12'h555;
rom[70710] = 12'h555;
rom[70711] = 12'h555;
rom[70712] = 12'h666;
rom[70713] = 12'h777;
rom[70714] = 12'h777;
rom[70715] = 12'h888;
rom[70716] = 12'h999;
rom[70717] = 12'haaa;
rom[70718] = 12'haaa;
rom[70719] = 12'haaa;
rom[70720] = 12'hbbb;
rom[70721] = 12'hbbb;
rom[70722] = 12'hbbb;
rom[70723] = 12'hbbb;
rom[70724] = 12'hbbb;
rom[70725] = 12'hbbb;
rom[70726] = 12'hccc;
rom[70727] = 12'hccc;
rom[70728] = 12'hccc;
rom[70729] = 12'hccc;
rom[70730] = 12'hddd;
rom[70731] = 12'hddd;
rom[70732] = 12'heee;
rom[70733] = 12'hfff;
rom[70734] = 12'hfff;
rom[70735] = 12'hfff;
rom[70736] = 12'hfff;
rom[70737] = 12'hfff;
rom[70738] = 12'hfff;
rom[70739] = 12'hfff;
rom[70740] = 12'hfff;
rom[70741] = 12'hfff;
rom[70742] = 12'heee;
rom[70743] = 12'heee;
rom[70744] = 12'hddd;
rom[70745] = 12'hccc;
rom[70746] = 12'hbbb;
rom[70747] = 12'hbbb;
rom[70748] = 12'haaa;
rom[70749] = 12'haaa;
rom[70750] = 12'haaa;
rom[70751] = 12'h999;
rom[70752] = 12'h999;
rom[70753] = 12'h999;
rom[70754] = 12'h888;
rom[70755] = 12'h888;
rom[70756] = 12'h888;
rom[70757] = 12'h888;
rom[70758] = 12'h777;
rom[70759] = 12'h777;
rom[70760] = 12'h666;
rom[70761] = 12'h666;
rom[70762] = 12'h666;
rom[70763] = 12'h666;
rom[70764] = 12'h666;
rom[70765] = 12'h666;
rom[70766] = 12'h666;
rom[70767] = 12'h666;
rom[70768] = 12'h666;
rom[70769] = 12'h666;
rom[70770] = 12'h666;
rom[70771] = 12'h666;
rom[70772] = 12'h666;
rom[70773] = 12'h666;
rom[70774] = 12'h666;
rom[70775] = 12'h666;
rom[70776] = 12'h666;
rom[70777] = 12'h666;
rom[70778] = 12'h777;
rom[70779] = 12'h777;
rom[70780] = 12'h777;
rom[70781] = 12'h777;
rom[70782] = 12'h777;
rom[70783] = 12'h777;
rom[70784] = 12'h777;
rom[70785] = 12'h777;
rom[70786] = 12'h888;
rom[70787] = 12'h888;
rom[70788] = 12'h888;
rom[70789] = 12'h999;
rom[70790] = 12'h999;
rom[70791] = 12'h999;
rom[70792] = 12'h999;
rom[70793] = 12'h999;
rom[70794] = 12'h999;
rom[70795] = 12'h999;
rom[70796] = 12'h888;
rom[70797] = 12'h888;
rom[70798] = 12'h888;
rom[70799] = 12'h777;
rom[70800] = 12'hfff;
rom[70801] = 12'hfff;
rom[70802] = 12'hfff;
rom[70803] = 12'hfff;
rom[70804] = 12'hfff;
rom[70805] = 12'hfff;
rom[70806] = 12'hfff;
rom[70807] = 12'hfff;
rom[70808] = 12'hfff;
rom[70809] = 12'hfff;
rom[70810] = 12'hfff;
rom[70811] = 12'hfff;
rom[70812] = 12'hfff;
rom[70813] = 12'hfff;
rom[70814] = 12'hfff;
rom[70815] = 12'hfff;
rom[70816] = 12'hfff;
rom[70817] = 12'hfff;
rom[70818] = 12'hfff;
rom[70819] = 12'hfff;
rom[70820] = 12'hfff;
rom[70821] = 12'hfff;
rom[70822] = 12'hfff;
rom[70823] = 12'hfff;
rom[70824] = 12'hfff;
rom[70825] = 12'hfff;
rom[70826] = 12'hfff;
rom[70827] = 12'hfff;
rom[70828] = 12'hfff;
rom[70829] = 12'hfff;
rom[70830] = 12'hfff;
rom[70831] = 12'hfff;
rom[70832] = 12'hfff;
rom[70833] = 12'hfff;
rom[70834] = 12'hfff;
rom[70835] = 12'hfff;
rom[70836] = 12'hfff;
rom[70837] = 12'hfff;
rom[70838] = 12'hfff;
rom[70839] = 12'hfff;
rom[70840] = 12'hfff;
rom[70841] = 12'hfff;
rom[70842] = 12'hfff;
rom[70843] = 12'hfff;
rom[70844] = 12'hfff;
rom[70845] = 12'hfff;
rom[70846] = 12'hfff;
rom[70847] = 12'hfff;
rom[70848] = 12'hfff;
rom[70849] = 12'hfff;
rom[70850] = 12'hfff;
rom[70851] = 12'hfff;
rom[70852] = 12'hfff;
rom[70853] = 12'hfff;
rom[70854] = 12'hfff;
rom[70855] = 12'hfff;
rom[70856] = 12'hfff;
rom[70857] = 12'hfff;
rom[70858] = 12'hfff;
rom[70859] = 12'hfff;
rom[70860] = 12'hfff;
rom[70861] = 12'hfff;
rom[70862] = 12'hfff;
rom[70863] = 12'hfff;
rom[70864] = 12'hfff;
rom[70865] = 12'hfff;
rom[70866] = 12'hfff;
rom[70867] = 12'hfff;
rom[70868] = 12'hfff;
rom[70869] = 12'hfff;
rom[70870] = 12'hfff;
rom[70871] = 12'hfff;
rom[70872] = 12'hfff;
rom[70873] = 12'hfff;
rom[70874] = 12'hfff;
rom[70875] = 12'hfff;
rom[70876] = 12'hfff;
rom[70877] = 12'hfff;
rom[70878] = 12'hfff;
rom[70879] = 12'hfff;
rom[70880] = 12'hfff;
rom[70881] = 12'hfff;
rom[70882] = 12'hfff;
rom[70883] = 12'hfff;
rom[70884] = 12'hfff;
rom[70885] = 12'hfff;
rom[70886] = 12'hfff;
rom[70887] = 12'hfff;
rom[70888] = 12'hfff;
rom[70889] = 12'hfff;
rom[70890] = 12'hfff;
rom[70891] = 12'hfff;
rom[70892] = 12'hfff;
rom[70893] = 12'hfff;
rom[70894] = 12'hfff;
rom[70895] = 12'hfff;
rom[70896] = 12'hfff;
rom[70897] = 12'hfff;
rom[70898] = 12'hfff;
rom[70899] = 12'hfff;
rom[70900] = 12'hfff;
rom[70901] = 12'hfff;
rom[70902] = 12'hfff;
rom[70903] = 12'hfff;
rom[70904] = 12'hfff;
rom[70905] = 12'hfff;
rom[70906] = 12'hfff;
rom[70907] = 12'hfff;
rom[70908] = 12'hfff;
rom[70909] = 12'hfff;
rom[70910] = 12'heee;
rom[70911] = 12'hddd;
rom[70912] = 12'hccc;
rom[70913] = 12'hccc;
rom[70914] = 12'hccc;
rom[70915] = 12'hbbb;
rom[70916] = 12'hbbb;
rom[70917] = 12'haaa;
rom[70918] = 12'haaa;
rom[70919] = 12'h999;
rom[70920] = 12'h999;
rom[70921] = 12'h888;
rom[70922] = 12'h888;
rom[70923] = 12'h888;
rom[70924] = 12'h888;
rom[70925] = 12'h777;
rom[70926] = 12'h777;
rom[70927] = 12'h777;
rom[70928] = 12'h777;
rom[70929] = 12'h777;
rom[70930] = 12'h777;
rom[70931] = 12'h777;
rom[70932] = 12'h666;
rom[70933] = 12'h666;
rom[70934] = 12'h666;
rom[70935] = 12'h666;
rom[70936] = 12'h666;
rom[70937] = 12'h555;
rom[70938] = 12'h555;
rom[70939] = 12'h444;
rom[70940] = 12'h444;
rom[70941] = 12'h444;
rom[70942] = 12'h444;
rom[70943] = 12'h444;
rom[70944] = 12'h444;
rom[70945] = 12'h444;
rom[70946] = 12'h444;
rom[70947] = 12'h444;
rom[70948] = 12'h444;
rom[70949] = 12'h444;
rom[70950] = 12'h444;
rom[70951] = 12'h444;
rom[70952] = 12'h555;
rom[70953] = 12'h555;
rom[70954] = 12'h555;
rom[70955] = 12'h555;
rom[70956] = 12'h555;
rom[70957] = 12'h555;
rom[70958] = 12'h555;
rom[70959] = 12'h555;
rom[70960] = 12'h555;
rom[70961] = 12'h555;
rom[70962] = 12'h555;
rom[70963] = 12'h555;
rom[70964] = 12'h555;
rom[70965] = 12'h555;
rom[70966] = 12'h555;
rom[70967] = 12'h555;
rom[70968] = 12'h555;
rom[70969] = 12'h555;
rom[70970] = 12'h555;
rom[70971] = 12'h555;
rom[70972] = 12'h555;
rom[70973] = 12'h444;
rom[70974] = 12'h444;
rom[70975] = 12'h444;
rom[70976] = 12'h333;
rom[70977] = 12'h333;
rom[70978] = 12'h333;
rom[70979] = 12'h333;
rom[70980] = 12'h333;
rom[70981] = 12'h333;
rom[70982] = 12'h333;
rom[70983] = 12'h333;
rom[70984] = 12'h333;
rom[70985] = 12'h333;
rom[70986] = 12'h333;
rom[70987] = 12'h333;
rom[70988] = 12'h333;
rom[70989] = 12'h222;
rom[70990] = 12'h222;
rom[70991] = 12'h222;
rom[70992] = 12'h333;
rom[70993] = 12'h222;
rom[70994] = 12'h333;
rom[70995] = 12'h333;
rom[70996] = 12'h222;
rom[70997] = 12'h111;
rom[70998] = 12'h111;
rom[70999] = 12'h111;
rom[71000] = 12'h111;
rom[71001] = 12'h222;
rom[71002] = 12'h222;
rom[71003] = 12'h222;
rom[71004] = 12'h222;
rom[71005] = 12'h222;
rom[71006] = 12'h111;
rom[71007] = 12'h111;
rom[71008] = 12'h111;
rom[71009] = 12'h111;
rom[71010] = 12'h222;
rom[71011] = 12'h222;
rom[71012] = 12'h222;
rom[71013] = 12'h222;
rom[71014] = 12'h111;
rom[71015] = 12'h111;
rom[71016] = 12'h  0;
rom[71017] = 12'h  0;
rom[71018] = 12'h  0;
rom[71019] = 12'h  0;
rom[71020] = 12'h  0;
rom[71021] = 12'h  0;
rom[71022] = 12'h  0;
rom[71023] = 12'h  0;
rom[71024] = 12'h  0;
rom[71025] = 12'h  0;
rom[71026] = 12'h  0;
rom[71027] = 12'h  0;
rom[71028] = 12'h  0;
rom[71029] = 12'h  0;
rom[71030] = 12'h  0;
rom[71031] = 12'h  0;
rom[71032] = 12'h  0;
rom[71033] = 12'h  0;
rom[71034] = 12'h  0;
rom[71035] = 12'h  0;
rom[71036] = 12'h  0;
rom[71037] = 12'h  0;
rom[71038] = 12'h  0;
rom[71039] = 12'h  0;
rom[71040] = 12'h  0;
rom[71041] = 12'h  0;
rom[71042] = 12'h  0;
rom[71043] = 12'h  0;
rom[71044] = 12'h  0;
rom[71045] = 12'h  0;
rom[71046] = 12'h  0;
rom[71047] = 12'h  0;
rom[71048] = 12'h  0;
rom[71049] = 12'h  0;
rom[71050] = 12'h  0;
rom[71051] = 12'h  0;
rom[71052] = 12'h  0;
rom[71053] = 12'h  0;
rom[71054] = 12'h  0;
rom[71055] = 12'h  0;
rom[71056] = 12'h  0;
rom[71057] = 12'h  0;
rom[71058] = 12'h  0;
rom[71059] = 12'h  0;
rom[71060] = 12'h  0;
rom[71061] = 12'h  0;
rom[71062] = 12'h  0;
rom[71063] = 12'h  0;
rom[71064] = 12'h  0;
rom[71065] = 12'h  0;
rom[71066] = 12'h  0;
rom[71067] = 12'h  0;
rom[71068] = 12'h  0;
rom[71069] = 12'h  0;
rom[71070] = 12'h111;
rom[71071] = 12'h111;
rom[71072] = 12'h222;
rom[71073] = 12'h222;
rom[71074] = 12'h222;
rom[71075] = 12'h222;
rom[71076] = 12'h333;
rom[71077] = 12'h444;
rom[71078] = 12'h555;
rom[71079] = 12'h555;
rom[71080] = 12'h666;
rom[71081] = 12'h444;
rom[71082] = 12'h222;
rom[71083] = 12'h111;
rom[71084] = 12'h111;
rom[71085] = 12'h111;
rom[71086] = 12'h  0;
rom[71087] = 12'h  0;
rom[71088] = 12'h  0;
rom[71089] = 12'h  0;
rom[71090] = 12'h  0;
rom[71091] = 12'h  0;
rom[71092] = 12'h  0;
rom[71093] = 12'h  0;
rom[71094] = 12'h  0;
rom[71095] = 12'h  0;
rom[71096] = 12'h111;
rom[71097] = 12'h111;
rom[71098] = 12'h111;
rom[71099] = 12'h111;
rom[71100] = 12'h222;
rom[71101] = 12'h222;
rom[71102] = 12'h333;
rom[71103] = 12'h333;
rom[71104] = 12'h444;
rom[71105] = 12'h444;
rom[71106] = 12'h444;
rom[71107] = 12'h555;
rom[71108] = 12'h555;
rom[71109] = 12'h555;
rom[71110] = 12'h555;
rom[71111] = 12'h555;
rom[71112] = 12'h666;
rom[71113] = 12'h777;
rom[71114] = 12'h777;
rom[71115] = 12'h888;
rom[71116] = 12'h999;
rom[71117] = 12'haaa;
rom[71118] = 12'haaa;
rom[71119] = 12'hbbb;
rom[71120] = 12'hbbb;
rom[71121] = 12'hbbb;
rom[71122] = 12'hbbb;
rom[71123] = 12'hbbb;
rom[71124] = 12'hbbb;
rom[71125] = 12'hbbb;
rom[71126] = 12'hccc;
rom[71127] = 12'hccc;
rom[71128] = 12'hccc;
rom[71129] = 12'hddd;
rom[71130] = 12'hddd;
rom[71131] = 12'heee;
rom[71132] = 12'hfff;
rom[71133] = 12'hfff;
rom[71134] = 12'hfff;
rom[71135] = 12'hfff;
rom[71136] = 12'hfff;
rom[71137] = 12'hfff;
rom[71138] = 12'hfff;
rom[71139] = 12'hfff;
rom[71140] = 12'hfff;
rom[71141] = 12'heee;
rom[71142] = 12'heee;
rom[71143] = 12'hddd;
rom[71144] = 12'hccc;
rom[71145] = 12'hbbb;
rom[71146] = 12'hbbb;
rom[71147] = 12'haaa;
rom[71148] = 12'haaa;
rom[71149] = 12'haaa;
rom[71150] = 12'h999;
rom[71151] = 12'h999;
rom[71152] = 12'h999;
rom[71153] = 12'h999;
rom[71154] = 12'h888;
rom[71155] = 12'h888;
rom[71156] = 12'h888;
rom[71157] = 12'h777;
rom[71158] = 12'h777;
rom[71159] = 12'h777;
rom[71160] = 12'h666;
rom[71161] = 12'h666;
rom[71162] = 12'h666;
rom[71163] = 12'h666;
rom[71164] = 12'h666;
rom[71165] = 12'h666;
rom[71166] = 12'h666;
rom[71167] = 12'h666;
rom[71168] = 12'h666;
rom[71169] = 12'h666;
rom[71170] = 12'h666;
rom[71171] = 12'h666;
rom[71172] = 12'h666;
rom[71173] = 12'h666;
rom[71174] = 12'h666;
rom[71175] = 12'h666;
rom[71176] = 12'h666;
rom[71177] = 12'h666;
rom[71178] = 12'h666;
rom[71179] = 12'h666;
rom[71180] = 12'h666;
rom[71181] = 12'h777;
rom[71182] = 12'h777;
rom[71183] = 12'h777;
rom[71184] = 12'h777;
rom[71185] = 12'h777;
rom[71186] = 12'h777;
rom[71187] = 12'h888;
rom[71188] = 12'h888;
rom[71189] = 12'h888;
rom[71190] = 12'h999;
rom[71191] = 12'h999;
rom[71192] = 12'h999;
rom[71193] = 12'h999;
rom[71194] = 12'h999;
rom[71195] = 12'h999;
rom[71196] = 12'h888;
rom[71197] = 12'h888;
rom[71198] = 12'h888;
rom[71199] = 12'h888;
rom[71200] = 12'hfff;
rom[71201] = 12'hfff;
rom[71202] = 12'hfff;
rom[71203] = 12'hfff;
rom[71204] = 12'hfff;
rom[71205] = 12'hfff;
rom[71206] = 12'hfff;
rom[71207] = 12'hfff;
rom[71208] = 12'hfff;
rom[71209] = 12'hfff;
rom[71210] = 12'hfff;
rom[71211] = 12'hfff;
rom[71212] = 12'hfff;
rom[71213] = 12'hfff;
rom[71214] = 12'hfff;
rom[71215] = 12'hfff;
rom[71216] = 12'hfff;
rom[71217] = 12'hfff;
rom[71218] = 12'hfff;
rom[71219] = 12'hfff;
rom[71220] = 12'hfff;
rom[71221] = 12'hfff;
rom[71222] = 12'hfff;
rom[71223] = 12'hfff;
rom[71224] = 12'hfff;
rom[71225] = 12'hfff;
rom[71226] = 12'hfff;
rom[71227] = 12'hfff;
rom[71228] = 12'hfff;
rom[71229] = 12'hfff;
rom[71230] = 12'hfff;
rom[71231] = 12'hfff;
rom[71232] = 12'hfff;
rom[71233] = 12'hfff;
rom[71234] = 12'hfff;
rom[71235] = 12'hfff;
rom[71236] = 12'hfff;
rom[71237] = 12'hfff;
rom[71238] = 12'hfff;
rom[71239] = 12'hfff;
rom[71240] = 12'hfff;
rom[71241] = 12'hfff;
rom[71242] = 12'hfff;
rom[71243] = 12'hfff;
rom[71244] = 12'hfff;
rom[71245] = 12'hfff;
rom[71246] = 12'hfff;
rom[71247] = 12'hfff;
rom[71248] = 12'hfff;
rom[71249] = 12'hfff;
rom[71250] = 12'hfff;
rom[71251] = 12'hfff;
rom[71252] = 12'hfff;
rom[71253] = 12'hfff;
rom[71254] = 12'hfff;
rom[71255] = 12'hfff;
rom[71256] = 12'hfff;
rom[71257] = 12'hfff;
rom[71258] = 12'hfff;
rom[71259] = 12'hfff;
rom[71260] = 12'hfff;
rom[71261] = 12'hfff;
rom[71262] = 12'hfff;
rom[71263] = 12'hfff;
rom[71264] = 12'hfff;
rom[71265] = 12'hfff;
rom[71266] = 12'hfff;
rom[71267] = 12'hfff;
rom[71268] = 12'hfff;
rom[71269] = 12'hfff;
rom[71270] = 12'hfff;
rom[71271] = 12'hfff;
rom[71272] = 12'hfff;
rom[71273] = 12'hfff;
rom[71274] = 12'hfff;
rom[71275] = 12'hfff;
rom[71276] = 12'hfff;
rom[71277] = 12'hfff;
rom[71278] = 12'hfff;
rom[71279] = 12'hfff;
rom[71280] = 12'hfff;
rom[71281] = 12'hfff;
rom[71282] = 12'hfff;
rom[71283] = 12'hfff;
rom[71284] = 12'hfff;
rom[71285] = 12'hfff;
rom[71286] = 12'hfff;
rom[71287] = 12'hfff;
rom[71288] = 12'hfff;
rom[71289] = 12'hfff;
rom[71290] = 12'hfff;
rom[71291] = 12'hfff;
rom[71292] = 12'hfff;
rom[71293] = 12'hfff;
rom[71294] = 12'hfff;
rom[71295] = 12'hfff;
rom[71296] = 12'hfff;
rom[71297] = 12'hfff;
rom[71298] = 12'hfff;
rom[71299] = 12'hfff;
rom[71300] = 12'hfff;
rom[71301] = 12'hfff;
rom[71302] = 12'hfff;
rom[71303] = 12'hfff;
rom[71304] = 12'hfff;
rom[71305] = 12'hfff;
rom[71306] = 12'hfff;
rom[71307] = 12'hfff;
rom[71308] = 12'hfff;
rom[71309] = 12'hfff;
rom[71310] = 12'heee;
rom[71311] = 12'hddd;
rom[71312] = 12'hccc;
rom[71313] = 12'hccc;
rom[71314] = 12'hccc;
rom[71315] = 12'hbbb;
rom[71316] = 12'hbbb;
rom[71317] = 12'haaa;
rom[71318] = 12'haaa;
rom[71319] = 12'haaa;
rom[71320] = 12'h999;
rom[71321] = 12'h999;
rom[71322] = 12'h888;
rom[71323] = 12'h888;
rom[71324] = 12'h888;
rom[71325] = 12'h888;
rom[71326] = 12'h777;
rom[71327] = 12'h777;
rom[71328] = 12'h777;
rom[71329] = 12'h777;
rom[71330] = 12'h777;
rom[71331] = 12'h777;
rom[71332] = 12'h777;
rom[71333] = 12'h666;
rom[71334] = 12'h666;
rom[71335] = 12'h666;
rom[71336] = 12'h666;
rom[71337] = 12'h555;
rom[71338] = 12'h555;
rom[71339] = 12'h555;
rom[71340] = 12'h444;
rom[71341] = 12'h444;
rom[71342] = 12'h444;
rom[71343] = 12'h444;
rom[71344] = 12'h444;
rom[71345] = 12'h444;
rom[71346] = 12'h444;
rom[71347] = 12'h444;
rom[71348] = 12'h444;
rom[71349] = 12'h444;
rom[71350] = 12'h444;
rom[71351] = 12'h444;
rom[71352] = 12'h444;
rom[71353] = 12'h444;
rom[71354] = 12'h555;
rom[71355] = 12'h555;
rom[71356] = 12'h555;
rom[71357] = 12'h555;
rom[71358] = 12'h555;
rom[71359] = 12'h555;
rom[71360] = 12'h555;
rom[71361] = 12'h555;
rom[71362] = 12'h555;
rom[71363] = 12'h444;
rom[71364] = 12'h444;
rom[71365] = 12'h444;
rom[71366] = 12'h555;
rom[71367] = 12'h555;
rom[71368] = 12'h555;
rom[71369] = 12'h555;
rom[71370] = 12'h555;
rom[71371] = 12'h555;
rom[71372] = 12'h555;
rom[71373] = 12'h555;
rom[71374] = 12'h444;
rom[71375] = 12'h444;
rom[71376] = 12'h444;
rom[71377] = 12'h444;
rom[71378] = 12'h333;
rom[71379] = 12'h333;
rom[71380] = 12'h333;
rom[71381] = 12'h333;
rom[71382] = 12'h333;
rom[71383] = 12'h333;
rom[71384] = 12'h333;
rom[71385] = 12'h333;
rom[71386] = 12'h333;
rom[71387] = 12'h333;
rom[71388] = 12'h333;
rom[71389] = 12'h333;
rom[71390] = 12'h222;
rom[71391] = 12'h222;
rom[71392] = 12'h333;
rom[71393] = 12'h333;
rom[71394] = 12'h333;
rom[71395] = 12'h333;
rom[71396] = 12'h222;
rom[71397] = 12'h111;
rom[71398] = 12'h111;
rom[71399] = 12'h111;
rom[71400] = 12'h222;
rom[71401] = 12'h222;
rom[71402] = 12'h333;
rom[71403] = 12'h222;
rom[71404] = 12'h222;
rom[71405] = 12'h111;
rom[71406] = 12'h111;
rom[71407] = 12'h111;
rom[71408] = 12'h111;
rom[71409] = 12'h111;
rom[71410] = 12'h222;
rom[71411] = 12'h222;
rom[71412] = 12'h222;
rom[71413] = 12'h111;
rom[71414] = 12'h111;
rom[71415] = 12'h111;
rom[71416] = 12'h  0;
rom[71417] = 12'h  0;
rom[71418] = 12'h  0;
rom[71419] = 12'h  0;
rom[71420] = 12'h  0;
rom[71421] = 12'h  0;
rom[71422] = 12'h  0;
rom[71423] = 12'h  0;
rom[71424] = 12'h  0;
rom[71425] = 12'h  0;
rom[71426] = 12'h  0;
rom[71427] = 12'h  0;
rom[71428] = 12'h  0;
rom[71429] = 12'h  0;
rom[71430] = 12'h  0;
rom[71431] = 12'h  0;
rom[71432] = 12'h  0;
rom[71433] = 12'h  0;
rom[71434] = 12'h  0;
rom[71435] = 12'h  0;
rom[71436] = 12'h  0;
rom[71437] = 12'h  0;
rom[71438] = 12'h  0;
rom[71439] = 12'h  0;
rom[71440] = 12'h  0;
rom[71441] = 12'h  0;
rom[71442] = 12'h  0;
rom[71443] = 12'h  0;
rom[71444] = 12'h  0;
rom[71445] = 12'h  0;
rom[71446] = 12'h  0;
rom[71447] = 12'h  0;
rom[71448] = 12'h  0;
rom[71449] = 12'h  0;
rom[71450] = 12'h  0;
rom[71451] = 12'h  0;
rom[71452] = 12'h  0;
rom[71453] = 12'h  0;
rom[71454] = 12'h  0;
rom[71455] = 12'h  0;
rom[71456] = 12'h  0;
rom[71457] = 12'h  0;
rom[71458] = 12'h  0;
rom[71459] = 12'h  0;
rom[71460] = 12'h  0;
rom[71461] = 12'h  0;
rom[71462] = 12'h  0;
rom[71463] = 12'h  0;
rom[71464] = 12'h  0;
rom[71465] = 12'h  0;
rom[71466] = 12'h  0;
rom[71467] = 12'h  0;
rom[71468] = 12'h  0;
rom[71469] = 12'h  0;
rom[71470] = 12'h111;
rom[71471] = 12'h111;
rom[71472] = 12'h111;
rom[71473] = 12'h222;
rom[71474] = 12'h222;
rom[71475] = 12'h222;
rom[71476] = 12'h222;
rom[71477] = 12'h444;
rom[71478] = 12'h555;
rom[71479] = 12'h666;
rom[71480] = 12'h666;
rom[71481] = 12'h444;
rom[71482] = 12'h222;
rom[71483] = 12'h222;
rom[71484] = 12'h111;
rom[71485] = 12'h111;
rom[71486] = 12'h111;
rom[71487] = 12'h  0;
rom[71488] = 12'h  0;
rom[71489] = 12'h  0;
rom[71490] = 12'h  0;
rom[71491] = 12'h  0;
rom[71492] = 12'h  0;
rom[71493] = 12'h  0;
rom[71494] = 12'h  0;
rom[71495] = 12'h  0;
rom[71496] = 12'h111;
rom[71497] = 12'h111;
rom[71498] = 12'h111;
rom[71499] = 12'h111;
rom[71500] = 12'h222;
rom[71501] = 12'h222;
rom[71502] = 12'h333;
rom[71503] = 12'h333;
rom[71504] = 12'h333;
rom[71505] = 12'h444;
rom[71506] = 12'h444;
rom[71507] = 12'h555;
rom[71508] = 12'h555;
rom[71509] = 12'h555;
rom[71510] = 12'h666;
rom[71511] = 12'h666;
rom[71512] = 12'h777;
rom[71513] = 12'h777;
rom[71514] = 12'h777;
rom[71515] = 12'h888;
rom[71516] = 12'h999;
rom[71517] = 12'haaa;
rom[71518] = 12'hbbb;
rom[71519] = 12'hbbb;
rom[71520] = 12'hbbb;
rom[71521] = 12'hbbb;
rom[71522] = 12'hbbb;
rom[71523] = 12'hbbb;
rom[71524] = 12'hbbb;
rom[71525] = 12'hccc;
rom[71526] = 12'hccc;
rom[71527] = 12'hccc;
rom[71528] = 12'hddd;
rom[71529] = 12'hddd;
rom[71530] = 12'heee;
rom[71531] = 12'hfff;
rom[71532] = 12'hfff;
rom[71533] = 12'hfff;
rom[71534] = 12'hfff;
rom[71535] = 12'hfff;
rom[71536] = 12'hfff;
rom[71537] = 12'hfff;
rom[71538] = 12'hfff;
rom[71539] = 12'hfff;
rom[71540] = 12'hfff;
rom[71541] = 12'heee;
rom[71542] = 12'hddd;
rom[71543] = 12'hccc;
rom[71544] = 12'hbbb;
rom[71545] = 12'hbbb;
rom[71546] = 12'haaa;
rom[71547] = 12'haaa;
rom[71548] = 12'haaa;
rom[71549] = 12'h999;
rom[71550] = 12'h999;
rom[71551] = 12'h999;
rom[71552] = 12'h888;
rom[71553] = 12'h888;
rom[71554] = 12'h888;
rom[71555] = 12'h888;
rom[71556] = 12'h888;
rom[71557] = 12'h777;
rom[71558] = 12'h777;
rom[71559] = 12'h777;
rom[71560] = 12'h666;
rom[71561] = 12'h666;
rom[71562] = 12'h666;
rom[71563] = 12'h666;
rom[71564] = 12'h666;
rom[71565] = 12'h555;
rom[71566] = 12'h555;
rom[71567] = 12'h555;
rom[71568] = 12'h555;
rom[71569] = 12'h555;
rom[71570] = 12'h555;
rom[71571] = 12'h555;
rom[71572] = 12'h555;
rom[71573] = 12'h555;
rom[71574] = 12'h555;
rom[71575] = 12'h555;
rom[71576] = 12'h555;
rom[71577] = 12'h555;
rom[71578] = 12'h666;
rom[71579] = 12'h666;
rom[71580] = 12'h666;
rom[71581] = 12'h666;
rom[71582] = 12'h666;
rom[71583] = 12'h666;
rom[71584] = 12'h666;
rom[71585] = 12'h666;
rom[71586] = 12'h666;
rom[71587] = 12'h777;
rom[71588] = 12'h888;
rom[71589] = 12'h888;
rom[71590] = 12'h888;
rom[71591] = 12'h888;
rom[71592] = 12'h888;
rom[71593] = 12'h888;
rom[71594] = 12'h888;
rom[71595] = 12'h888;
rom[71596] = 12'h888;
rom[71597] = 12'h888;
rom[71598] = 12'h888;
rom[71599] = 12'h888;
rom[71600] = 12'hfff;
rom[71601] = 12'hfff;
rom[71602] = 12'hfff;
rom[71603] = 12'hfff;
rom[71604] = 12'hfff;
rom[71605] = 12'hfff;
rom[71606] = 12'hfff;
rom[71607] = 12'hfff;
rom[71608] = 12'hfff;
rom[71609] = 12'hfff;
rom[71610] = 12'hfff;
rom[71611] = 12'hfff;
rom[71612] = 12'hfff;
rom[71613] = 12'hfff;
rom[71614] = 12'hfff;
rom[71615] = 12'hfff;
rom[71616] = 12'hfff;
rom[71617] = 12'hfff;
rom[71618] = 12'hfff;
rom[71619] = 12'hfff;
rom[71620] = 12'hfff;
rom[71621] = 12'hfff;
rom[71622] = 12'hfff;
rom[71623] = 12'hfff;
rom[71624] = 12'hfff;
rom[71625] = 12'hfff;
rom[71626] = 12'hfff;
rom[71627] = 12'hfff;
rom[71628] = 12'hfff;
rom[71629] = 12'hfff;
rom[71630] = 12'hfff;
rom[71631] = 12'hfff;
rom[71632] = 12'hfff;
rom[71633] = 12'hfff;
rom[71634] = 12'hfff;
rom[71635] = 12'hfff;
rom[71636] = 12'hfff;
rom[71637] = 12'hfff;
rom[71638] = 12'hfff;
rom[71639] = 12'hfff;
rom[71640] = 12'hfff;
rom[71641] = 12'hfff;
rom[71642] = 12'hfff;
rom[71643] = 12'hfff;
rom[71644] = 12'hfff;
rom[71645] = 12'hfff;
rom[71646] = 12'hfff;
rom[71647] = 12'hfff;
rom[71648] = 12'hfff;
rom[71649] = 12'hfff;
rom[71650] = 12'hfff;
rom[71651] = 12'hfff;
rom[71652] = 12'hfff;
rom[71653] = 12'hfff;
rom[71654] = 12'hfff;
rom[71655] = 12'hfff;
rom[71656] = 12'hfff;
rom[71657] = 12'hfff;
rom[71658] = 12'hfff;
rom[71659] = 12'hfff;
rom[71660] = 12'hfff;
rom[71661] = 12'hfff;
rom[71662] = 12'hfff;
rom[71663] = 12'hfff;
rom[71664] = 12'hfff;
rom[71665] = 12'hfff;
rom[71666] = 12'hfff;
rom[71667] = 12'hfff;
rom[71668] = 12'hfff;
rom[71669] = 12'hfff;
rom[71670] = 12'hfff;
rom[71671] = 12'hfff;
rom[71672] = 12'hfff;
rom[71673] = 12'hfff;
rom[71674] = 12'hfff;
rom[71675] = 12'hfff;
rom[71676] = 12'hfff;
rom[71677] = 12'hfff;
rom[71678] = 12'hfff;
rom[71679] = 12'hfff;
rom[71680] = 12'hfff;
rom[71681] = 12'hfff;
rom[71682] = 12'hfff;
rom[71683] = 12'hfff;
rom[71684] = 12'hfff;
rom[71685] = 12'hfff;
rom[71686] = 12'hfff;
rom[71687] = 12'hfff;
rom[71688] = 12'hfff;
rom[71689] = 12'hfff;
rom[71690] = 12'hfff;
rom[71691] = 12'hfff;
rom[71692] = 12'hfff;
rom[71693] = 12'hfff;
rom[71694] = 12'hfff;
rom[71695] = 12'hfff;
rom[71696] = 12'hfff;
rom[71697] = 12'hfff;
rom[71698] = 12'hfff;
rom[71699] = 12'hfff;
rom[71700] = 12'hfff;
rom[71701] = 12'hfff;
rom[71702] = 12'hfff;
rom[71703] = 12'hfff;
rom[71704] = 12'hfff;
rom[71705] = 12'hfff;
rom[71706] = 12'hfff;
rom[71707] = 12'hfff;
rom[71708] = 12'hfff;
rom[71709] = 12'hfff;
rom[71710] = 12'heee;
rom[71711] = 12'hddd;
rom[71712] = 12'hddd;
rom[71713] = 12'hccc;
rom[71714] = 12'hccc;
rom[71715] = 12'hbbb;
rom[71716] = 12'haaa;
rom[71717] = 12'haaa;
rom[71718] = 12'haaa;
rom[71719] = 12'h999;
rom[71720] = 12'h999;
rom[71721] = 12'h999;
rom[71722] = 12'h888;
rom[71723] = 12'h888;
rom[71724] = 12'h888;
rom[71725] = 12'h888;
rom[71726] = 12'h888;
rom[71727] = 12'h777;
rom[71728] = 12'h777;
rom[71729] = 12'h777;
rom[71730] = 12'h777;
rom[71731] = 12'h777;
rom[71732] = 12'h777;
rom[71733] = 12'h666;
rom[71734] = 12'h666;
rom[71735] = 12'h666;
rom[71736] = 12'h666;
rom[71737] = 12'h666;
rom[71738] = 12'h555;
rom[71739] = 12'h555;
rom[71740] = 12'h555;
rom[71741] = 12'h444;
rom[71742] = 12'h444;
rom[71743] = 12'h444;
rom[71744] = 12'h444;
rom[71745] = 12'h444;
rom[71746] = 12'h444;
rom[71747] = 12'h444;
rom[71748] = 12'h444;
rom[71749] = 12'h444;
rom[71750] = 12'h444;
rom[71751] = 12'h444;
rom[71752] = 12'h444;
rom[71753] = 12'h444;
rom[71754] = 12'h444;
rom[71755] = 12'h444;
rom[71756] = 12'h555;
rom[71757] = 12'h555;
rom[71758] = 12'h555;
rom[71759] = 12'h555;
rom[71760] = 12'h555;
rom[71761] = 12'h555;
rom[71762] = 12'h444;
rom[71763] = 12'h444;
rom[71764] = 12'h444;
rom[71765] = 12'h444;
rom[71766] = 12'h555;
rom[71767] = 12'h555;
rom[71768] = 12'h555;
rom[71769] = 12'h555;
rom[71770] = 12'h555;
rom[71771] = 12'h555;
rom[71772] = 12'h555;
rom[71773] = 12'h555;
rom[71774] = 12'h555;
rom[71775] = 12'h555;
rom[71776] = 12'h555;
rom[71777] = 12'h444;
rom[71778] = 12'h444;
rom[71779] = 12'h444;
rom[71780] = 12'h444;
rom[71781] = 12'h333;
rom[71782] = 12'h333;
rom[71783] = 12'h333;
rom[71784] = 12'h333;
rom[71785] = 12'h333;
rom[71786] = 12'h333;
rom[71787] = 12'h333;
rom[71788] = 12'h333;
rom[71789] = 12'h333;
rom[71790] = 12'h222;
rom[71791] = 12'h222;
rom[71792] = 12'h333;
rom[71793] = 12'h333;
rom[71794] = 12'h333;
rom[71795] = 12'h333;
rom[71796] = 12'h333;
rom[71797] = 12'h222;
rom[71798] = 12'h111;
rom[71799] = 12'h111;
rom[71800] = 12'h222;
rom[71801] = 12'h222;
rom[71802] = 12'h333;
rom[71803] = 12'h222;
rom[71804] = 12'h222;
rom[71805] = 12'h111;
rom[71806] = 12'h111;
rom[71807] = 12'h111;
rom[71808] = 12'h111;
rom[71809] = 12'h222;
rom[71810] = 12'h222;
rom[71811] = 12'h333;
rom[71812] = 12'h222;
rom[71813] = 12'h111;
rom[71814] = 12'h111;
rom[71815] = 12'h  0;
rom[71816] = 12'h  0;
rom[71817] = 12'h  0;
rom[71818] = 12'h  0;
rom[71819] = 12'h  0;
rom[71820] = 12'h  0;
rom[71821] = 12'h  0;
rom[71822] = 12'h  0;
rom[71823] = 12'h  0;
rom[71824] = 12'h  0;
rom[71825] = 12'h  0;
rom[71826] = 12'h  0;
rom[71827] = 12'h  0;
rom[71828] = 12'h  0;
rom[71829] = 12'h  0;
rom[71830] = 12'h  0;
rom[71831] = 12'h111;
rom[71832] = 12'h  0;
rom[71833] = 12'h  0;
rom[71834] = 12'h  0;
rom[71835] = 12'h  0;
rom[71836] = 12'h  0;
rom[71837] = 12'h  0;
rom[71838] = 12'h  0;
rom[71839] = 12'h  0;
rom[71840] = 12'h  0;
rom[71841] = 12'h  0;
rom[71842] = 12'h  0;
rom[71843] = 12'h  0;
rom[71844] = 12'h  0;
rom[71845] = 12'h  0;
rom[71846] = 12'h  0;
rom[71847] = 12'h  0;
rom[71848] = 12'h  0;
rom[71849] = 12'h  0;
rom[71850] = 12'h  0;
rom[71851] = 12'h  0;
rom[71852] = 12'h  0;
rom[71853] = 12'h  0;
rom[71854] = 12'h  0;
rom[71855] = 12'h  0;
rom[71856] = 12'h  0;
rom[71857] = 12'h  0;
rom[71858] = 12'h  0;
rom[71859] = 12'h  0;
rom[71860] = 12'h  0;
rom[71861] = 12'h  0;
rom[71862] = 12'h  0;
rom[71863] = 12'h  0;
rom[71864] = 12'h  0;
rom[71865] = 12'h  0;
rom[71866] = 12'h  0;
rom[71867] = 12'h  0;
rom[71868] = 12'h  0;
rom[71869] = 12'h  0;
rom[71870] = 12'h111;
rom[71871] = 12'h111;
rom[71872] = 12'h111;
rom[71873] = 12'h111;
rom[71874] = 12'h222;
rom[71875] = 12'h222;
rom[71876] = 12'h222;
rom[71877] = 12'h444;
rom[71878] = 12'h555;
rom[71879] = 12'h666;
rom[71880] = 12'h666;
rom[71881] = 12'h444;
rom[71882] = 12'h222;
rom[71883] = 12'h222;
rom[71884] = 12'h111;
rom[71885] = 12'h111;
rom[71886] = 12'h111;
rom[71887] = 12'h  0;
rom[71888] = 12'h  0;
rom[71889] = 12'h  0;
rom[71890] = 12'h  0;
rom[71891] = 12'h  0;
rom[71892] = 12'h  0;
rom[71893] = 12'h  0;
rom[71894] = 12'h  0;
rom[71895] = 12'h  0;
rom[71896] = 12'h111;
rom[71897] = 12'h111;
rom[71898] = 12'h111;
rom[71899] = 12'h111;
rom[71900] = 12'h222;
rom[71901] = 12'h222;
rom[71902] = 12'h333;
rom[71903] = 12'h333;
rom[71904] = 12'h333;
rom[71905] = 12'h444;
rom[71906] = 12'h444;
rom[71907] = 12'h555;
rom[71908] = 12'h555;
rom[71909] = 12'h555;
rom[71910] = 12'h666;
rom[71911] = 12'h666;
rom[71912] = 12'h777;
rom[71913] = 12'h777;
rom[71914] = 12'h888;
rom[71915] = 12'h888;
rom[71916] = 12'haaa;
rom[71917] = 12'haaa;
rom[71918] = 12'hbbb;
rom[71919] = 12'hbbb;
rom[71920] = 12'hbbb;
rom[71921] = 12'hbbb;
rom[71922] = 12'hbbb;
rom[71923] = 12'hbbb;
rom[71924] = 12'hccc;
rom[71925] = 12'hccc;
rom[71926] = 12'hccc;
rom[71927] = 12'hddd;
rom[71928] = 12'hddd;
rom[71929] = 12'heee;
rom[71930] = 12'heee;
rom[71931] = 12'hfff;
rom[71932] = 12'hfff;
rom[71933] = 12'hfff;
rom[71934] = 12'hfff;
rom[71935] = 12'hfff;
rom[71936] = 12'hfff;
rom[71937] = 12'hfff;
rom[71938] = 12'hfff;
rom[71939] = 12'hfff;
rom[71940] = 12'heee;
rom[71941] = 12'hddd;
rom[71942] = 12'hccc;
rom[71943] = 12'hbbb;
rom[71944] = 12'hbbb;
rom[71945] = 12'haaa;
rom[71946] = 12'haaa;
rom[71947] = 12'haaa;
rom[71948] = 12'h999;
rom[71949] = 12'h999;
rom[71950] = 12'h999;
rom[71951] = 12'h888;
rom[71952] = 12'h888;
rom[71953] = 12'h888;
rom[71954] = 12'h888;
rom[71955] = 12'h777;
rom[71956] = 12'h777;
rom[71957] = 12'h777;
rom[71958] = 12'h777;
rom[71959] = 12'h777;
rom[71960] = 12'h666;
rom[71961] = 12'h666;
rom[71962] = 12'h666;
rom[71963] = 12'h666;
rom[71964] = 12'h555;
rom[71965] = 12'h555;
rom[71966] = 12'h555;
rom[71967] = 12'h555;
rom[71968] = 12'h555;
rom[71969] = 12'h555;
rom[71970] = 12'h555;
rom[71971] = 12'h555;
rom[71972] = 12'h555;
rom[71973] = 12'h555;
rom[71974] = 12'h555;
rom[71975] = 12'h555;
rom[71976] = 12'h555;
rom[71977] = 12'h555;
rom[71978] = 12'h555;
rom[71979] = 12'h555;
rom[71980] = 12'h555;
rom[71981] = 12'h555;
rom[71982] = 12'h666;
rom[71983] = 12'h666;
rom[71984] = 12'h666;
rom[71985] = 12'h666;
rom[71986] = 12'h666;
rom[71987] = 12'h666;
rom[71988] = 12'h777;
rom[71989] = 12'h888;
rom[71990] = 12'h888;
rom[71991] = 12'h888;
rom[71992] = 12'h888;
rom[71993] = 12'h888;
rom[71994] = 12'h888;
rom[71995] = 12'h777;
rom[71996] = 12'h777;
rom[71997] = 12'h888;
rom[71998] = 12'h888;
rom[71999] = 12'h888;
rom[72000] = 12'hfff;
rom[72001] = 12'hfff;
rom[72002] = 12'hfff;
rom[72003] = 12'hfff;
rom[72004] = 12'hfff;
rom[72005] = 12'hfff;
rom[72006] = 12'hfff;
rom[72007] = 12'hfff;
rom[72008] = 12'hfff;
rom[72009] = 12'hfff;
rom[72010] = 12'hfff;
rom[72011] = 12'hfff;
rom[72012] = 12'hfff;
rom[72013] = 12'hfff;
rom[72014] = 12'hfff;
rom[72015] = 12'hfff;
rom[72016] = 12'hfff;
rom[72017] = 12'hfff;
rom[72018] = 12'hfff;
rom[72019] = 12'hfff;
rom[72020] = 12'hfff;
rom[72021] = 12'hfff;
rom[72022] = 12'hfff;
rom[72023] = 12'hfff;
rom[72024] = 12'hfff;
rom[72025] = 12'hfff;
rom[72026] = 12'hfff;
rom[72027] = 12'hfff;
rom[72028] = 12'hfff;
rom[72029] = 12'hfff;
rom[72030] = 12'hfff;
rom[72031] = 12'hfff;
rom[72032] = 12'hfff;
rom[72033] = 12'hfff;
rom[72034] = 12'hfff;
rom[72035] = 12'hfff;
rom[72036] = 12'hfff;
rom[72037] = 12'hfff;
rom[72038] = 12'hfff;
rom[72039] = 12'hfff;
rom[72040] = 12'hfff;
rom[72041] = 12'hfff;
rom[72042] = 12'hfff;
rom[72043] = 12'hfff;
rom[72044] = 12'hfff;
rom[72045] = 12'hfff;
rom[72046] = 12'hfff;
rom[72047] = 12'hfff;
rom[72048] = 12'hfff;
rom[72049] = 12'hfff;
rom[72050] = 12'hfff;
rom[72051] = 12'hfff;
rom[72052] = 12'hfff;
rom[72053] = 12'hfff;
rom[72054] = 12'hfff;
rom[72055] = 12'hfff;
rom[72056] = 12'hfff;
rom[72057] = 12'hfff;
rom[72058] = 12'hfff;
rom[72059] = 12'hfff;
rom[72060] = 12'hfff;
rom[72061] = 12'hfff;
rom[72062] = 12'hfff;
rom[72063] = 12'hfff;
rom[72064] = 12'hfff;
rom[72065] = 12'hfff;
rom[72066] = 12'hfff;
rom[72067] = 12'hfff;
rom[72068] = 12'hfff;
rom[72069] = 12'hfff;
rom[72070] = 12'hfff;
rom[72071] = 12'hfff;
rom[72072] = 12'hfff;
rom[72073] = 12'hfff;
rom[72074] = 12'hfff;
rom[72075] = 12'hfff;
rom[72076] = 12'hfff;
rom[72077] = 12'hfff;
rom[72078] = 12'hfff;
rom[72079] = 12'hfff;
rom[72080] = 12'hfff;
rom[72081] = 12'hfff;
rom[72082] = 12'hfff;
rom[72083] = 12'hfff;
rom[72084] = 12'hfff;
rom[72085] = 12'hfff;
rom[72086] = 12'hfff;
rom[72087] = 12'hfff;
rom[72088] = 12'hfff;
rom[72089] = 12'hfff;
rom[72090] = 12'hfff;
rom[72091] = 12'hfff;
rom[72092] = 12'hfff;
rom[72093] = 12'hfff;
rom[72094] = 12'hfff;
rom[72095] = 12'hfff;
rom[72096] = 12'hfff;
rom[72097] = 12'hfff;
rom[72098] = 12'hfff;
rom[72099] = 12'hfff;
rom[72100] = 12'hfff;
rom[72101] = 12'hfff;
rom[72102] = 12'hfff;
rom[72103] = 12'hfff;
rom[72104] = 12'hfff;
rom[72105] = 12'hfff;
rom[72106] = 12'hfff;
rom[72107] = 12'hfff;
rom[72108] = 12'hfff;
rom[72109] = 12'hfff;
rom[72110] = 12'heee;
rom[72111] = 12'hddd;
rom[72112] = 12'hccc;
rom[72113] = 12'hccc;
rom[72114] = 12'hbbb;
rom[72115] = 12'hbbb;
rom[72116] = 12'haaa;
rom[72117] = 12'haaa;
rom[72118] = 12'h999;
rom[72119] = 12'h999;
rom[72120] = 12'h999;
rom[72121] = 12'h999;
rom[72122] = 12'h888;
rom[72123] = 12'h888;
rom[72124] = 12'h888;
rom[72125] = 12'h888;
rom[72126] = 12'h777;
rom[72127] = 12'h777;
rom[72128] = 12'h777;
rom[72129] = 12'h777;
rom[72130] = 12'h777;
rom[72131] = 12'h666;
rom[72132] = 12'h666;
rom[72133] = 12'h666;
rom[72134] = 12'h666;
rom[72135] = 12'h666;
rom[72136] = 12'h666;
rom[72137] = 12'h666;
rom[72138] = 12'h555;
rom[72139] = 12'h555;
rom[72140] = 12'h555;
rom[72141] = 12'h444;
rom[72142] = 12'h444;
rom[72143] = 12'h444;
rom[72144] = 12'h444;
rom[72145] = 12'h444;
rom[72146] = 12'h444;
rom[72147] = 12'h444;
rom[72148] = 12'h444;
rom[72149] = 12'h444;
rom[72150] = 12'h444;
rom[72151] = 12'h444;
rom[72152] = 12'h444;
rom[72153] = 12'h444;
rom[72154] = 12'h444;
rom[72155] = 12'h444;
rom[72156] = 12'h555;
rom[72157] = 12'h555;
rom[72158] = 12'h555;
rom[72159] = 12'h555;
rom[72160] = 12'h555;
rom[72161] = 12'h444;
rom[72162] = 12'h444;
rom[72163] = 12'h444;
rom[72164] = 12'h444;
rom[72165] = 12'h444;
rom[72166] = 12'h555;
rom[72167] = 12'h555;
rom[72168] = 12'h444;
rom[72169] = 12'h444;
rom[72170] = 12'h555;
rom[72171] = 12'h555;
rom[72172] = 12'h555;
rom[72173] = 12'h555;
rom[72174] = 12'h555;
rom[72175] = 12'h555;
rom[72176] = 12'h555;
rom[72177] = 12'h555;
rom[72178] = 12'h444;
rom[72179] = 12'h444;
rom[72180] = 12'h444;
rom[72181] = 12'h444;
rom[72182] = 12'h333;
rom[72183] = 12'h333;
rom[72184] = 12'h333;
rom[72185] = 12'h333;
rom[72186] = 12'h333;
rom[72187] = 12'h333;
rom[72188] = 12'h333;
rom[72189] = 12'h333;
rom[72190] = 12'h333;
rom[72191] = 12'h222;
rom[72192] = 12'h222;
rom[72193] = 12'h333;
rom[72194] = 12'h333;
rom[72195] = 12'h444;
rom[72196] = 12'h333;
rom[72197] = 12'h222;
rom[72198] = 12'h111;
rom[72199] = 12'h111;
rom[72200] = 12'h222;
rom[72201] = 12'h333;
rom[72202] = 12'h333;
rom[72203] = 12'h222;
rom[72204] = 12'h111;
rom[72205] = 12'h111;
rom[72206] = 12'h111;
rom[72207] = 12'h111;
rom[72208] = 12'h111;
rom[72209] = 12'h222;
rom[72210] = 12'h333;
rom[72211] = 12'h333;
rom[72212] = 12'h222;
rom[72213] = 12'h111;
rom[72214] = 12'h  0;
rom[72215] = 12'h  0;
rom[72216] = 12'h  0;
rom[72217] = 12'h  0;
rom[72218] = 12'h  0;
rom[72219] = 12'h  0;
rom[72220] = 12'h  0;
rom[72221] = 12'h  0;
rom[72222] = 12'h  0;
rom[72223] = 12'h  0;
rom[72224] = 12'h  0;
rom[72225] = 12'h  0;
rom[72226] = 12'h  0;
rom[72227] = 12'h  0;
rom[72228] = 12'h  0;
rom[72229] = 12'h  0;
rom[72230] = 12'h  0;
rom[72231] = 12'h111;
rom[72232] = 12'h  0;
rom[72233] = 12'h  0;
rom[72234] = 12'h  0;
rom[72235] = 12'h  0;
rom[72236] = 12'h  0;
rom[72237] = 12'h  0;
rom[72238] = 12'h  0;
rom[72239] = 12'h  0;
rom[72240] = 12'h  0;
rom[72241] = 12'h  0;
rom[72242] = 12'h  0;
rom[72243] = 12'h  0;
rom[72244] = 12'h  0;
rom[72245] = 12'h  0;
rom[72246] = 12'h  0;
rom[72247] = 12'h  0;
rom[72248] = 12'h  0;
rom[72249] = 12'h  0;
rom[72250] = 12'h  0;
rom[72251] = 12'h  0;
rom[72252] = 12'h  0;
rom[72253] = 12'h  0;
rom[72254] = 12'h  0;
rom[72255] = 12'h  0;
rom[72256] = 12'h  0;
rom[72257] = 12'h  0;
rom[72258] = 12'h  0;
rom[72259] = 12'h  0;
rom[72260] = 12'h  0;
rom[72261] = 12'h  0;
rom[72262] = 12'h  0;
rom[72263] = 12'h  0;
rom[72264] = 12'h  0;
rom[72265] = 12'h  0;
rom[72266] = 12'h  0;
rom[72267] = 12'h  0;
rom[72268] = 12'h  0;
rom[72269] = 12'h  0;
rom[72270] = 12'h111;
rom[72271] = 12'h111;
rom[72272] = 12'h111;
rom[72273] = 12'h222;
rom[72274] = 12'h222;
rom[72275] = 12'h222;
rom[72276] = 12'h333;
rom[72277] = 12'h444;
rom[72278] = 12'h555;
rom[72279] = 12'h666;
rom[72280] = 12'h666;
rom[72281] = 12'h444;
rom[72282] = 12'h222;
rom[72283] = 12'h222;
rom[72284] = 12'h111;
rom[72285] = 12'h111;
rom[72286] = 12'h111;
rom[72287] = 12'h111;
rom[72288] = 12'h  0;
rom[72289] = 12'h  0;
rom[72290] = 12'h  0;
rom[72291] = 12'h  0;
rom[72292] = 12'h  0;
rom[72293] = 12'h  0;
rom[72294] = 12'h  0;
rom[72295] = 12'h  0;
rom[72296] = 12'h111;
rom[72297] = 12'h111;
rom[72298] = 12'h111;
rom[72299] = 12'h111;
rom[72300] = 12'h222;
rom[72301] = 12'h222;
rom[72302] = 12'h222;
rom[72303] = 12'h333;
rom[72304] = 12'h333;
rom[72305] = 12'h333;
rom[72306] = 12'h444;
rom[72307] = 12'h555;
rom[72308] = 12'h555;
rom[72309] = 12'h555;
rom[72310] = 12'h666;
rom[72311] = 12'h666;
rom[72312] = 12'h666;
rom[72313] = 12'h777;
rom[72314] = 12'h888;
rom[72315] = 12'h999;
rom[72316] = 12'haaa;
rom[72317] = 12'haaa;
rom[72318] = 12'hbbb;
rom[72319] = 12'hbbb;
rom[72320] = 12'hbbb;
rom[72321] = 12'hbbb;
rom[72322] = 12'hccc;
rom[72323] = 12'hccc;
rom[72324] = 12'hccc;
rom[72325] = 12'hccc;
rom[72326] = 12'hddd;
rom[72327] = 12'hddd;
rom[72328] = 12'heee;
rom[72329] = 12'heee;
rom[72330] = 12'hfff;
rom[72331] = 12'hfff;
rom[72332] = 12'hfff;
rom[72333] = 12'hfff;
rom[72334] = 12'hfff;
rom[72335] = 12'hfff;
rom[72336] = 12'hfff;
rom[72337] = 12'hfff;
rom[72338] = 12'hfff;
rom[72339] = 12'heee;
rom[72340] = 12'hddd;
rom[72341] = 12'hccc;
rom[72342] = 12'hccc;
rom[72343] = 12'hbbb;
rom[72344] = 12'haaa;
rom[72345] = 12'haaa;
rom[72346] = 12'haaa;
rom[72347] = 12'h999;
rom[72348] = 12'h999;
rom[72349] = 12'h999;
rom[72350] = 12'h888;
rom[72351] = 12'h888;
rom[72352] = 12'h888;
rom[72353] = 12'h777;
rom[72354] = 12'h777;
rom[72355] = 12'h777;
rom[72356] = 12'h777;
rom[72357] = 12'h777;
rom[72358] = 12'h777;
rom[72359] = 12'h777;
rom[72360] = 12'h666;
rom[72361] = 12'h666;
rom[72362] = 12'h666;
rom[72363] = 12'h666;
rom[72364] = 12'h555;
rom[72365] = 12'h555;
rom[72366] = 12'h555;
rom[72367] = 12'h555;
rom[72368] = 12'h555;
rom[72369] = 12'h555;
rom[72370] = 12'h555;
rom[72371] = 12'h555;
rom[72372] = 12'h555;
rom[72373] = 12'h555;
rom[72374] = 12'h555;
rom[72375] = 12'h555;
rom[72376] = 12'h555;
rom[72377] = 12'h555;
rom[72378] = 12'h555;
rom[72379] = 12'h555;
rom[72380] = 12'h555;
rom[72381] = 12'h555;
rom[72382] = 12'h555;
rom[72383] = 12'h555;
rom[72384] = 12'h666;
rom[72385] = 12'h555;
rom[72386] = 12'h555;
rom[72387] = 12'h555;
rom[72388] = 12'h666;
rom[72389] = 12'h777;
rom[72390] = 12'h777;
rom[72391] = 12'h777;
rom[72392] = 12'h777;
rom[72393] = 12'h777;
rom[72394] = 12'h777;
rom[72395] = 12'h777;
rom[72396] = 12'h777;
rom[72397] = 12'h777;
rom[72398] = 12'h777;
rom[72399] = 12'h777;
rom[72400] = 12'hfff;
rom[72401] = 12'hfff;
rom[72402] = 12'hfff;
rom[72403] = 12'hfff;
rom[72404] = 12'hfff;
rom[72405] = 12'hfff;
rom[72406] = 12'hfff;
rom[72407] = 12'hfff;
rom[72408] = 12'hfff;
rom[72409] = 12'hfff;
rom[72410] = 12'hfff;
rom[72411] = 12'hfff;
rom[72412] = 12'hfff;
rom[72413] = 12'hfff;
rom[72414] = 12'hfff;
rom[72415] = 12'hfff;
rom[72416] = 12'hfff;
rom[72417] = 12'hfff;
rom[72418] = 12'hfff;
rom[72419] = 12'hfff;
rom[72420] = 12'hfff;
rom[72421] = 12'hfff;
rom[72422] = 12'hfff;
rom[72423] = 12'hfff;
rom[72424] = 12'hfff;
rom[72425] = 12'hfff;
rom[72426] = 12'hfff;
rom[72427] = 12'hfff;
rom[72428] = 12'hfff;
rom[72429] = 12'hfff;
rom[72430] = 12'hfff;
rom[72431] = 12'hfff;
rom[72432] = 12'hfff;
rom[72433] = 12'hfff;
rom[72434] = 12'hfff;
rom[72435] = 12'hfff;
rom[72436] = 12'hfff;
rom[72437] = 12'hfff;
rom[72438] = 12'hfff;
rom[72439] = 12'hfff;
rom[72440] = 12'hfff;
rom[72441] = 12'hfff;
rom[72442] = 12'hfff;
rom[72443] = 12'hfff;
rom[72444] = 12'hfff;
rom[72445] = 12'hfff;
rom[72446] = 12'hfff;
rom[72447] = 12'hfff;
rom[72448] = 12'hfff;
rom[72449] = 12'hfff;
rom[72450] = 12'hfff;
rom[72451] = 12'hfff;
rom[72452] = 12'hfff;
rom[72453] = 12'hfff;
rom[72454] = 12'hfff;
rom[72455] = 12'hfff;
rom[72456] = 12'hfff;
rom[72457] = 12'hfff;
rom[72458] = 12'hfff;
rom[72459] = 12'hfff;
rom[72460] = 12'hfff;
rom[72461] = 12'hfff;
rom[72462] = 12'hfff;
rom[72463] = 12'hfff;
rom[72464] = 12'hfff;
rom[72465] = 12'hfff;
rom[72466] = 12'hfff;
rom[72467] = 12'hfff;
rom[72468] = 12'hfff;
rom[72469] = 12'hfff;
rom[72470] = 12'hfff;
rom[72471] = 12'hfff;
rom[72472] = 12'hfff;
rom[72473] = 12'hfff;
rom[72474] = 12'hfff;
rom[72475] = 12'hfff;
rom[72476] = 12'hfff;
rom[72477] = 12'hfff;
rom[72478] = 12'hfff;
rom[72479] = 12'hfff;
rom[72480] = 12'hfff;
rom[72481] = 12'hfff;
rom[72482] = 12'hfff;
rom[72483] = 12'hfff;
rom[72484] = 12'hfff;
rom[72485] = 12'hfff;
rom[72486] = 12'hfff;
rom[72487] = 12'hfff;
rom[72488] = 12'hfff;
rom[72489] = 12'hfff;
rom[72490] = 12'hfff;
rom[72491] = 12'hfff;
rom[72492] = 12'hfff;
rom[72493] = 12'hfff;
rom[72494] = 12'hfff;
rom[72495] = 12'hfff;
rom[72496] = 12'hfff;
rom[72497] = 12'hfff;
rom[72498] = 12'hfff;
rom[72499] = 12'hfff;
rom[72500] = 12'hfff;
rom[72501] = 12'hfff;
rom[72502] = 12'hfff;
rom[72503] = 12'hfff;
rom[72504] = 12'hfff;
rom[72505] = 12'hfff;
rom[72506] = 12'hfff;
rom[72507] = 12'hfff;
rom[72508] = 12'hfff;
rom[72509] = 12'hfff;
rom[72510] = 12'heee;
rom[72511] = 12'hddd;
rom[72512] = 12'hccc;
rom[72513] = 12'hccc;
rom[72514] = 12'hbbb;
rom[72515] = 12'hbbb;
rom[72516] = 12'haaa;
rom[72517] = 12'haaa;
rom[72518] = 12'haaa;
rom[72519] = 12'h999;
rom[72520] = 12'h999;
rom[72521] = 12'h999;
rom[72522] = 12'h888;
rom[72523] = 12'h888;
rom[72524] = 12'h888;
rom[72525] = 12'h777;
rom[72526] = 12'h777;
rom[72527] = 12'h777;
rom[72528] = 12'h777;
rom[72529] = 12'h777;
rom[72530] = 12'h777;
rom[72531] = 12'h777;
rom[72532] = 12'h777;
rom[72533] = 12'h777;
rom[72534] = 12'h666;
rom[72535] = 12'h666;
rom[72536] = 12'h666;
rom[72537] = 12'h666;
rom[72538] = 12'h555;
rom[72539] = 12'h555;
rom[72540] = 12'h555;
rom[72541] = 12'h555;
rom[72542] = 12'h444;
rom[72543] = 12'h444;
rom[72544] = 12'h444;
rom[72545] = 12'h444;
rom[72546] = 12'h444;
rom[72547] = 12'h444;
rom[72548] = 12'h444;
rom[72549] = 12'h444;
rom[72550] = 12'h444;
rom[72551] = 12'h444;
rom[72552] = 12'h444;
rom[72553] = 12'h444;
rom[72554] = 12'h444;
rom[72555] = 12'h444;
rom[72556] = 12'h555;
rom[72557] = 12'h555;
rom[72558] = 12'h555;
rom[72559] = 12'h555;
rom[72560] = 12'h555;
rom[72561] = 12'h555;
rom[72562] = 12'h555;
rom[72563] = 12'h444;
rom[72564] = 12'h444;
rom[72565] = 12'h444;
rom[72566] = 12'h444;
rom[72567] = 12'h444;
rom[72568] = 12'h444;
rom[72569] = 12'h444;
rom[72570] = 12'h444;
rom[72571] = 12'h444;
rom[72572] = 12'h444;
rom[72573] = 12'h555;
rom[72574] = 12'h555;
rom[72575] = 12'h555;
rom[72576] = 12'h555;
rom[72577] = 12'h555;
rom[72578] = 12'h555;
rom[72579] = 12'h555;
rom[72580] = 12'h444;
rom[72581] = 12'h444;
rom[72582] = 12'h444;
rom[72583] = 12'h444;
rom[72584] = 12'h333;
rom[72585] = 12'h333;
rom[72586] = 12'h333;
rom[72587] = 12'h333;
rom[72588] = 12'h333;
rom[72589] = 12'h333;
rom[72590] = 12'h333;
rom[72591] = 12'h333;
rom[72592] = 12'h333;
rom[72593] = 12'h333;
rom[72594] = 12'h333;
rom[72595] = 12'h444;
rom[72596] = 12'h333;
rom[72597] = 12'h333;
rom[72598] = 12'h222;
rom[72599] = 12'h222;
rom[72600] = 12'h222;
rom[72601] = 12'h333;
rom[72602] = 12'h333;
rom[72603] = 12'h222;
rom[72604] = 12'h111;
rom[72605] = 12'h111;
rom[72606] = 12'h111;
rom[72607] = 12'h111;
rom[72608] = 12'h222;
rom[72609] = 12'h222;
rom[72610] = 12'h333;
rom[72611] = 12'h222;
rom[72612] = 12'h222;
rom[72613] = 12'h111;
rom[72614] = 12'h  0;
rom[72615] = 12'h  0;
rom[72616] = 12'h  0;
rom[72617] = 12'h  0;
rom[72618] = 12'h  0;
rom[72619] = 12'h  0;
rom[72620] = 12'h  0;
rom[72621] = 12'h  0;
rom[72622] = 12'h  0;
rom[72623] = 12'h  0;
rom[72624] = 12'h  0;
rom[72625] = 12'h  0;
rom[72626] = 12'h  0;
rom[72627] = 12'h  0;
rom[72628] = 12'h  0;
rom[72629] = 12'h  0;
rom[72630] = 12'h111;
rom[72631] = 12'h111;
rom[72632] = 12'h111;
rom[72633] = 12'h  0;
rom[72634] = 12'h  0;
rom[72635] = 12'h  0;
rom[72636] = 12'h  0;
rom[72637] = 12'h  0;
rom[72638] = 12'h  0;
rom[72639] = 12'h  0;
rom[72640] = 12'h  0;
rom[72641] = 12'h  0;
rom[72642] = 12'h  0;
rom[72643] = 12'h  0;
rom[72644] = 12'h  0;
rom[72645] = 12'h  0;
rom[72646] = 12'h  0;
rom[72647] = 12'h  0;
rom[72648] = 12'h  0;
rom[72649] = 12'h  0;
rom[72650] = 12'h  0;
rom[72651] = 12'h  0;
rom[72652] = 12'h  0;
rom[72653] = 12'h  0;
rom[72654] = 12'h  0;
rom[72655] = 12'h  0;
rom[72656] = 12'h  0;
rom[72657] = 12'h  0;
rom[72658] = 12'h  0;
rom[72659] = 12'h  0;
rom[72660] = 12'h  0;
rom[72661] = 12'h  0;
rom[72662] = 12'h  0;
rom[72663] = 12'h  0;
rom[72664] = 12'h  0;
rom[72665] = 12'h  0;
rom[72666] = 12'h  0;
rom[72667] = 12'h  0;
rom[72668] = 12'h  0;
rom[72669] = 12'h  0;
rom[72670] = 12'h111;
rom[72671] = 12'h111;
rom[72672] = 12'h111;
rom[72673] = 12'h222;
rom[72674] = 12'h222;
rom[72675] = 12'h222;
rom[72676] = 12'h333;
rom[72677] = 12'h444;
rom[72678] = 12'h555;
rom[72679] = 12'h666;
rom[72680] = 12'h666;
rom[72681] = 12'h444;
rom[72682] = 12'h222;
rom[72683] = 12'h222;
rom[72684] = 12'h222;
rom[72685] = 12'h111;
rom[72686] = 12'h111;
rom[72687] = 12'h111;
rom[72688] = 12'h111;
rom[72689] = 12'h  0;
rom[72690] = 12'h  0;
rom[72691] = 12'h  0;
rom[72692] = 12'h  0;
rom[72693] = 12'h  0;
rom[72694] = 12'h111;
rom[72695] = 12'h111;
rom[72696] = 12'h111;
rom[72697] = 12'h111;
rom[72698] = 12'h111;
rom[72699] = 12'h222;
rom[72700] = 12'h222;
rom[72701] = 12'h222;
rom[72702] = 12'h222;
rom[72703] = 12'h333;
rom[72704] = 12'h333;
rom[72705] = 12'h333;
rom[72706] = 12'h444;
rom[72707] = 12'h555;
rom[72708] = 12'h555;
rom[72709] = 12'h555;
rom[72710] = 12'h666;
rom[72711] = 12'h666;
rom[72712] = 12'h666;
rom[72713] = 12'h777;
rom[72714] = 12'h888;
rom[72715] = 12'h999;
rom[72716] = 12'haaa;
rom[72717] = 12'hbbb;
rom[72718] = 12'hbbb;
rom[72719] = 12'hbbb;
rom[72720] = 12'hbbb;
rom[72721] = 12'hccc;
rom[72722] = 12'hccc;
rom[72723] = 12'hccc;
rom[72724] = 12'hccc;
rom[72725] = 12'hddd;
rom[72726] = 12'hddd;
rom[72727] = 12'heee;
rom[72728] = 12'heee;
rom[72729] = 12'hfff;
rom[72730] = 12'hfff;
rom[72731] = 12'hfff;
rom[72732] = 12'hfff;
rom[72733] = 12'hfff;
rom[72734] = 12'hfff;
rom[72735] = 12'hfff;
rom[72736] = 12'hfff;
rom[72737] = 12'hfff;
rom[72738] = 12'heee;
rom[72739] = 12'hddd;
rom[72740] = 12'hccc;
rom[72741] = 12'hccc;
rom[72742] = 12'hbbb;
rom[72743] = 12'hbbb;
rom[72744] = 12'haaa;
rom[72745] = 12'h999;
rom[72746] = 12'h999;
rom[72747] = 12'h999;
rom[72748] = 12'h999;
rom[72749] = 12'h888;
rom[72750] = 12'h888;
rom[72751] = 12'h888;
rom[72752] = 12'h777;
rom[72753] = 12'h777;
rom[72754] = 12'h777;
rom[72755] = 12'h777;
rom[72756] = 12'h777;
rom[72757] = 12'h777;
rom[72758] = 12'h666;
rom[72759] = 12'h666;
rom[72760] = 12'h666;
rom[72761] = 12'h666;
rom[72762] = 12'h666;
rom[72763] = 12'h666;
rom[72764] = 12'h555;
rom[72765] = 12'h555;
rom[72766] = 12'h555;
rom[72767] = 12'h555;
rom[72768] = 12'h555;
rom[72769] = 12'h555;
rom[72770] = 12'h555;
rom[72771] = 12'h555;
rom[72772] = 12'h555;
rom[72773] = 12'h555;
rom[72774] = 12'h555;
rom[72775] = 12'h555;
rom[72776] = 12'h555;
rom[72777] = 12'h555;
rom[72778] = 12'h555;
rom[72779] = 12'h555;
rom[72780] = 12'h555;
rom[72781] = 12'h555;
rom[72782] = 12'h555;
rom[72783] = 12'h555;
rom[72784] = 12'h666;
rom[72785] = 12'h555;
rom[72786] = 12'h555;
rom[72787] = 12'h555;
rom[72788] = 12'h555;
rom[72789] = 12'h666;
rom[72790] = 12'h777;
rom[72791] = 12'h777;
rom[72792] = 12'h777;
rom[72793] = 12'h777;
rom[72794] = 12'h777;
rom[72795] = 12'h777;
rom[72796] = 12'h777;
rom[72797] = 12'h777;
rom[72798] = 12'h777;
rom[72799] = 12'h777;
rom[72800] = 12'hfff;
rom[72801] = 12'hfff;
rom[72802] = 12'hfff;
rom[72803] = 12'hfff;
rom[72804] = 12'hfff;
rom[72805] = 12'hfff;
rom[72806] = 12'hfff;
rom[72807] = 12'hfff;
rom[72808] = 12'hfff;
rom[72809] = 12'hfff;
rom[72810] = 12'hfff;
rom[72811] = 12'hfff;
rom[72812] = 12'hfff;
rom[72813] = 12'hfff;
rom[72814] = 12'hfff;
rom[72815] = 12'hfff;
rom[72816] = 12'hfff;
rom[72817] = 12'hfff;
rom[72818] = 12'hfff;
rom[72819] = 12'hfff;
rom[72820] = 12'hfff;
rom[72821] = 12'hfff;
rom[72822] = 12'hfff;
rom[72823] = 12'hfff;
rom[72824] = 12'hfff;
rom[72825] = 12'hfff;
rom[72826] = 12'hfff;
rom[72827] = 12'hfff;
rom[72828] = 12'hfff;
rom[72829] = 12'hfff;
rom[72830] = 12'hfff;
rom[72831] = 12'hfff;
rom[72832] = 12'hfff;
rom[72833] = 12'hfff;
rom[72834] = 12'hfff;
rom[72835] = 12'hfff;
rom[72836] = 12'hfff;
rom[72837] = 12'hfff;
rom[72838] = 12'hfff;
rom[72839] = 12'hfff;
rom[72840] = 12'hfff;
rom[72841] = 12'hfff;
rom[72842] = 12'hfff;
rom[72843] = 12'hfff;
rom[72844] = 12'hfff;
rom[72845] = 12'hfff;
rom[72846] = 12'hfff;
rom[72847] = 12'hfff;
rom[72848] = 12'hfff;
rom[72849] = 12'hfff;
rom[72850] = 12'hfff;
rom[72851] = 12'hfff;
rom[72852] = 12'hfff;
rom[72853] = 12'hfff;
rom[72854] = 12'hfff;
rom[72855] = 12'hfff;
rom[72856] = 12'hfff;
rom[72857] = 12'hfff;
rom[72858] = 12'hfff;
rom[72859] = 12'hfff;
rom[72860] = 12'hfff;
rom[72861] = 12'hfff;
rom[72862] = 12'hfff;
rom[72863] = 12'hfff;
rom[72864] = 12'hfff;
rom[72865] = 12'hfff;
rom[72866] = 12'hfff;
rom[72867] = 12'hfff;
rom[72868] = 12'hfff;
rom[72869] = 12'hfff;
rom[72870] = 12'hfff;
rom[72871] = 12'hfff;
rom[72872] = 12'hfff;
rom[72873] = 12'hfff;
rom[72874] = 12'hfff;
rom[72875] = 12'hfff;
rom[72876] = 12'hfff;
rom[72877] = 12'hfff;
rom[72878] = 12'hfff;
rom[72879] = 12'hfff;
rom[72880] = 12'hfff;
rom[72881] = 12'hfff;
rom[72882] = 12'hfff;
rom[72883] = 12'hfff;
rom[72884] = 12'hfff;
rom[72885] = 12'hfff;
rom[72886] = 12'hfff;
rom[72887] = 12'hfff;
rom[72888] = 12'hfff;
rom[72889] = 12'hfff;
rom[72890] = 12'hfff;
rom[72891] = 12'hfff;
rom[72892] = 12'hfff;
rom[72893] = 12'hfff;
rom[72894] = 12'hfff;
rom[72895] = 12'hfff;
rom[72896] = 12'hfff;
rom[72897] = 12'hfff;
rom[72898] = 12'hfff;
rom[72899] = 12'hfff;
rom[72900] = 12'hfff;
rom[72901] = 12'hfff;
rom[72902] = 12'hfff;
rom[72903] = 12'hfff;
rom[72904] = 12'hfff;
rom[72905] = 12'hfff;
rom[72906] = 12'hfff;
rom[72907] = 12'hfff;
rom[72908] = 12'hfff;
rom[72909] = 12'hfff;
rom[72910] = 12'heee;
rom[72911] = 12'heee;
rom[72912] = 12'hddd;
rom[72913] = 12'hddd;
rom[72914] = 12'hccc;
rom[72915] = 12'hbbb;
rom[72916] = 12'haaa;
rom[72917] = 12'haaa;
rom[72918] = 12'haaa;
rom[72919] = 12'h999;
rom[72920] = 12'h999;
rom[72921] = 12'h888;
rom[72922] = 12'h888;
rom[72923] = 12'h888;
rom[72924] = 12'h888;
rom[72925] = 12'h888;
rom[72926] = 12'h777;
rom[72927] = 12'h777;
rom[72928] = 12'h777;
rom[72929] = 12'h777;
rom[72930] = 12'h777;
rom[72931] = 12'h777;
rom[72932] = 12'h777;
rom[72933] = 12'h777;
rom[72934] = 12'h777;
rom[72935] = 12'h777;
rom[72936] = 12'h666;
rom[72937] = 12'h666;
rom[72938] = 12'h666;
rom[72939] = 12'h555;
rom[72940] = 12'h555;
rom[72941] = 12'h555;
rom[72942] = 12'h555;
rom[72943] = 12'h555;
rom[72944] = 12'h444;
rom[72945] = 12'h444;
rom[72946] = 12'h444;
rom[72947] = 12'h444;
rom[72948] = 12'h444;
rom[72949] = 12'h444;
rom[72950] = 12'h444;
rom[72951] = 12'h444;
rom[72952] = 12'h444;
rom[72953] = 12'h444;
rom[72954] = 12'h444;
rom[72955] = 12'h555;
rom[72956] = 12'h555;
rom[72957] = 12'h555;
rom[72958] = 12'h555;
rom[72959] = 12'h555;
rom[72960] = 12'h555;
rom[72961] = 12'h555;
rom[72962] = 12'h555;
rom[72963] = 12'h555;
rom[72964] = 12'h555;
rom[72965] = 12'h444;
rom[72966] = 12'h444;
rom[72967] = 12'h444;
rom[72968] = 12'h444;
rom[72969] = 12'h444;
rom[72970] = 12'h444;
rom[72971] = 12'h444;
rom[72972] = 12'h555;
rom[72973] = 12'h555;
rom[72974] = 12'h555;
rom[72975] = 12'h555;
rom[72976] = 12'h555;
rom[72977] = 12'h555;
rom[72978] = 12'h555;
rom[72979] = 12'h555;
rom[72980] = 12'h555;
rom[72981] = 12'h555;
rom[72982] = 12'h555;
rom[72983] = 12'h444;
rom[72984] = 12'h444;
rom[72985] = 12'h444;
rom[72986] = 12'h333;
rom[72987] = 12'h333;
rom[72988] = 12'h333;
rom[72989] = 12'h333;
rom[72990] = 12'h333;
rom[72991] = 12'h333;
rom[72992] = 12'h333;
rom[72993] = 12'h333;
rom[72994] = 12'h333;
rom[72995] = 12'h444;
rom[72996] = 12'h444;
rom[72997] = 12'h333;
rom[72998] = 12'h333;
rom[72999] = 12'h222;
rom[73000] = 12'h333;
rom[73001] = 12'h333;
rom[73002] = 12'h333;
rom[73003] = 12'h222;
rom[73004] = 12'h222;
rom[73005] = 12'h222;
rom[73006] = 12'h111;
rom[73007] = 12'h111;
rom[73008] = 12'h222;
rom[73009] = 12'h222;
rom[73010] = 12'h222;
rom[73011] = 12'h222;
rom[73012] = 12'h111;
rom[73013] = 12'h111;
rom[73014] = 12'h111;
rom[73015] = 12'h111;
rom[73016] = 12'h111;
rom[73017] = 12'h  0;
rom[73018] = 12'h  0;
rom[73019] = 12'h  0;
rom[73020] = 12'h  0;
rom[73021] = 12'h111;
rom[73022] = 12'h  0;
rom[73023] = 12'h  0;
rom[73024] = 12'h  0;
rom[73025] = 12'h  0;
rom[73026] = 12'h  0;
rom[73027] = 12'h  0;
rom[73028] = 12'h  0;
rom[73029] = 12'h111;
rom[73030] = 12'h111;
rom[73031] = 12'h111;
rom[73032] = 12'h111;
rom[73033] = 12'h111;
rom[73034] = 12'h  0;
rom[73035] = 12'h  0;
rom[73036] = 12'h  0;
rom[73037] = 12'h  0;
rom[73038] = 12'h  0;
rom[73039] = 12'h  0;
rom[73040] = 12'h  0;
rom[73041] = 12'h  0;
rom[73042] = 12'h  0;
rom[73043] = 12'h  0;
rom[73044] = 12'h  0;
rom[73045] = 12'h  0;
rom[73046] = 12'h  0;
rom[73047] = 12'h  0;
rom[73048] = 12'h  0;
rom[73049] = 12'h  0;
rom[73050] = 12'h  0;
rom[73051] = 12'h  0;
rom[73052] = 12'h  0;
rom[73053] = 12'h  0;
rom[73054] = 12'h  0;
rom[73055] = 12'h  0;
rom[73056] = 12'h  0;
rom[73057] = 12'h  0;
rom[73058] = 12'h  0;
rom[73059] = 12'h  0;
rom[73060] = 12'h  0;
rom[73061] = 12'h  0;
rom[73062] = 12'h  0;
rom[73063] = 12'h  0;
rom[73064] = 12'h  0;
rom[73065] = 12'h  0;
rom[73066] = 12'h  0;
rom[73067] = 12'h  0;
rom[73068] = 12'h  0;
rom[73069] = 12'h  0;
rom[73070] = 12'h111;
rom[73071] = 12'h111;
rom[73072] = 12'h111;
rom[73073] = 12'h222;
rom[73074] = 12'h222;
rom[73075] = 12'h222;
rom[73076] = 12'h333;
rom[73077] = 12'h444;
rom[73078] = 12'h555;
rom[73079] = 12'h666;
rom[73080] = 12'h666;
rom[73081] = 12'h444;
rom[73082] = 12'h222;
rom[73083] = 12'h222;
rom[73084] = 12'h222;
rom[73085] = 12'h111;
rom[73086] = 12'h111;
rom[73087] = 12'h111;
rom[73088] = 12'h111;
rom[73089] = 12'h111;
rom[73090] = 12'h111;
rom[73091] = 12'h  0;
rom[73092] = 12'h  0;
rom[73093] = 12'h111;
rom[73094] = 12'h111;
rom[73095] = 12'h111;
rom[73096] = 12'h111;
rom[73097] = 12'h111;
rom[73098] = 12'h111;
rom[73099] = 12'h222;
rom[73100] = 12'h222;
rom[73101] = 12'h222;
rom[73102] = 12'h333;
rom[73103] = 12'h333;
rom[73104] = 12'h333;
rom[73105] = 12'h444;
rom[73106] = 12'h444;
rom[73107] = 12'h555;
rom[73108] = 12'h555;
rom[73109] = 12'h666;
rom[73110] = 12'h666;
rom[73111] = 12'h777;
rom[73112] = 12'h777;
rom[73113] = 12'h777;
rom[73114] = 12'h888;
rom[73115] = 12'h999;
rom[73116] = 12'haaa;
rom[73117] = 12'hbbb;
rom[73118] = 12'hbbb;
rom[73119] = 12'hbbb;
rom[73120] = 12'hccc;
rom[73121] = 12'hccc;
rom[73122] = 12'hccc;
rom[73123] = 12'hccc;
rom[73124] = 12'hddd;
rom[73125] = 12'hddd;
rom[73126] = 12'heee;
rom[73127] = 12'hfff;
rom[73128] = 12'hfff;
rom[73129] = 12'hfff;
rom[73130] = 12'hfff;
rom[73131] = 12'hfff;
rom[73132] = 12'hfff;
rom[73133] = 12'hfff;
rom[73134] = 12'hfff;
rom[73135] = 12'hfff;
rom[73136] = 12'hfff;
rom[73137] = 12'heee;
rom[73138] = 12'hddd;
rom[73139] = 12'hccc;
rom[73140] = 12'hbbb;
rom[73141] = 12'hbbb;
rom[73142] = 12'hbbb;
rom[73143] = 12'haaa;
rom[73144] = 12'haaa;
rom[73145] = 12'h999;
rom[73146] = 12'h999;
rom[73147] = 12'h888;
rom[73148] = 12'h888;
rom[73149] = 12'h888;
rom[73150] = 12'h888;
rom[73151] = 12'h777;
rom[73152] = 12'h777;
rom[73153] = 12'h777;
rom[73154] = 12'h777;
rom[73155] = 12'h777;
rom[73156] = 12'h777;
rom[73157] = 12'h666;
rom[73158] = 12'h666;
rom[73159] = 12'h666;
rom[73160] = 12'h666;
rom[73161] = 12'h666;
rom[73162] = 12'h666;
rom[73163] = 12'h555;
rom[73164] = 12'h555;
rom[73165] = 12'h555;
rom[73166] = 12'h555;
rom[73167] = 12'h555;
rom[73168] = 12'h555;
rom[73169] = 12'h555;
rom[73170] = 12'h555;
rom[73171] = 12'h555;
rom[73172] = 12'h555;
rom[73173] = 12'h555;
rom[73174] = 12'h555;
rom[73175] = 12'h555;
rom[73176] = 12'h555;
rom[73177] = 12'h555;
rom[73178] = 12'h555;
rom[73179] = 12'h555;
rom[73180] = 12'h555;
rom[73181] = 12'h555;
rom[73182] = 12'h555;
rom[73183] = 12'h555;
rom[73184] = 12'h555;
rom[73185] = 12'h555;
rom[73186] = 12'h555;
rom[73187] = 12'h555;
rom[73188] = 12'h555;
rom[73189] = 12'h666;
rom[73190] = 12'h666;
rom[73191] = 12'h777;
rom[73192] = 12'h777;
rom[73193] = 12'h777;
rom[73194] = 12'h777;
rom[73195] = 12'h777;
rom[73196] = 12'h777;
rom[73197] = 12'h777;
rom[73198] = 12'h666;
rom[73199] = 12'h666;
rom[73200] = 12'hfff;
rom[73201] = 12'hfff;
rom[73202] = 12'hfff;
rom[73203] = 12'hfff;
rom[73204] = 12'hfff;
rom[73205] = 12'hfff;
rom[73206] = 12'hfff;
rom[73207] = 12'hfff;
rom[73208] = 12'hfff;
rom[73209] = 12'hfff;
rom[73210] = 12'hfff;
rom[73211] = 12'hfff;
rom[73212] = 12'hfff;
rom[73213] = 12'hfff;
rom[73214] = 12'hfff;
rom[73215] = 12'hfff;
rom[73216] = 12'hfff;
rom[73217] = 12'hfff;
rom[73218] = 12'hfff;
rom[73219] = 12'hfff;
rom[73220] = 12'hfff;
rom[73221] = 12'hfff;
rom[73222] = 12'hfff;
rom[73223] = 12'hfff;
rom[73224] = 12'hfff;
rom[73225] = 12'hfff;
rom[73226] = 12'hfff;
rom[73227] = 12'hfff;
rom[73228] = 12'hfff;
rom[73229] = 12'hfff;
rom[73230] = 12'hfff;
rom[73231] = 12'hfff;
rom[73232] = 12'hfff;
rom[73233] = 12'hfff;
rom[73234] = 12'hfff;
rom[73235] = 12'hfff;
rom[73236] = 12'hfff;
rom[73237] = 12'hfff;
rom[73238] = 12'hfff;
rom[73239] = 12'hfff;
rom[73240] = 12'hfff;
rom[73241] = 12'hfff;
rom[73242] = 12'hfff;
rom[73243] = 12'hfff;
rom[73244] = 12'hfff;
rom[73245] = 12'hfff;
rom[73246] = 12'hfff;
rom[73247] = 12'hfff;
rom[73248] = 12'hfff;
rom[73249] = 12'hfff;
rom[73250] = 12'hfff;
rom[73251] = 12'hfff;
rom[73252] = 12'hfff;
rom[73253] = 12'hfff;
rom[73254] = 12'hfff;
rom[73255] = 12'hfff;
rom[73256] = 12'hfff;
rom[73257] = 12'hfff;
rom[73258] = 12'hfff;
rom[73259] = 12'hfff;
rom[73260] = 12'hfff;
rom[73261] = 12'hfff;
rom[73262] = 12'hfff;
rom[73263] = 12'hfff;
rom[73264] = 12'hfff;
rom[73265] = 12'hfff;
rom[73266] = 12'hfff;
rom[73267] = 12'hfff;
rom[73268] = 12'hfff;
rom[73269] = 12'hfff;
rom[73270] = 12'hfff;
rom[73271] = 12'hfff;
rom[73272] = 12'hfff;
rom[73273] = 12'hfff;
rom[73274] = 12'hfff;
rom[73275] = 12'hfff;
rom[73276] = 12'hfff;
rom[73277] = 12'hfff;
rom[73278] = 12'hfff;
rom[73279] = 12'hfff;
rom[73280] = 12'hfff;
rom[73281] = 12'hfff;
rom[73282] = 12'hfff;
rom[73283] = 12'hfff;
rom[73284] = 12'hfff;
rom[73285] = 12'hfff;
rom[73286] = 12'hfff;
rom[73287] = 12'hfff;
rom[73288] = 12'hfff;
rom[73289] = 12'hfff;
rom[73290] = 12'hfff;
rom[73291] = 12'hfff;
rom[73292] = 12'hfff;
rom[73293] = 12'hfff;
rom[73294] = 12'hfff;
rom[73295] = 12'hfff;
rom[73296] = 12'hfff;
rom[73297] = 12'hfff;
rom[73298] = 12'hfff;
rom[73299] = 12'hfff;
rom[73300] = 12'hfff;
rom[73301] = 12'hfff;
rom[73302] = 12'hfff;
rom[73303] = 12'hfff;
rom[73304] = 12'hfff;
rom[73305] = 12'hfff;
rom[73306] = 12'hfff;
rom[73307] = 12'hfff;
rom[73308] = 12'hfff;
rom[73309] = 12'hfff;
rom[73310] = 12'hfff;
rom[73311] = 12'hfff;
rom[73312] = 12'heee;
rom[73313] = 12'heee;
rom[73314] = 12'hddd;
rom[73315] = 12'hccc;
rom[73316] = 12'hbbb;
rom[73317] = 12'haaa;
rom[73318] = 12'h999;
rom[73319] = 12'h999;
rom[73320] = 12'h888;
rom[73321] = 12'h888;
rom[73322] = 12'h888;
rom[73323] = 12'h888;
rom[73324] = 12'h888;
rom[73325] = 12'h888;
rom[73326] = 12'h888;
rom[73327] = 12'h888;
rom[73328] = 12'h777;
rom[73329] = 12'h777;
rom[73330] = 12'h777;
rom[73331] = 12'h777;
rom[73332] = 12'h777;
rom[73333] = 12'h777;
rom[73334] = 12'h777;
rom[73335] = 12'h777;
rom[73336] = 12'h777;
rom[73337] = 12'h666;
rom[73338] = 12'h666;
rom[73339] = 12'h666;
rom[73340] = 12'h666;
rom[73341] = 12'h666;
rom[73342] = 12'h666;
rom[73343] = 12'h555;
rom[73344] = 12'h555;
rom[73345] = 12'h555;
rom[73346] = 12'h555;
rom[73347] = 12'h555;
rom[73348] = 12'h444;
rom[73349] = 12'h444;
rom[73350] = 12'h444;
rom[73351] = 12'h444;
rom[73352] = 12'h444;
rom[73353] = 12'h444;
rom[73354] = 12'h444;
rom[73355] = 12'h555;
rom[73356] = 12'h555;
rom[73357] = 12'h555;
rom[73358] = 12'h555;
rom[73359] = 12'h555;
rom[73360] = 12'h444;
rom[73361] = 12'h555;
rom[73362] = 12'h555;
rom[73363] = 12'h555;
rom[73364] = 12'h555;
rom[73365] = 12'h555;
rom[73366] = 12'h555;
rom[73367] = 12'h444;
rom[73368] = 12'h555;
rom[73369] = 12'h555;
rom[73370] = 12'h555;
rom[73371] = 12'h555;
rom[73372] = 12'h555;
rom[73373] = 12'h555;
rom[73374] = 12'h555;
rom[73375] = 12'h444;
rom[73376] = 12'h555;
rom[73377] = 12'h555;
rom[73378] = 12'h555;
rom[73379] = 12'h555;
rom[73380] = 12'h555;
rom[73381] = 12'h555;
rom[73382] = 12'h555;
rom[73383] = 12'h555;
rom[73384] = 12'h555;
rom[73385] = 12'h444;
rom[73386] = 12'h444;
rom[73387] = 12'h333;
rom[73388] = 12'h333;
rom[73389] = 12'h333;
rom[73390] = 12'h333;
rom[73391] = 12'h333;
rom[73392] = 12'h333;
rom[73393] = 12'h333;
rom[73394] = 12'h333;
rom[73395] = 12'h444;
rom[73396] = 12'h444;
rom[73397] = 12'h444;
rom[73398] = 12'h333;
rom[73399] = 12'h333;
rom[73400] = 12'h333;
rom[73401] = 12'h333;
rom[73402] = 12'h333;
rom[73403] = 12'h222;
rom[73404] = 12'h222;
rom[73405] = 12'h222;
rom[73406] = 12'h222;
rom[73407] = 12'h111;
rom[73408] = 12'h333;
rom[73409] = 12'h333;
rom[73410] = 12'h222;
rom[73411] = 12'h222;
rom[73412] = 12'h111;
rom[73413] = 12'h111;
rom[73414] = 12'h111;
rom[73415] = 12'h111;
rom[73416] = 12'h111;
rom[73417] = 12'h111;
rom[73418] = 12'h  0;
rom[73419] = 12'h  0;
rom[73420] = 12'h111;
rom[73421] = 12'h111;
rom[73422] = 12'h  0;
rom[73423] = 12'h  0;
rom[73424] = 12'h  0;
rom[73425] = 12'h  0;
rom[73426] = 12'h  0;
rom[73427] = 12'h  0;
rom[73428] = 12'h  0;
rom[73429] = 12'h111;
rom[73430] = 12'h111;
rom[73431] = 12'h111;
rom[73432] = 12'h111;
rom[73433] = 12'h111;
rom[73434] = 12'h  0;
rom[73435] = 12'h  0;
rom[73436] = 12'h  0;
rom[73437] = 12'h  0;
rom[73438] = 12'h  0;
rom[73439] = 12'h  0;
rom[73440] = 12'h  0;
rom[73441] = 12'h  0;
rom[73442] = 12'h  0;
rom[73443] = 12'h  0;
rom[73444] = 12'h  0;
rom[73445] = 12'h  0;
rom[73446] = 12'h  0;
rom[73447] = 12'h  0;
rom[73448] = 12'h  0;
rom[73449] = 12'h  0;
rom[73450] = 12'h  0;
rom[73451] = 12'h  0;
rom[73452] = 12'h  0;
rom[73453] = 12'h  0;
rom[73454] = 12'h  0;
rom[73455] = 12'h  0;
rom[73456] = 12'h  0;
rom[73457] = 12'h  0;
rom[73458] = 12'h  0;
rom[73459] = 12'h  0;
rom[73460] = 12'h  0;
rom[73461] = 12'h  0;
rom[73462] = 12'h  0;
rom[73463] = 12'h  0;
rom[73464] = 12'h  0;
rom[73465] = 12'h  0;
rom[73466] = 12'h  0;
rom[73467] = 12'h  0;
rom[73468] = 12'h  0;
rom[73469] = 12'h  0;
rom[73470] = 12'h111;
rom[73471] = 12'h111;
rom[73472] = 12'h111;
rom[73473] = 12'h222;
rom[73474] = 12'h222;
rom[73475] = 12'h222;
rom[73476] = 12'h333;
rom[73477] = 12'h444;
rom[73478] = 12'h555;
rom[73479] = 12'h777;
rom[73480] = 12'h666;
rom[73481] = 12'h444;
rom[73482] = 12'h222;
rom[73483] = 12'h222;
rom[73484] = 12'h222;
rom[73485] = 12'h222;
rom[73486] = 12'h111;
rom[73487] = 12'h111;
rom[73488] = 12'h111;
rom[73489] = 12'h111;
rom[73490] = 12'h111;
rom[73491] = 12'h111;
rom[73492] = 12'h111;
rom[73493] = 12'h111;
rom[73494] = 12'h111;
rom[73495] = 12'h111;
rom[73496] = 12'h111;
rom[73497] = 12'h111;
rom[73498] = 12'h222;
rom[73499] = 12'h222;
rom[73500] = 12'h222;
rom[73501] = 12'h222;
rom[73502] = 12'h333;
rom[73503] = 12'h333;
rom[73504] = 12'h333;
rom[73505] = 12'h444;
rom[73506] = 12'h444;
rom[73507] = 12'h555;
rom[73508] = 12'h555;
rom[73509] = 12'h666;
rom[73510] = 12'h666;
rom[73511] = 12'h777;
rom[73512] = 12'h777;
rom[73513] = 12'h777;
rom[73514] = 12'h888;
rom[73515] = 12'h999;
rom[73516] = 12'haaa;
rom[73517] = 12'hbbb;
rom[73518] = 12'hbbb;
rom[73519] = 12'hbbb;
rom[73520] = 12'hccc;
rom[73521] = 12'hccc;
rom[73522] = 12'hccc;
rom[73523] = 12'hccc;
rom[73524] = 12'hddd;
rom[73525] = 12'heee;
rom[73526] = 12'hfff;
rom[73527] = 12'hfff;
rom[73528] = 12'hfff;
rom[73529] = 12'hfff;
rom[73530] = 12'hfff;
rom[73531] = 12'hfff;
rom[73532] = 12'hfff;
rom[73533] = 12'hfff;
rom[73534] = 12'hfff;
rom[73535] = 12'hfff;
rom[73536] = 12'heee;
rom[73537] = 12'heee;
rom[73538] = 12'hddd;
rom[73539] = 12'hccc;
rom[73540] = 12'hbbb;
rom[73541] = 12'hbbb;
rom[73542] = 12'haaa;
rom[73543] = 12'haaa;
rom[73544] = 12'haaa;
rom[73545] = 12'h999;
rom[73546] = 12'h999;
rom[73547] = 12'h888;
rom[73548] = 12'h888;
rom[73549] = 12'h888;
rom[73550] = 12'h777;
rom[73551] = 12'h777;
rom[73552] = 12'h777;
rom[73553] = 12'h777;
rom[73554] = 12'h777;
rom[73555] = 12'h777;
rom[73556] = 12'h666;
rom[73557] = 12'h666;
rom[73558] = 12'h666;
rom[73559] = 12'h666;
rom[73560] = 12'h666;
rom[73561] = 12'h666;
rom[73562] = 12'h555;
rom[73563] = 12'h555;
rom[73564] = 12'h555;
rom[73565] = 12'h555;
rom[73566] = 12'h555;
rom[73567] = 12'h555;
rom[73568] = 12'h555;
rom[73569] = 12'h444;
rom[73570] = 12'h444;
rom[73571] = 12'h444;
rom[73572] = 12'h444;
rom[73573] = 12'h444;
rom[73574] = 12'h444;
rom[73575] = 12'h444;
rom[73576] = 12'h555;
rom[73577] = 12'h555;
rom[73578] = 12'h555;
rom[73579] = 12'h555;
rom[73580] = 12'h555;
rom[73581] = 12'h555;
rom[73582] = 12'h555;
rom[73583] = 12'h555;
rom[73584] = 12'h444;
rom[73585] = 12'h555;
rom[73586] = 12'h555;
rom[73587] = 12'h555;
rom[73588] = 12'h555;
rom[73589] = 12'h555;
rom[73590] = 12'h666;
rom[73591] = 12'h666;
rom[73592] = 12'h666;
rom[73593] = 12'h666;
rom[73594] = 12'h666;
rom[73595] = 12'h666;
rom[73596] = 12'h666;
rom[73597] = 12'h666;
rom[73598] = 12'h666;
rom[73599] = 12'h666;
rom[73600] = 12'hfff;
rom[73601] = 12'hfff;
rom[73602] = 12'hfff;
rom[73603] = 12'hfff;
rom[73604] = 12'hfff;
rom[73605] = 12'hfff;
rom[73606] = 12'hfff;
rom[73607] = 12'hfff;
rom[73608] = 12'hfff;
rom[73609] = 12'hfff;
rom[73610] = 12'hfff;
rom[73611] = 12'hfff;
rom[73612] = 12'hfff;
rom[73613] = 12'hfff;
rom[73614] = 12'hfff;
rom[73615] = 12'hfff;
rom[73616] = 12'hfff;
rom[73617] = 12'hfff;
rom[73618] = 12'hfff;
rom[73619] = 12'hfff;
rom[73620] = 12'hfff;
rom[73621] = 12'hfff;
rom[73622] = 12'hfff;
rom[73623] = 12'hfff;
rom[73624] = 12'hfff;
rom[73625] = 12'hfff;
rom[73626] = 12'hfff;
rom[73627] = 12'hfff;
rom[73628] = 12'hfff;
rom[73629] = 12'hfff;
rom[73630] = 12'hfff;
rom[73631] = 12'hfff;
rom[73632] = 12'hfff;
rom[73633] = 12'hfff;
rom[73634] = 12'hfff;
rom[73635] = 12'hfff;
rom[73636] = 12'hfff;
rom[73637] = 12'hfff;
rom[73638] = 12'hfff;
rom[73639] = 12'hfff;
rom[73640] = 12'hfff;
rom[73641] = 12'hfff;
rom[73642] = 12'hfff;
rom[73643] = 12'hfff;
rom[73644] = 12'hfff;
rom[73645] = 12'hfff;
rom[73646] = 12'hfff;
rom[73647] = 12'hfff;
rom[73648] = 12'hfff;
rom[73649] = 12'hfff;
rom[73650] = 12'hfff;
rom[73651] = 12'hfff;
rom[73652] = 12'hfff;
rom[73653] = 12'hfff;
rom[73654] = 12'hfff;
rom[73655] = 12'hfff;
rom[73656] = 12'hfff;
rom[73657] = 12'hfff;
rom[73658] = 12'hfff;
rom[73659] = 12'hfff;
rom[73660] = 12'hfff;
rom[73661] = 12'hfff;
rom[73662] = 12'hfff;
rom[73663] = 12'hfff;
rom[73664] = 12'hfff;
rom[73665] = 12'hfff;
rom[73666] = 12'hfff;
rom[73667] = 12'hfff;
rom[73668] = 12'hfff;
rom[73669] = 12'hfff;
rom[73670] = 12'hfff;
rom[73671] = 12'hfff;
rom[73672] = 12'hfff;
rom[73673] = 12'hfff;
rom[73674] = 12'hfff;
rom[73675] = 12'hfff;
rom[73676] = 12'hfff;
rom[73677] = 12'hfff;
rom[73678] = 12'hfff;
rom[73679] = 12'hfff;
rom[73680] = 12'hfff;
rom[73681] = 12'hfff;
rom[73682] = 12'hfff;
rom[73683] = 12'hfff;
rom[73684] = 12'hfff;
rom[73685] = 12'hfff;
rom[73686] = 12'hfff;
rom[73687] = 12'hfff;
rom[73688] = 12'hfff;
rom[73689] = 12'hfff;
rom[73690] = 12'hfff;
rom[73691] = 12'hfff;
rom[73692] = 12'hfff;
rom[73693] = 12'hfff;
rom[73694] = 12'hfff;
rom[73695] = 12'hfff;
rom[73696] = 12'hfff;
rom[73697] = 12'hfff;
rom[73698] = 12'hfff;
rom[73699] = 12'hfff;
rom[73700] = 12'hfff;
rom[73701] = 12'hfff;
rom[73702] = 12'hfff;
rom[73703] = 12'hfff;
rom[73704] = 12'hfff;
rom[73705] = 12'hfff;
rom[73706] = 12'hfff;
rom[73707] = 12'hfff;
rom[73708] = 12'hfff;
rom[73709] = 12'hfff;
rom[73710] = 12'hfff;
rom[73711] = 12'hfff;
rom[73712] = 12'hfff;
rom[73713] = 12'heee;
rom[73714] = 12'heee;
rom[73715] = 12'hddd;
rom[73716] = 12'hddd;
rom[73717] = 12'hccc;
rom[73718] = 12'hbbb;
rom[73719] = 12'haaa;
rom[73720] = 12'h999;
rom[73721] = 12'h999;
rom[73722] = 12'h888;
rom[73723] = 12'h888;
rom[73724] = 12'h888;
rom[73725] = 12'h888;
rom[73726] = 12'h888;
rom[73727] = 12'h777;
rom[73728] = 12'h777;
rom[73729] = 12'h777;
rom[73730] = 12'h777;
rom[73731] = 12'h777;
rom[73732] = 12'h777;
rom[73733] = 12'h777;
rom[73734] = 12'h777;
rom[73735] = 12'h777;
rom[73736] = 12'h777;
rom[73737] = 12'h777;
rom[73738] = 12'h777;
rom[73739] = 12'h666;
rom[73740] = 12'h666;
rom[73741] = 12'h666;
rom[73742] = 12'h666;
rom[73743] = 12'h666;
rom[73744] = 12'h666;
rom[73745] = 12'h555;
rom[73746] = 12'h555;
rom[73747] = 12'h555;
rom[73748] = 12'h444;
rom[73749] = 12'h444;
rom[73750] = 12'h444;
rom[73751] = 12'h444;
rom[73752] = 12'h555;
rom[73753] = 12'h555;
rom[73754] = 12'h555;
rom[73755] = 12'h555;
rom[73756] = 12'h555;
rom[73757] = 12'h555;
rom[73758] = 12'h555;
rom[73759] = 12'h555;
rom[73760] = 12'h555;
rom[73761] = 12'h555;
rom[73762] = 12'h555;
rom[73763] = 12'h555;
rom[73764] = 12'h555;
rom[73765] = 12'h555;
rom[73766] = 12'h555;
rom[73767] = 12'h555;
rom[73768] = 12'h555;
rom[73769] = 12'h555;
rom[73770] = 12'h555;
rom[73771] = 12'h555;
rom[73772] = 12'h555;
rom[73773] = 12'h555;
rom[73774] = 12'h444;
rom[73775] = 12'h444;
rom[73776] = 12'h555;
rom[73777] = 12'h555;
rom[73778] = 12'h555;
rom[73779] = 12'h555;
rom[73780] = 12'h555;
rom[73781] = 12'h555;
rom[73782] = 12'h555;
rom[73783] = 12'h666;
rom[73784] = 12'h666;
rom[73785] = 12'h555;
rom[73786] = 12'h555;
rom[73787] = 12'h444;
rom[73788] = 12'h444;
rom[73789] = 12'h444;
rom[73790] = 12'h444;
rom[73791] = 12'h444;
rom[73792] = 12'h333;
rom[73793] = 12'h333;
rom[73794] = 12'h333;
rom[73795] = 12'h333;
rom[73796] = 12'h444;
rom[73797] = 12'h555;
rom[73798] = 12'h444;
rom[73799] = 12'h333;
rom[73800] = 12'h333;
rom[73801] = 12'h333;
rom[73802] = 12'h333;
rom[73803] = 12'h222;
rom[73804] = 12'h222;
rom[73805] = 12'h222;
rom[73806] = 12'h222;
rom[73807] = 12'h222;
rom[73808] = 12'h333;
rom[73809] = 12'h333;
rom[73810] = 12'h222;
rom[73811] = 12'h111;
rom[73812] = 12'h111;
rom[73813] = 12'h111;
rom[73814] = 12'h111;
rom[73815] = 12'h111;
rom[73816] = 12'h111;
rom[73817] = 12'h111;
rom[73818] = 12'h111;
rom[73819] = 12'h  0;
rom[73820] = 12'h  0;
rom[73821] = 12'h  0;
rom[73822] = 12'h111;
rom[73823] = 12'h111;
rom[73824] = 12'h111;
rom[73825] = 12'h111;
rom[73826] = 12'h  0;
rom[73827] = 12'h111;
rom[73828] = 12'h111;
rom[73829] = 12'h111;
rom[73830] = 12'h111;
rom[73831] = 12'h111;
rom[73832] = 12'h111;
rom[73833] = 12'h  0;
rom[73834] = 12'h  0;
rom[73835] = 12'h  0;
rom[73836] = 12'h  0;
rom[73837] = 12'h  0;
rom[73838] = 12'h  0;
rom[73839] = 12'h  0;
rom[73840] = 12'h  0;
rom[73841] = 12'h  0;
rom[73842] = 12'h  0;
rom[73843] = 12'h  0;
rom[73844] = 12'h  0;
rom[73845] = 12'h  0;
rom[73846] = 12'h  0;
rom[73847] = 12'h  0;
rom[73848] = 12'h  0;
rom[73849] = 12'h  0;
rom[73850] = 12'h  0;
rom[73851] = 12'h  0;
rom[73852] = 12'h  0;
rom[73853] = 12'h  0;
rom[73854] = 12'h  0;
rom[73855] = 12'h  0;
rom[73856] = 12'h  0;
rom[73857] = 12'h  0;
rom[73858] = 12'h  0;
rom[73859] = 12'h  0;
rom[73860] = 12'h  0;
rom[73861] = 12'h  0;
rom[73862] = 12'h  0;
rom[73863] = 12'h  0;
rom[73864] = 12'h  0;
rom[73865] = 12'h  0;
rom[73866] = 12'h  0;
rom[73867] = 12'h  0;
rom[73868] = 12'h  0;
rom[73869] = 12'h  0;
rom[73870] = 12'h  0;
rom[73871] = 12'h111;
rom[73872] = 12'h111;
rom[73873] = 12'h111;
rom[73874] = 12'h222;
rom[73875] = 12'h333;
rom[73876] = 12'h333;
rom[73877] = 12'h444;
rom[73878] = 12'h555;
rom[73879] = 12'h777;
rom[73880] = 12'h666;
rom[73881] = 12'h555;
rom[73882] = 12'h333;
rom[73883] = 12'h222;
rom[73884] = 12'h222;
rom[73885] = 12'h111;
rom[73886] = 12'h111;
rom[73887] = 12'h111;
rom[73888] = 12'h111;
rom[73889] = 12'h111;
rom[73890] = 12'h111;
rom[73891] = 12'h111;
rom[73892] = 12'h111;
rom[73893] = 12'h111;
rom[73894] = 12'h111;
rom[73895] = 12'h111;
rom[73896] = 12'h111;
rom[73897] = 12'h111;
rom[73898] = 12'h222;
rom[73899] = 12'h222;
rom[73900] = 12'h222;
rom[73901] = 12'h333;
rom[73902] = 12'h333;
rom[73903] = 12'h333;
rom[73904] = 12'h444;
rom[73905] = 12'h444;
rom[73906] = 12'h555;
rom[73907] = 12'h555;
rom[73908] = 12'h555;
rom[73909] = 12'h666;
rom[73910] = 12'h666;
rom[73911] = 12'h777;
rom[73912] = 12'h777;
rom[73913] = 12'h777;
rom[73914] = 12'h888;
rom[73915] = 12'haaa;
rom[73916] = 12'hbbb;
rom[73917] = 12'hbbb;
rom[73918] = 12'hbbb;
rom[73919] = 12'hccc;
rom[73920] = 12'hccc;
rom[73921] = 12'hccc;
rom[73922] = 12'hccc;
rom[73923] = 12'hddd;
rom[73924] = 12'heee;
rom[73925] = 12'hfff;
rom[73926] = 12'hfff;
rom[73927] = 12'hfff;
rom[73928] = 12'hfff;
rom[73929] = 12'hfff;
rom[73930] = 12'hfff;
rom[73931] = 12'hfff;
rom[73932] = 12'hfff;
rom[73933] = 12'hfff;
rom[73934] = 12'hfff;
rom[73935] = 12'heee;
rom[73936] = 12'hddd;
rom[73937] = 12'hccc;
rom[73938] = 12'hccc;
rom[73939] = 12'hbbb;
rom[73940] = 12'haaa;
rom[73941] = 12'haaa;
rom[73942] = 12'haaa;
rom[73943] = 12'h999;
rom[73944] = 12'haaa;
rom[73945] = 12'h999;
rom[73946] = 12'h999;
rom[73947] = 12'h999;
rom[73948] = 12'h888;
rom[73949] = 12'h888;
rom[73950] = 12'h777;
rom[73951] = 12'h666;
rom[73952] = 12'h777;
rom[73953] = 12'h666;
rom[73954] = 12'h666;
rom[73955] = 12'h666;
rom[73956] = 12'h666;
rom[73957] = 12'h666;
rom[73958] = 12'h666;
rom[73959] = 12'h666;
rom[73960] = 12'h555;
rom[73961] = 12'h555;
rom[73962] = 12'h555;
rom[73963] = 12'h555;
rom[73964] = 12'h555;
rom[73965] = 12'h555;
rom[73966] = 12'h555;
rom[73967] = 12'h444;
rom[73968] = 12'h444;
rom[73969] = 12'h444;
rom[73970] = 12'h444;
rom[73971] = 12'h444;
rom[73972] = 12'h444;
rom[73973] = 12'h444;
rom[73974] = 12'h444;
rom[73975] = 12'h444;
rom[73976] = 12'h444;
rom[73977] = 12'h444;
rom[73978] = 12'h444;
rom[73979] = 12'h444;
rom[73980] = 12'h444;
rom[73981] = 12'h444;
rom[73982] = 12'h444;
rom[73983] = 12'h444;
rom[73984] = 12'h444;
rom[73985] = 12'h444;
rom[73986] = 12'h444;
rom[73987] = 12'h555;
rom[73988] = 12'h555;
rom[73989] = 12'h555;
rom[73990] = 12'h555;
rom[73991] = 12'h555;
rom[73992] = 12'h666;
rom[73993] = 12'h666;
rom[73994] = 12'h666;
rom[73995] = 12'h666;
rom[73996] = 12'h555;
rom[73997] = 12'h666;
rom[73998] = 12'h666;
rom[73999] = 12'h666;
rom[74000] = 12'hfff;
rom[74001] = 12'hfff;
rom[74002] = 12'hfff;
rom[74003] = 12'hfff;
rom[74004] = 12'hfff;
rom[74005] = 12'hfff;
rom[74006] = 12'hfff;
rom[74007] = 12'hfff;
rom[74008] = 12'hfff;
rom[74009] = 12'hfff;
rom[74010] = 12'hfff;
rom[74011] = 12'hfff;
rom[74012] = 12'hfff;
rom[74013] = 12'hfff;
rom[74014] = 12'hfff;
rom[74015] = 12'hfff;
rom[74016] = 12'hfff;
rom[74017] = 12'hfff;
rom[74018] = 12'hfff;
rom[74019] = 12'hfff;
rom[74020] = 12'hfff;
rom[74021] = 12'hfff;
rom[74022] = 12'hfff;
rom[74023] = 12'hfff;
rom[74024] = 12'hfff;
rom[74025] = 12'hfff;
rom[74026] = 12'hfff;
rom[74027] = 12'hfff;
rom[74028] = 12'hfff;
rom[74029] = 12'hfff;
rom[74030] = 12'hfff;
rom[74031] = 12'hfff;
rom[74032] = 12'hfff;
rom[74033] = 12'hfff;
rom[74034] = 12'hfff;
rom[74035] = 12'hfff;
rom[74036] = 12'hfff;
rom[74037] = 12'hfff;
rom[74038] = 12'hfff;
rom[74039] = 12'hfff;
rom[74040] = 12'hfff;
rom[74041] = 12'hfff;
rom[74042] = 12'hfff;
rom[74043] = 12'hfff;
rom[74044] = 12'hfff;
rom[74045] = 12'hfff;
rom[74046] = 12'hfff;
rom[74047] = 12'hfff;
rom[74048] = 12'hfff;
rom[74049] = 12'hfff;
rom[74050] = 12'hfff;
rom[74051] = 12'hfff;
rom[74052] = 12'hfff;
rom[74053] = 12'hfff;
rom[74054] = 12'hfff;
rom[74055] = 12'hfff;
rom[74056] = 12'hfff;
rom[74057] = 12'hfff;
rom[74058] = 12'hfff;
rom[74059] = 12'hfff;
rom[74060] = 12'hfff;
rom[74061] = 12'hfff;
rom[74062] = 12'hfff;
rom[74063] = 12'hfff;
rom[74064] = 12'hfff;
rom[74065] = 12'hfff;
rom[74066] = 12'hfff;
rom[74067] = 12'hfff;
rom[74068] = 12'hfff;
rom[74069] = 12'hfff;
rom[74070] = 12'hfff;
rom[74071] = 12'hfff;
rom[74072] = 12'hfff;
rom[74073] = 12'hfff;
rom[74074] = 12'hfff;
rom[74075] = 12'hfff;
rom[74076] = 12'hfff;
rom[74077] = 12'hfff;
rom[74078] = 12'hfff;
rom[74079] = 12'hfff;
rom[74080] = 12'hfff;
rom[74081] = 12'hfff;
rom[74082] = 12'hfff;
rom[74083] = 12'hfff;
rom[74084] = 12'hfff;
rom[74085] = 12'hfff;
rom[74086] = 12'hfff;
rom[74087] = 12'hfff;
rom[74088] = 12'hfff;
rom[74089] = 12'hfff;
rom[74090] = 12'hfff;
rom[74091] = 12'hfff;
rom[74092] = 12'hfff;
rom[74093] = 12'hfff;
rom[74094] = 12'hfff;
rom[74095] = 12'hfff;
rom[74096] = 12'hfff;
rom[74097] = 12'hfff;
rom[74098] = 12'hfff;
rom[74099] = 12'hfff;
rom[74100] = 12'hfff;
rom[74101] = 12'hfff;
rom[74102] = 12'hfff;
rom[74103] = 12'hfff;
rom[74104] = 12'hfff;
rom[74105] = 12'hfff;
rom[74106] = 12'hfff;
rom[74107] = 12'hfff;
rom[74108] = 12'hfff;
rom[74109] = 12'hfff;
rom[74110] = 12'hfff;
rom[74111] = 12'hfff;
rom[74112] = 12'heee;
rom[74113] = 12'heee;
rom[74114] = 12'heee;
rom[74115] = 12'heee;
rom[74116] = 12'heee;
rom[74117] = 12'hddd;
rom[74118] = 12'hccc;
rom[74119] = 12'hccc;
rom[74120] = 12'hbbb;
rom[74121] = 12'haaa;
rom[74122] = 12'haaa;
rom[74123] = 12'h999;
rom[74124] = 12'h888;
rom[74125] = 12'h888;
rom[74126] = 12'h777;
rom[74127] = 12'h777;
rom[74128] = 12'h777;
rom[74129] = 12'h777;
rom[74130] = 12'h666;
rom[74131] = 12'h666;
rom[74132] = 12'h666;
rom[74133] = 12'h666;
rom[74134] = 12'h777;
rom[74135] = 12'h777;
rom[74136] = 12'h777;
rom[74137] = 12'h777;
rom[74138] = 12'h777;
rom[74139] = 12'h777;
rom[74140] = 12'h777;
rom[74141] = 12'h777;
rom[74142] = 12'h777;
rom[74143] = 12'h777;
rom[74144] = 12'h777;
rom[74145] = 12'h666;
rom[74146] = 12'h666;
rom[74147] = 12'h666;
rom[74148] = 12'h666;
rom[74149] = 12'h555;
rom[74150] = 12'h555;
rom[74151] = 12'h555;
rom[74152] = 12'h555;
rom[74153] = 12'h555;
rom[74154] = 12'h555;
rom[74155] = 12'h555;
rom[74156] = 12'h555;
rom[74157] = 12'h555;
rom[74158] = 12'h555;
rom[74159] = 12'h555;
rom[74160] = 12'h555;
rom[74161] = 12'h555;
rom[74162] = 12'h555;
rom[74163] = 12'h555;
rom[74164] = 12'h555;
rom[74165] = 12'h555;
rom[74166] = 12'h555;
rom[74167] = 12'h555;
rom[74168] = 12'h555;
rom[74169] = 12'h555;
rom[74170] = 12'h555;
rom[74171] = 12'h555;
rom[74172] = 12'h444;
rom[74173] = 12'h444;
rom[74174] = 12'h444;
rom[74175] = 12'h444;
rom[74176] = 12'h444;
rom[74177] = 12'h444;
rom[74178] = 12'h444;
rom[74179] = 12'h444;
rom[74180] = 12'h444;
rom[74181] = 12'h444;
rom[74182] = 12'h555;
rom[74183] = 12'h555;
rom[74184] = 12'h666;
rom[74185] = 12'h555;
rom[74186] = 12'h555;
rom[74187] = 12'h555;
rom[74188] = 12'h555;
rom[74189] = 12'h444;
rom[74190] = 12'h444;
rom[74191] = 12'h444;
rom[74192] = 12'h333;
rom[74193] = 12'h333;
rom[74194] = 12'h333;
rom[74195] = 12'h333;
rom[74196] = 12'h444;
rom[74197] = 12'h555;
rom[74198] = 12'h555;
rom[74199] = 12'h444;
rom[74200] = 12'h333;
rom[74201] = 12'h333;
rom[74202] = 12'h333;
rom[74203] = 12'h333;
rom[74204] = 12'h222;
rom[74205] = 12'h222;
rom[74206] = 12'h222;
rom[74207] = 12'h333;
rom[74208] = 12'h333;
rom[74209] = 12'h333;
rom[74210] = 12'h222;
rom[74211] = 12'h111;
rom[74212] = 12'h111;
rom[74213] = 12'h111;
rom[74214] = 12'h111;
rom[74215] = 12'h111;
rom[74216] = 12'h111;
rom[74217] = 12'h111;
rom[74218] = 12'h111;
rom[74219] = 12'h  0;
rom[74220] = 12'h  0;
rom[74221] = 12'h  0;
rom[74222] = 12'h111;
rom[74223] = 12'h111;
rom[74224] = 12'h111;
rom[74225] = 12'h111;
rom[74226] = 12'h111;
rom[74227] = 12'h111;
rom[74228] = 12'h111;
rom[74229] = 12'h111;
rom[74230] = 12'h111;
rom[74231] = 12'h111;
rom[74232] = 12'h111;
rom[74233] = 12'h  0;
rom[74234] = 12'h  0;
rom[74235] = 12'h  0;
rom[74236] = 12'h  0;
rom[74237] = 12'h  0;
rom[74238] = 12'h  0;
rom[74239] = 12'h  0;
rom[74240] = 12'h  0;
rom[74241] = 12'h  0;
rom[74242] = 12'h  0;
rom[74243] = 12'h  0;
rom[74244] = 12'h  0;
rom[74245] = 12'h  0;
rom[74246] = 12'h  0;
rom[74247] = 12'h  0;
rom[74248] = 12'h  0;
rom[74249] = 12'h  0;
rom[74250] = 12'h  0;
rom[74251] = 12'h  0;
rom[74252] = 12'h  0;
rom[74253] = 12'h  0;
rom[74254] = 12'h  0;
rom[74255] = 12'h  0;
rom[74256] = 12'h  0;
rom[74257] = 12'h  0;
rom[74258] = 12'h  0;
rom[74259] = 12'h  0;
rom[74260] = 12'h  0;
rom[74261] = 12'h  0;
rom[74262] = 12'h  0;
rom[74263] = 12'h  0;
rom[74264] = 12'h  0;
rom[74265] = 12'h  0;
rom[74266] = 12'h  0;
rom[74267] = 12'h  0;
rom[74268] = 12'h  0;
rom[74269] = 12'h  0;
rom[74270] = 12'h111;
rom[74271] = 12'h111;
rom[74272] = 12'h111;
rom[74273] = 12'h111;
rom[74274] = 12'h222;
rom[74275] = 12'h333;
rom[74276] = 12'h333;
rom[74277] = 12'h444;
rom[74278] = 12'h555;
rom[74279] = 12'h777;
rom[74280] = 12'h666;
rom[74281] = 12'h555;
rom[74282] = 12'h333;
rom[74283] = 12'h222;
rom[74284] = 12'h222;
rom[74285] = 12'h222;
rom[74286] = 12'h111;
rom[74287] = 12'h111;
rom[74288] = 12'h111;
rom[74289] = 12'h111;
rom[74290] = 12'h111;
rom[74291] = 12'h111;
rom[74292] = 12'h111;
rom[74293] = 12'h111;
rom[74294] = 12'h111;
rom[74295] = 12'h111;
rom[74296] = 12'h222;
rom[74297] = 12'h222;
rom[74298] = 12'h222;
rom[74299] = 12'h222;
rom[74300] = 12'h222;
rom[74301] = 12'h333;
rom[74302] = 12'h333;
rom[74303] = 12'h333;
rom[74304] = 12'h444;
rom[74305] = 12'h444;
rom[74306] = 12'h555;
rom[74307] = 12'h555;
rom[74308] = 12'h555;
rom[74309] = 12'h666;
rom[74310] = 12'h666;
rom[74311] = 12'h777;
rom[74312] = 12'h777;
rom[74313] = 12'h777;
rom[74314] = 12'h888;
rom[74315] = 12'haaa;
rom[74316] = 12'hbbb;
rom[74317] = 12'hbbb;
rom[74318] = 12'hbbb;
rom[74319] = 12'hccc;
rom[74320] = 12'hccc;
rom[74321] = 12'hccc;
rom[74322] = 12'hddd;
rom[74323] = 12'heee;
rom[74324] = 12'heee;
rom[74325] = 12'hfff;
rom[74326] = 12'hfff;
rom[74327] = 12'hfff;
rom[74328] = 12'hfff;
rom[74329] = 12'hfff;
rom[74330] = 12'hfff;
rom[74331] = 12'hfff;
rom[74332] = 12'hfff;
rom[74333] = 12'hfff;
rom[74334] = 12'heee;
rom[74335] = 12'heee;
rom[74336] = 12'hccc;
rom[74337] = 12'hccc;
rom[74338] = 12'hbbb;
rom[74339] = 12'haaa;
rom[74340] = 12'haaa;
rom[74341] = 12'haaa;
rom[74342] = 12'h999;
rom[74343] = 12'h999;
rom[74344] = 12'h999;
rom[74345] = 12'h999;
rom[74346] = 12'h999;
rom[74347] = 12'h999;
rom[74348] = 12'h999;
rom[74349] = 12'h888;
rom[74350] = 12'h777;
rom[74351] = 12'h777;
rom[74352] = 12'h666;
rom[74353] = 12'h666;
rom[74354] = 12'h666;
rom[74355] = 12'h555;
rom[74356] = 12'h555;
rom[74357] = 12'h666;
rom[74358] = 12'h666;
rom[74359] = 12'h666;
rom[74360] = 12'h555;
rom[74361] = 12'h555;
rom[74362] = 12'h555;
rom[74363] = 12'h555;
rom[74364] = 12'h555;
rom[74365] = 12'h555;
rom[74366] = 12'h555;
rom[74367] = 12'h444;
rom[74368] = 12'h444;
rom[74369] = 12'h444;
rom[74370] = 12'h444;
rom[74371] = 12'h444;
rom[74372] = 12'h444;
rom[74373] = 12'h444;
rom[74374] = 12'h444;
rom[74375] = 12'h444;
rom[74376] = 12'h444;
rom[74377] = 12'h444;
rom[74378] = 12'h444;
rom[74379] = 12'h444;
rom[74380] = 12'h444;
rom[74381] = 12'h444;
rom[74382] = 12'h444;
rom[74383] = 12'h444;
rom[74384] = 12'h444;
rom[74385] = 12'h444;
rom[74386] = 12'h444;
rom[74387] = 12'h444;
rom[74388] = 12'h444;
rom[74389] = 12'h555;
rom[74390] = 12'h555;
rom[74391] = 12'h555;
rom[74392] = 12'h666;
rom[74393] = 12'h666;
rom[74394] = 12'h666;
rom[74395] = 12'h555;
rom[74396] = 12'h555;
rom[74397] = 12'h555;
rom[74398] = 12'h555;
rom[74399] = 12'h555;
rom[74400] = 12'hfff;
rom[74401] = 12'hfff;
rom[74402] = 12'hfff;
rom[74403] = 12'hfff;
rom[74404] = 12'hfff;
rom[74405] = 12'hfff;
rom[74406] = 12'hfff;
rom[74407] = 12'hfff;
rom[74408] = 12'hfff;
rom[74409] = 12'hfff;
rom[74410] = 12'hfff;
rom[74411] = 12'hfff;
rom[74412] = 12'hfff;
rom[74413] = 12'hfff;
rom[74414] = 12'hfff;
rom[74415] = 12'hfff;
rom[74416] = 12'hfff;
rom[74417] = 12'hfff;
rom[74418] = 12'hfff;
rom[74419] = 12'hfff;
rom[74420] = 12'hfff;
rom[74421] = 12'hfff;
rom[74422] = 12'hfff;
rom[74423] = 12'hfff;
rom[74424] = 12'hfff;
rom[74425] = 12'hfff;
rom[74426] = 12'hfff;
rom[74427] = 12'hfff;
rom[74428] = 12'hfff;
rom[74429] = 12'hfff;
rom[74430] = 12'hfff;
rom[74431] = 12'hfff;
rom[74432] = 12'hfff;
rom[74433] = 12'hfff;
rom[74434] = 12'hfff;
rom[74435] = 12'hfff;
rom[74436] = 12'hfff;
rom[74437] = 12'hfff;
rom[74438] = 12'hfff;
rom[74439] = 12'hfff;
rom[74440] = 12'hfff;
rom[74441] = 12'hfff;
rom[74442] = 12'hfff;
rom[74443] = 12'hfff;
rom[74444] = 12'hfff;
rom[74445] = 12'hfff;
rom[74446] = 12'hfff;
rom[74447] = 12'hfff;
rom[74448] = 12'hfff;
rom[74449] = 12'hfff;
rom[74450] = 12'hfff;
rom[74451] = 12'hfff;
rom[74452] = 12'hfff;
rom[74453] = 12'hfff;
rom[74454] = 12'hfff;
rom[74455] = 12'hfff;
rom[74456] = 12'hfff;
rom[74457] = 12'hfff;
rom[74458] = 12'hfff;
rom[74459] = 12'hfff;
rom[74460] = 12'hfff;
rom[74461] = 12'hfff;
rom[74462] = 12'hfff;
rom[74463] = 12'hfff;
rom[74464] = 12'hfff;
rom[74465] = 12'hfff;
rom[74466] = 12'hfff;
rom[74467] = 12'hfff;
rom[74468] = 12'hfff;
rom[74469] = 12'hfff;
rom[74470] = 12'hfff;
rom[74471] = 12'hfff;
rom[74472] = 12'hfff;
rom[74473] = 12'hfff;
rom[74474] = 12'hfff;
rom[74475] = 12'hfff;
rom[74476] = 12'hfff;
rom[74477] = 12'hfff;
rom[74478] = 12'hfff;
rom[74479] = 12'hfff;
rom[74480] = 12'hfff;
rom[74481] = 12'hfff;
rom[74482] = 12'hfff;
rom[74483] = 12'hfff;
rom[74484] = 12'hfff;
rom[74485] = 12'hfff;
rom[74486] = 12'hfff;
rom[74487] = 12'hfff;
rom[74488] = 12'hfff;
rom[74489] = 12'hfff;
rom[74490] = 12'hfff;
rom[74491] = 12'hfff;
rom[74492] = 12'hfff;
rom[74493] = 12'hfff;
rom[74494] = 12'hfff;
rom[74495] = 12'hfff;
rom[74496] = 12'hfff;
rom[74497] = 12'hfff;
rom[74498] = 12'hfff;
rom[74499] = 12'hfff;
rom[74500] = 12'hfff;
rom[74501] = 12'hfff;
rom[74502] = 12'hfff;
rom[74503] = 12'hfff;
rom[74504] = 12'hfff;
rom[74505] = 12'hfff;
rom[74506] = 12'hfff;
rom[74507] = 12'hfff;
rom[74508] = 12'hfff;
rom[74509] = 12'hfff;
rom[74510] = 12'hfff;
rom[74511] = 12'heee;
rom[74512] = 12'heee;
rom[74513] = 12'heee;
rom[74514] = 12'hddd;
rom[74515] = 12'hddd;
rom[74516] = 12'hddd;
rom[74517] = 12'hddd;
rom[74518] = 12'hccc;
rom[74519] = 12'hccc;
rom[74520] = 12'hccc;
rom[74521] = 12'hbbb;
rom[74522] = 12'hbbb;
rom[74523] = 12'haaa;
rom[74524] = 12'h999;
rom[74525] = 12'h999;
rom[74526] = 12'h888;
rom[74527] = 12'h888;
rom[74528] = 12'h777;
rom[74529] = 12'h777;
rom[74530] = 12'h777;
rom[74531] = 12'h666;
rom[74532] = 12'h666;
rom[74533] = 12'h666;
rom[74534] = 12'h666;
rom[74535] = 12'h666;
rom[74536] = 12'h777;
rom[74537] = 12'h777;
rom[74538] = 12'h777;
rom[74539] = 12'h777;
rom[74540] = 12'h777;
rom[74541] = 12'h777;
rom[74542] = 12'h777;
rom[74543] = 12'h777;
rom[74544] = 12'h777;
rom[74545] = 12'h777;
rom[74546] = 12'h777;
rom[74547] = 12'h777;
rom[74548] = 12'h777;
rom[74549] = 12'h777;
rom[74550] = 12'h666;
rom[74551] = 12'h666;
rom[74552] = 12'h666;
rom[74553] = 12'h666;
rom[74554] = 12'h666;
rom[74555] = 12'h555;
rom[74556] = 12'h555;
rom[74557] = 12'h555;
rom[74558] = 12'h555;
rom[74559] = 12'h555;
rom[74560] = 12'h555;
rom[74561] = 12'h555;
rom[74562] = 12'h555;
rom[74563] = 12'h555;
rom[74564] = 12'h555;
rom[74565] = 12'h555;
rom[74566] = 12'h555;
rom[74567] = 12'h555;
rom[74568] = 12'h555;
rom[74569] = 12'h555;
rom[74570] = 12'h555;
rom[74571] = 12'h444;
rom[74572] = 12'h444;
rom[74573] = 12'h444;
rom[74574] = 12'h444;
rom[74575] = 12'h444;
rom[74576] = 12'h444;
rom[74577] = 12'h444;
rom[74578] = 12'h444;
rom[74579] = 12'h444;
rom[74580] = 12'h444;
rom[74581] = 12'h444;
rom[74582] = 12'h444;
rom[74583] = 12'h444;
rom[74584] = 12'h555;
rom[74585] = 12'h555;
rom[74586] = 12'h666;
rom[74587] = 12'h666;
rom[74588] = 12'h666;
rom[74589] = 12'h555;
rom[74590] = 12'h555;
rom[74591] = 12'h444;
rom[74592] = 12'h444;
rom[74593] = 12'h444;
rom[74594] = 12'h333;
rom[74595] = 12'h333;
rom[74596] = 12'h444;
rom[74597] = 12'h555;
rom[74598] = 12'h555;
rom[74599] = 12'h555;
rom[74600] = 12'h444;
rom[74601] = 12'h444;
rom[74602] = 12'h333;
rom[74603] = 12'h333;
rom[74604] = 12'h333;
rom[74605] = 12'h333;
rom[74606] = 12'h333;
rom[74607] = 12'h333;
rom[74608] = 12'h333;
rom[74609] = 12'h333;
rom[74610] = 12'h222;
rom[74611] = 12'h222;
rom[74612] = 12'h111;
rom[74613] = 12'h111;
rom[74614] = 12'h111;
rom[74615] = 12'h111;
rom[74616] = 12'h111;
rom[74617] = 12'h111;
rom[74618] = 12'h111;
rom[74619] = 12'h111;
rom[74620] = 12'h  0;
rom[74621] = 12'h111;
rom[74622] = 12'h111;
rom[74623] = 12'h111;
rom[74624] = 12'h111;
rom[74625] = 12'h111;
rom[74626] = 12'h111;
rom[74627] = 12'h111;
rom[74628] = 12'h111;
rom[74629] = 12'h111;
rom[74630] = 12'h111;
rom[74631] = 12'h111;
rom[74632] = 12'h111;
rom[74633] = 12'h  0;
rom[74634] = 12'h  0;
rom[74635] = 12'h  0;
rom[74636] = 12'h  0;
rom[74637] = 12'h  0;
rom[74638] = 12'h  0;
rom[74639] = 12'h  0;
rom[74640] = 12'h  0;
rom[74641] = 12'h  0;
rom[74642] = 12'h  0;
rom[74643] = 12'h  0;
rom[74644] = 12'h  0;
rom[74645] = 12'h  0;
rom[74646] = 12'h  0;
rom[74647] = 12'h  0;
rom[74648] = 12'h  0;
rom[74649] = 12'h  0;
rom[74650] = 12'h  0;
rom[74651] = 12'h  0;
rom[74652] = 12'h  0;
rom[74653] = 12'h  0;
rom[74654] = 12'h  0;
rom[74655] = 12'h  0;
rom[74656] = 12'h  0;
rom[74657] = 12'h  0;
rom[74658] = 12'h  0;
rom[74659] = 12'h  0;
rom[74660] = 12'h  0;
rom[74661] = 12'h  0;
rom[74662] = 12'h  0;
rom[74663] = 12'h  0;
rom[74664] = 12'h  0;
rom[74665] = 12'h  0;
rom[74666] = 12'h  0;
rom[74667] = 12'h  0;
rom[74668] = 12'h  0;
rom[74669] = 12'h  0;
rom[74670] = 12'h111;
rom[74671] = 12'h111;
rom[74672] = 12'h111;
rom[74673] = 12'h111;
rom[74674] = 12'h222;
rom[74675] = 12'h333;
rom[74676] = 12'h333;
rom[74677] = 12'h444;
rom[74678] = 12'h666;
rom[74679] = 12'h777;
rom[74680] = 12'h666;
rom[74681] = 12'h555;
rom[74682] = 12'h333;
rom[74683] = 12'h222;
rom[74684] = 12'h222;
rom[74685] = 12'h222;
rom[74686] = 12'h111;
rom[74687] = 12'h111;
rom[74688] = 12'h111;
rom[74689] = 12'h111;
rom[74690] = 12'h111;
rom[74691] = 12'h111;
rom[74692] = 12'h111;
rom[74693] = 12'h111;
rom[74694] = 12'h111;
rom[74695] = 12'h111;
rom[74696] = 12'h222;
rom[74697] = 12'h222;
rom[74698] = 12'h222;
rom[74699] = 12'h222;
rom[74700] = 12'h333;
rom[74701] = 12'h333;
rom[74702] = 12'h333;
rom[74703] = 12'h444;
rom[74704] = 12'h444;
rom[74705] = 12'h444;
rom[74706] = 12'h555;
rom[74707] = 12'h555;
rom[74708] = 12'h555;
rom[74709] = 12'h666;
rom[74710] = 12'h666;
rom[74711] = 12'h777;
rom[74712] = 12'h777;
rom[74713] = 12'h888;
rom[74714] = 12'h999;
rom[74715] = 12'haaa;
rom[74716] = 12'hbbb;
rom[74717] = 12'hbbb;
rom[74718] = 12'hccc;
rom[74719] = 12'hccc;
rom[74720] = 12'hddd;
rom[74721] = 12'hddd;
rom[74722] = 12'heee;
rom[74723] = 12'heee;
rom[74724] = 12'hfff;
rom[74725] = 12'hfff;
rom[74726] = 12'hfff;
rom[74727] = 12'hfff;
rom[74728] = 12'hfff;
rom[74729] = 12'hfff;
rom[74730] = 12'hfff;
rom[74731] = 12'hfff;
rom[74732] = 12'hfff;
rom[74733] = 12'heee;
rom[74734] = 12'hddd;
rom[74735] = 12'hddd;
rom[74736] = 12'hbbb;
rom[74737] = 12'hbbb;
rom[74738] = 12'haaa;
rom[74739] = 12'haaa;
rom[74740] = 12'haaa;
rom[74741] = 12'h999;
rom[74742] = 12'h999;
rom[74743] = 12'h999;
rom[74744] = 12'h888;
rom[74745] = 12'h999;
rom[74746] = 12'h999;
rom[74747] = 12'h999;
rom[74748] = 12'h888;
rom[74749] = 12'h888;
rom[74750] = 12'h777;
rom[74751] = 12'h777;
rom[74752] = 12'h666;
rom[74753] = 12'h666;
rom[74754] = 12'h555;
rom[74755] = 12'h555;
rom[74756] = 12'h555;
rom[74757] = 12'h555;
rom[74758] = 12'h555;
rom[74759] = 12'h555;
rom[74760] = 12'h555;
rom[74761] = 12'h555;
rom[74762] = 12'h555;
rom[74763] = 12'h555;
rom[74764] = 12'h555;
rom[74765] = 12'h555;
rom[74766] = 12'h555;
rom[74767] = 12'h444;
rom[74768] = 12'h444;
rom[74769] = 12'h444;
rom[74770] = 12'h444;
rom[74771] = 12'h444;
rom[74772] = 12'h444;
rom[74773] = 12'h444;
rom[74774] = 12'h444;
rom[74775] = 12'h444;
rom[74776] = 12'h444;
rom[74777] = 12'h444;
rom[74778] = 12'h444;
rom[74779] = 12'h444;
rom[74780] = 12'h444;
rom[74781] = 12'h444;
rom[74782] = 12'h444;
rom[74783] = 12'h444;
rom[74784] = 12'h444;
rom[74785] = 12'h444;
rom[74786] = 12'h444;
rom[74787] = 12'h444;
rom[74788] = 12'h444;
rom[74789] = 12'h444;
rom[74790] = 12'h444;
rom[74791] = 12'h555;
rom[74792] = 12'h555;
rom[74793] = 12'h555;
rom[74794] = 12'h666;
rom[74795] = 12'h555;
rom[74796] = 12'h555;
rom[74797] = 12'h555;
rom[74798] = 12'h555;
rom[74799] = 12'h555;
rom[74800] = 12'hfff;
rom[74801] = 12'hfff;
rom[74802] = 12'hfff;
rom[74803] = 12'hfff;
rom[74804] = 12'hfff;
rom[74805] = 12'hfff;
rom[74806] = 12'hfff;
rom[74807] = 12'hfff;
rom[74808] = 12'hfff;
rom[74809] = 12'hfff;
rom[74810] = 12'hfff;
rom[74811] = 12'hfff;
rom[74812] = 12'hfff;
rom[74813] = 12'hfff;
rom[74814] = 12'hfff;
rom[74815] = 12'hfff;
rom[74816] = 12'hfff;
rom[74817] = 12'hfff;
rom[74818] = 12'hfff;
rom[74819] = 12'hfff;
rom[74820] = 12'hfff;
rom[74821] = 12'hfff;
rom[74822] = 12'hfff;
rom[74823] = 12'hfff;
rom[74824] = 12'hfff;
rom[74825] = 12'hfff;
rom[74826] = 12'hfff;
rom[74827] = 12'hfff;
rom[74828] = 12'hfff;
rom[74829] = 12'hfff;
rom[74830] = 12'hfff;
rom[74831] = 12'hfff;
rom[74832] = 12'hfff;
rom[74833] = 12'hfff;
rom[74834] = 12'hfff;
rom[74835] = 12'hfff;
rom[74836] = 12'hfff;
rom[74837] = 12'hfff;
rom[74838] = 12'hfff;
rom[74839] = 12'hfff;
rom[74840] = 12'hfff;
rom[74841] = 12'hfff;
rom[74842] = 12'hfff;
rom[74843] = 12'hfff;
rom[74844] = 12'hfff;
rom[74845] = 12'hfff;
rom[74846] = 12'hfff;
rom[74847] = 12'hfff;
rom[74848] = 12'hfff;
rom[74849] = 12'hfff;
rom[74850] = 12'hfff;
rom[74851] = 12'hfff;
rom[74852] = 12'hfff;
rom[74853] = 12'hfff;
rom[74854] = 12'hfff;
rom[74855] = 12'hfff;
rom[74856] = 12'hfff;
rom[74857] = 12'hfff;
rom[74858] = 12'hfff;
rom[74859] = 12'hfff;
rom[74860] = 12'hfff;
rom[74861] = 12'hfff;
rom[74862] = 12'hfff;
rom[74863] = 12'hfff;
rom[74864] = 12'hfff;
rom[74865] = 12'hfff;
rom[74866] = 12'hfff;
rom[74867] = 12'hfff;
rom[74868] = 12'hfff;
rom[74869] = 12'hfff;
rom[74870] = 12'hfff;
rom[74871] = 12'hfff;
rom[74872] = 12'hfff;
rom[74873] = 12'hfff;
rom[74874] = 12'hfff;
rom[74875] = 12'hfff;
rom[74876] = 12'hfff;
rom[74877] = 12'hfff;
rom[74878] = 12'hfff;
rom[74879] = 12'hfff;
rom[74880] = 12'hfff;
rom[74881] = 12'hfff;
rom[74882] = 12'hfff;
rom[74883] = 12'hfff;
rom[74884] = 12'hfff;
rom[74885] = 12'hfff;
rom[74886] = 12'hfff;
rom[74887] = 12'hfff;
rom[74888] = 12'hfff;
rom[74889] = 12'hfff;
rom[74890] = 12'hfff;
rom[74891] = 12'hfff;
rom[74892] = 12'hfff;
rom[74893] = 12'hfff;
rom[74894] = 12'hfff;
rom[74895] = 12'hfff;
rom[74896] = 12'hfff;
rom[74897] = 12'hfff;
rom[74898] = 12'hfff;
rom[74899] = 12'hfff;
rom[74900] = 12'hfff;
rom[74901] = 12'hfff;
rom[74902] = 12'hfff;
rom[74903] = 12'hfff;
rom[74904] = 12'hfff;
rom[74905] = 12'hfff;
rom[74906] = 12'hfff;
rom[74907] = 12'hfff;
rom[74908] = 12'hfff;
rom[74909] = 12'hfff;
rom[74910] = 12'hfff;
rom[74911] = 12'heee;
rom[74912] = 12'heee;
rom[74913] = 12'hddd;
rom[74914] = 12'hccc;
rom[74915] = 12'hccc;
rom[74916] = 12'hbbb;
rom[74917] = 12'hbbb;
rom[74918] = 12'hbbb;
rom[74919] = 12'hbbb;
rom[74920] = 12'hbbb;
rom[74921] = 12'hbbb;
rom[74922] = 12'haaa;
rom[74923] = 12'haaa;
rom[74924] = 12'haaa;
rom[74925] = 12'haaa;
rom[74926] = 12'h999;
rom[74927] = 12'h999;
rom[74928] = 12'h888;
rom[74929] = 12'h888;
rom[74930] = 12'h888;
rom[74931] = 12'h777;
rom[74932] = 12'h777;
rom[74933] = 12'h666;
rom[74934] = 12'h666;
rom[74935] = 12'h666;
rom[74936] = 12'h666;
rom[74937] = 12'h666;
rom[74938] = 12'h666;
rom[74939] = 12'h666;
rom[74940] = 12'h666;
rom[74941] = 12'h666;
rom[74942] = 12'h666;
rom[74943] = 12'h777;
rom[74944] = 12'h777;
rom[74945] = 12'h777;
rom[74946] = 12'h777;
rom[74947] = 12'h777;
rom[74948] = 12'h777;
rom[74949] = 12'h777;
rom[74950] = 12'h777;
rom[74951] = 12'h777;
rom[74952] = 12'h777;
rom[74953] = 12'h777;
rom[74954] = 12'h777;
rom[74955] = 12'h666;
rom[74956] = 12'h666;
rom[74957] = 12'h666;
rom[74958] = 12'h555;
rom[74959] = 12'h555;
rom[74960] = 12'h555;
rom[74961] = 12'h555;
rom[74962] = 12'h555;
rom[74963] = 12'h555;
rom[74964] = 12'h555;
rom[74965] = 12'h555;
rom[74966] = 12'h555;
rom[74967] = 12'h555;
rom[74968] = 12'h555;
rom[74969] = 12'h555;
rom[74970] = 12'h555;
rom[74971] = 12'h444;
rom[74972] = 12'h444;
rom[74973] = 12'h444;
rom[74974] = 12'h444;
rom[74975] = 12'h444;
rom[74976] = 12'h444;
rom[74977] = 12'h444;
rom[74978] = 12'h444;
rom[74979] = 12'h444;
rom[74980] = 12'h444;
rom[74981] = 12'h444;
rom[74982] = 12'h444;
rom[74983] = 12'h444;
rom[74984] = 12'h444;
rom[74985] = 12'h555;
rom[74986] = 12'h555;
rom[74987] = 12'h666;
rom[74988] = 12'h666;
rom[74989] = 12'h666;
rom[74990] = 12'h555;
rom[74991] = 12'h555;
rom[74992] = 12'h555;
rom[74993] = 12'h444;
rom[74994] = 12'h444;
rom[74995] = 12'h333;
rom[74996] = 12'h444;
rom[74997] = 12'h555;
rom[74998] = 12'h666;
rom[74999] = 12'h555;
rom[75000] = 12'h444;
rom[75001] = 12'h444;
rom[75002] = 12'h444;
rom[75003] = 12'h444;
rom[75004] = 12'h333;
rom[75005] = 12'h333;
rom[75006] = 12'h333;
rom[75007] = 12'h444;
rom[75008] = 12'h444;
rom[75009] = 12'h333;
rom[75010] = 12'h222;
rom[75011] = 12'h222;
rom[75012] = 12'h111;
rom[75013] = 12'h111;
rom[75014] = 12'h222;
rom[75015] = 12'h111;
rom[75016] = 12'h111;
rom[75017] = 12'h111;
rom[75018] = 12'h111;
rom[75019] = 12'h111;
rom[75020] = 12'h111;
rom[75021] = 12'h111;
rom[75022] = 12'h111;
rom[75023] = 12'h111;
rom[75024] = 12'h111;
rom[75025] = 12'h111;
rom[75026] = 12'h111;
rom[75027] = 12'h111;
rom[75028] = 12'h111;
rom[75029] = 12'h111;
rom[75030] = 12'h111;
rom[75031] = 12'h111;
rom[75032] = 12'h111;
rom[75033] = 12'h111;
rom[75034] = 12'h  0;
rom[75035] = 12'h  0;
rom[75036] = 12'h  0;
rom[75037] = 12'h  0;
rom[75038] = 12'h  0;
rom[75039] = 12'h  0;
rom[75040] = 12'h  0;
rom[75041] = 12'h  0;
rom[75042] = 12'h  0;
rom[75043] = 12'h  0;
rom[75044] = 12'h  0;
rom[75045] = 12'h  0;
rom[75046] = 12'h  0;
rom[75047] = 12'h  0;
rom[75048] = 12'h  0;
rom[75049] = 12'h  0;
rom[75050] = 12'h  0;
rom[75051] = 12'h  0;
rom[75052] = 12'h  0;
rom[75053] = 12'h  0;
rom[75054] = 12'h  0;
rom[75055] = 12'h  0;
rom[75056] = 12'h  0;
rom[75057] = 12'h  0;
rom[75058] = 12'h  0;
rom[75059] = 12'h  0;
rom[75060] = 12'h  0;
rom[75061] = 12'h  0;
rom[75062] = 12'h  0;
rom[75063] = 12'h  0;
rom[75064] = 12'h  0;
rom[75065] = 12'h  0;
rom[75066] = 12'h  0;
rom[75067] = 12'h  0;
rom[75068] = 12'h  0;
rom[75069] = 12'h  0;
rom[75070] = 12'h111;
rom[75071] = 12'h111;
rom[75072] = 12'h111;
rom[75073] = 12'h111;
rom[75074] = 12'h222;
rom[75075] = 12'h333;
rom[75076] = 12'h444;
rom[75077] = 12'h444;
rom[75078] = 12'h666;
rom[75079] = 12'h777;
rom[75080] = 12'h777;
rom[75081] = 12'h555;
rom[75082] = 12'h333;
rom[75083] = 12'h222;
rom[75084] = 12'h222;
rom[75085] = 12'h222;
rom[75086] = 12'h222;
rom[75087] = 12'h222;
rom[75088] = 12'h111;
rom[75089] = 12'h111;
rom[75090] = 12'h111;
rom[75091] = 12'h111;
rom[75092] = 12'h222;
rom[75093] = 12'h222;
rom[75094] = 12'h222;
rom[75095] = 12'h222;
rom[75096] = 12'h222;
rom[75097] = 12'h222;
rom[75098] = 12'h222;
rom[75099] = 12'h333;
rom[75100] = 12'h333;
rom[75101] = 12'h333;
rom[75102] = 12'h444;
rom[75103] = 12'h444;
rom[75104] = 12'h444;
rom[75105] = 12'h444;
rom[75106] = 12'h555;
rom[75107] = 12'h555;
rom[75108] = 12'h555;
rom[75109] = 12'h666;
rom[75110] = 12'h666;
rom[75111] = 12'h777;
rom[75112] = 12'h777;
rom[75113] = 12'h888;
rom[75114] = 12'h999;
rom[75115] = 12'haaa;
rom[75116] = 12'hbbb;
rom[75117] = 12'hbbb;
rom[75118] = 12'hccc;
rom[75119] = 12'hddd;
rom[75120] = 12'hddd;
rom[75121] = 12'heee;
rom[75122] = 12'hfff;
rom[75123] = 12'hfff;
rom[75124] = 12'hfff;
rom[75125] = 12'hfff;
rom[75126] = 12'hfff;
rom[75127] = 12'hfff;
rom[75128] = 12'hfff;
rom[75129] = 12'hfff;
rom[75130] = 12'hfff;
rom[75131] = 12'hfff;
rom[75132] = 12'heee;
rom[75133] = 12'hddd;
rom[75134] = 12'hccc;
rom[75135] = 12'hccc;
rom[75136] = 12'hbbb;
rom[75137] = 12'haaa;
rom[75138] = 12'haaa;
rom[75139] = 12'h999;
rom[75140] = 12'h999;
rom[75141] = 12'h999;
rom[75142] = 12'h888;
rom[75143] = 12'h888;
rom[75144] = 12'h888;
rom[75145] = 12'h888;
rom[75146] = 12'h888;
rom[75147] = 12'h888;
rom[75148] = 12'h888;
rom[75149] = 12'h888;
rom[75150] = 12'h777;
rom[75151] = 12'h777;
rom[75152] = 12'h666;
rom[75153] = 12'h666;
rom[75154] = 12'h666;
rom[75155] = 12'h555;
rom[75156] = 12'h555;
rom[75157] = 12'h555;
rom[75158] = 12'h555;
rom[75159] = 12'h555;
rom[75160] = 12'h555;
rom[75161] = 12'h555;
rom[75162] = 12'h555;
rom[75163] = 12'h555;
rom[75164] = 12'h555;
rom[75165] = 12'h555;
rom[75166] = 12'h444;
rom[75167] = 12'h444;
rom[75168] = 12'h444;
rom[75169] = 12'h444;
rom[75170] = 12'h444;
rom[75171] = 12'h444;
rom[75172] = 12'h444;
rom[75173] = 12'h444;
rom[75174] = 12'h444;
rom[75175] = 12'h444;
rom[75176] = 12'h444;
rom[75177] = 12'h444;
rom[75178] = 12'h444;
rom[75179] = 12'h444;
rom[75180] = 12'h444;
rom[75181] = 12'h444;
rom[75182] = 12'h444;
rom[75183] = 12'h444;
rom[75184] = 12'h444;
rom[75185] = 12'h444;
rom[75186] = 12'h444;
rom[75187] = 12'h444;
rom[75188] = 12'h444;
rom[75189] = 12'h444;
rom[75190] = 12'h444;
rom[75191] = 12'h444;
rom[75192] = 12'h555;
rom[75193] = 12'h555;
rom[75194] = 12'h555;
rom[75195] = 12'h555;
rom[75196] = 12'h555;
rom[75197] = 12'h555;
rom[75198] = 12'h555;
rom[75199] = 12'h555;
rom[75200] = 12'hfff;
rom[75201] = 12'hfff;
rom[75202] = 12'hfff;
rom[75203] = 12'hfff;
rom[75204] = 12'hfff;
rom[75205] = 12'hfff;
rom[75206] = 12'hfff;
rom[75207] = 12'hfff;
rom[75208] = 12'hfff;
rom[75209] = 12'hfff;
rom[75210] = 12'hfff;
rom[75211] = 12'hfff;
rom[75212] = 12'hfff;
rom[75213] = 12'hfff;
rom[75214] = 12'hfff;
rom[75215] = 12'hfff;
rom[75216] = 12'hfff;
rom[75217] = 12'hfff;
rom[75218] = 12'hfff;
rom[75219] = 12'hfff;
rom[75220] = 12'hfff;
rom[75221] = 12'hfff;
rom[75222] = 12'hfff;
rom[75223] = 12'hfff;
rom[75224] = 12'hfff;
rom[75225] = 12'hfff;
rom[75226] = 12'hfff;
rom[75227] = 12'hfff;
rom[75228] = 12'hfff;
rom[75229] = 12'hfff;
rom[75230] = 12'hfff;
rom[75231] = 12'hfff;
rom[75232] = 12'hfff;
rom[75233] = 12'hfff;
rom[75234] = 12'hfff;
rom[75235] = 12'hfff;
rom[75236] = 12'hfff;
rom[75237] = 12'hfff;
rom[75238] = 12'hfff;
rom[75239] = 12'hfff;
rom[75240] = 12'hfff;
rom[75241] = 12'hfff;
rom[75242] = 12'hfff;
rom[75243] = 12'hfff;
rom[75244] = 12'hfff;
rom[75245] = 12'hfff;
rom[75246] = 12'hfff;
rom[75247] = 12'hfff;
rom[75248] = 12'hfff;
rom[75249] = 12'hfff;
rom[75250] = 12'hfff;
rom[75251] = 12'hfff;
rom[75252] = 12'hfff;
rom[75253] = 12'hfff;
rom[75254] = 12'hfff;
rom[75255] = 12'hfff;
rom[75256] = 12'hfff;
rom[75257] = 12'hfff;
rom[75258] = 12'hfff;
rom[75259] = 12'hfff;
rom[75260] = 12'hfff;
rom[75261] = 12'hfff;
rom[75262] = 12'hfff;
rom[75263] = 12'hfff;
rom[75264] = 12'hfff;
rom[75265] = 12'hfff;
rom[75266] = 12'hfff;
rom[75267] = 12'hfff;
rom[75268] = 12'hfff;
rom[75269] = 12'hfff;
rom[75270] = 12'hfff;
rom[75271] = 12'hfff;
rom[75272] = 12'hfff;
rom[75273] = 12'hfff;
rom[75274] = 12'hfff;
rom[75275] = 12'hfff;
rom[75276] = 12'hfff;
rom[75277] = 12'hfff;
rom[75278] = 12'hfff;
rom[75279] = 12'hfff;
rom[75280] = 12'hfff;
rom[75281] = 12'hfff;
rom[75282] = 12'hfff;
rom[75283] = 12'hfff;
rom[75284] = 12'hfff;
rom[75285] = 12'hfff;
rom[75286] = 12'hfff;
rom[75287] = 12'hfff;
rom[75288] = 12'hfff;
rom[75289] = 12'hfff;
rom[75290] = 12'hfff;
rom[75291] = 12'hfff;
rom[75292] = 12'hfff;
rom[75293] = 12'hfff;
rom[75294] = 12'hfff;
rom[75295] = 12'hfff;
rom[75296] = 12'hfff;
rom[75297] = 12'hfff;
rom[75298] = 12'hfff;
rom[75299] = 12'hfff;
rom[75300] = 12'hfff;
rom[75301] = 12'hfff;
rom[75302] = 12'hfff;
rom[75303] = 12'hfff;
rom[75304] = 12'hfff;
rom[75305] = 12'hfff;
rom[75306] = 12'hfff;
rom[75307] = 12'hfff;
rom[75308] = 12'hfff;
rom[75309] = 12'hfff;
rom[75310] = 12'hfff;
rom[75311] = 12'hfff;
rom[75312] = 12'hfff;
rom[75313] = 12'heee;
rom[75314] = 12'hddd;
rom[75315] = 12'hccc;
rom[75316] = 12'hbbb;
rom[75317] = 12'hbbb;
rom[75318] = 12'hbbb;
rom[75319] = 12'haaa;
rom[75320] = 12'haaa;
rom[75321] = 12'haaa;
rom[75322] = 12'haaa;
rom[75323] = 12'haaa;
rom[75324] = 12'haaa;
rom[75325] = 12'haaa;
rom[75326] = 12'haaa;
rom[75327] = 12'h999;
rom[75328] = 12'h999;
rom[75329] = 12'h999;
rom[75330] = 12'h888;
rom[75331] = 12'h888;
rom[75332] = 12'h888;
rom[75333] = 12'h888;
rom[75334] = 12'h777;
rom[75335] = 12'h777;
rom[75336] = 12'h666;
rom[75337] = 12'h666;
rom[75338] = 12'h666;
rom[75339] = 12'h666;
rom[75340] = 12'h666;
rom[75341] = 12'h666;
rom[75342] = 12'h666;
rom[75343] = 12'h666;
rom[75344] = 12'h666;
rom[75345] = 12'h666;
rom[75346] = 12'h666;
rom[75347] = 12'h666;
rom[75348] = 12'h777;
rom[75349] = 12'h777;
rom[75350] = 12'h777;
rom[75351] = 12'h777;
rom[75352] = 12'h777;
rom[75353] = 12'h777;
rom[75354] = 12'h777;
rom[75355] = 12'h777;
rom[75356] = 12'h777;
rom[75357] = 12'h777;
rom[75358] = 12'h777;
rom[75359] = 12'h777;
rom[75360] = 12'h666;
rom[75361] = 12'h666;
rom[75362] = 12'h666;
rom[75363] = 12'h666;
rom[75364] = 12'h666;
rom[75365] = 12'h555;
rom[75366] = 12'h555;
rom[75367] = 12'h555;
rom[75368] = 12'h555;
rom[75369] = 12'h555;
rom[75370] = 12'h444;
rom[75371] = 12'h444;
rom[75372] = 12'h444;
rom[75373] = 12'h444;
rom[75374] = 12'h444;
rom[75375] = 12'h444;
rom[75376] = 12'h444;
rom[75377] = 12'h444;
rom[75378] = 12'h444;
rom[75379] = 12'h444;
rom[75380] = 12'h444;
rom[75381] = 12'h444;
rom[75382] = 12'h444;
rom[75383] = 12'h444;
rom[75384] = 12'h444;
rom[75385] = 12'h444;
rom[75386] = 12'h444;
rom[75387] = 12'h555;
rom[75388] = 12'h555;
rom[75389] = 12'h666;
rom[75390] = 12'h666;
rom[75391] = 12'h666;
rom[75392] = 12'h666;
rom[75393] = 12'h555;
rom[75394] = 12'h444;
rom[75395] = 12'h444;
rom[75396] = 12'h444;
rom[75397] = 12'h555;
rom[75398] = 12'h666;
rom[75399] = 12'h666;
rom[75400] = 12'h555;
rom[75401] = 12'h555;
rom[75402] = 12'h444;
rom[75403] = 12'h444;
rom[75404] = 12'h444;
rom[75405] = 12'h333;
rom[75406] = 12'h333;
rom[75407] = 12'h444;
rom[75408] = 12'h444;
rom[75409] = 12'h333;
rom[75410] = 12'h222;
rom[75411] = 12'h222;
rom[75412] = 12'h222;
rom[75413] = 12'h222;
rom[75414] = 12'h222;
rom[75415] = 12'h222;
rom[75416] = 12'h111;
rom[75417] = 12'h111;
rom[75418] = 12'h111;
rom[75419] = 12'h111;
rom[75420] = 12'h111;
rom[75421] = 12'h111;
rom[75422] = 12'h111;
rom[75423] = 12'h111;
rom[75424] = 12'h111;
rom[75425] = 12'h111;
rom[75426] = 12'h111;
rom[75427] = 12'h111;
rom[75428] = 12'h111;
rom[75429] = 12'h111;
rom[75430] = 12'h111;
rom[75431] = 12'h111;
rom[75432] = 12'h111;
rom[75433] = 12'h111;
rom[75434] = 12'h  0;
rom[75435] = 12'h  0;
rom[75436] = 12'h  0;
rom[75437] = 12'h  0;
rom[75438] = 12'h  0;
rom[75439] = 12'h  0;
rom[75440] = 12'h  0;
rom[75441] = 12'h  0;
rom[75442] = 12'h  0;
rom[75443] = 12'h  0;
rom[75444] = 12'h  0;
rom[75445] = 12'h  0;
rom[75446] = 12'h  0;
rom[75447] = 12'h  0;
rom[75448] = 12'h  0;
rom[75449] = 12'h  0;
rom[75450] = 12'h  0;
rom[75451] = 12'h  0;
rom[75452] = 12'h  0;
rom[75453] = 12'h  0;
rom[75454] = 12'h  0;
rom[75455] = 12'h  0;
rom[75456] = 12'h  0;
rom[75457] = 12'h  0;
rom[75458] = 12'h  0;
rom[75459] = 12'h  0;
rom[75460] = 12'h  0;
rom[75461] = 12'h  0;
rom[75462] = 12'h  0;
rom[75463] = 12'h  0;
rom[75464] = 12'h  0;
rom[75465] = 12'h  0;
rom[75466] = 12'h  0;
rom[75467] = 12'h  0;
rom[75468] = 12'h  0;
rom[75469] = 12'h  0;
rom[75470] = 12'h111;
rom[75471] = 12'h111;
rom[75472] = 12'h111;
rom[75473] = 12'h111;
rom[75474] = 12'h222;
rom[75475] = 12'h333;
rom[75476] = 12'h444;
rom[75477] = 12'h444;
rom[75478] = 12'h666;
rom[75479] = 12'h777;
rom[75480] = 12'h777;
rom[75481] = 12'h555;
rom[75482] = 12'h333;
rom[75483] = 12'h222;
rom[75484] = 12'h222;
rom[75485] = 12'h222;
rom[75486] = 12'h222;
rom[75487] = 12'h222;
rom[75488] = 12'h222;
rom[75489] = 12'h222;
rom[75490] = 12'h222;
rom[75491] = 12'h222;
rom[75492] = 12'h222;
rom[75493] = 12'h222;
rom[75494] = 12'h222;
rom[75495] = 12'h222;
rom[75496] = 12'h222;
rom[75497] = 12'h222;
rom[75498] = 12'h333;
rom[75499] = 12'h333;
rom[75500] = 12'h333;
rom[75501] = 12'h444;
rom[75502] = 12'h444;
rom[75503] = 12'h444;
rom[75504] = 12'h444;
rom[75505] = 12'h444;
rom[75506] = 12'h555;
rom[75507] = 12'h555;
rom[75508] = 12'h555;
rom[75509] = 12'h666;
rom[75510] = 12'h666;
rom[75511] = 12'h777;
rom[75512] = 12'h777;
rom[75513] = 12'h888;
rom[75514] = 12'h999;
rom[75515] = 12'haaa;
rom[75516] = 12'hbbb;
rom[75517] = 12'hccc;
rom[75518] = 12'hccc;
rom[75519] = 12'hddd;
rom[75520] = 12'hddd;
rom[75521] = 12'heee;
rom[75522] = 12'hfff;
rom[75523] = 12'hfff;
rom[75524] = 12'hfff;
rom[75525] = 12'hfff;
rom[75526] = 12'hfff;
rom[75527] = 12'hfff;
rom[75528] = 12'hfff;
rom[75529] = 12'hfff;
rom[75530] = 12'hfff;
rom[75531] = 12'heee;
rom[75532] = 12'hddd;
rom[75533] = 12'hccc;
rom[75534] = 12'hbbb;
rom[75535] = 12'hbbb;
rom[75536] = 12'haaa;
rom[75537] = 12'haaa;
rom[75538] = 12'h999;
rom[75539] = 12'h999;
rom[75540] = 12'h888;
rom[75541] = 12'h888;
rom[75542] = 12'h888;
rom[75543] = 12'h777;
rom[75544] = 12'h777;
rom[75545] = 12'h777;
rom[75546] = 12'h777;
rom[75547] = 12'h777;
rom[75548] = 12'h777;
rom[75549] = 12'h777;
rom[75550] = 12'h777;
rom[75551] = 12'h777;
rom[75552] = 12'h777;
rom[75553] = 12'h666;
rom[75554] = 12'h666;
rom[75555] = 12'h666;
rom[75556] = 12'h555;
rom[75557] = 12'h555;
rom[75558] = 12'h555;
rom[75559] = 12'h555;
rom[75560] = 12'h555;
rom[75561] = 12'h555;
rom[75562] = 12'h555;
rom[75563] = 12'h555;
rom[75564] = 12'h555;
rom[75565] = 12'h555;
rom[75566] = 12'h444;
rom[75567] = 12'h444;
rom[75568] = 12'h444;
rom[75569] = 12'h444;
rom[75570] = 12'h444;
rom[75571] = 12'h444;
rom[75572] = 12'h444;
rom[75573] = 12'h444;
rom[75574] = 12'h444;
rom[75575] = 12'h444;
rom[75576] = 12'h444;
rom[75577] = 12'h444;
rom[75578] = 12'h444;
rom[75579] = 12'h444;
rom[75580] = 12'h444;
rom[75581] = 12'h444;
rom[75582] = 12'h444;
rom[75583] = 12'h444;
rom[75584] = 12'h444;
rom[75585] = 12'h444;
rom[75586] = 12'h444;
rom[75587] = 12'h444;
rom[75588] = 12'h444;
rom[75589] = 12'h444;
rom[75590] = 12'h444;
rom[75591] = 12'h444;
rom[75592] = 12'h444;
rom[75593] = 12'h555;
rom[75594] = 12'h555;
rom[75595] = 12'h555;
rom[75596] = 12'h555;
rom[75597] = 12'h555;
rom[75598] = 12'h444;
rom[75599] = 12'h444;
rom[75600] = 12'hfff;
rom[75601] = 12'hfff;
rom[75602] = 12'hfff;
rom[75603] = 12'hfff;
rom[75604] = 12'hfff;
rom[75605] = 12'hfff;
rom[75606] = 12'hfff;
rom[75607] = 12'hfff;
rom[75608] = 12'hfff;
rom[75609] = 12'hfff;
rom[75610] = 12'hfff;
rom[75611] = 12'hfff;
rom[75612] = 12'hfff;
rom[75613] = 12'hfff;
rom[75614] = 12'hfff;
rom[75615] = 12'hfff;
rom[75616] = 12'hfff;
rom[75617] = 12'hfff;
rom[75618] = 12'hfff;
rom[75619] = 12'hfff;
rom[75620] = 12'hfff;
rom[75621] = 12'hfff;
rom[75622] = 12'hfff;
rom[75623] = 12'hfff;
rom[75624] = 12'hfff;
rom[75625] = 12'hfff;
rom[75626] = 12'hfff;
rom[75627] = 12'hfff;
rom[75628] = 12'hfff;
rom[75629] = 12'hfff;
rom[75630] = 12'hfff;
rom[75631] = 12'hfff;
rom[75632] = 12'hfff;
rom[75633] = 12'hfff;
rom[75634] = 12'hfff;
rom[75635] = 12'hfff;
rom[75636] = 12'hfff;
rom[75637] = 12'hfff;
rom[75638] = 12'hfff;
rom[75639] = 12'hfff;
rom[75640] = 12'hfff;
rom[75641] = 12'hfff;
rom[75642] = 12'hfff;
rom[75643] = 12'hfff;
rom[75644] = 12'hfff;
rom[75645] = 12'hfff;
rom[75646] = 12'hfff;
rom[75647] = 12'hfff;
rom[75648] = 12'hfff;
rom[75649] = 12'hfff;
rom[75650] = 12'hfff;
rom[75651] = 12'hfff;
rom[75652] = 12'hfff;
rom[75653] = 12'hfff;
rom[75654] = 12'hfff;
rom[75655] = 12'hfff;
rom[75656] = 12'hfff;
rom[75657] = 12'hfff;
rom[75658] = 12'hfff;
rom[75659] = 12'hfff;
rom[75660] = 12'hfff;
rom[75661] = 12'hfff;
rom[75662] = 12'hfff;
rom[75663] = 12'hfff;
rom[75664] = 12'hfff;
rom[75665] = 12'hfff;
rom[75666] = 12'hfff;
rom[75667] = 12'hfff;
rom[75668] = 12'hfff;
rom[75669] = 12'hfff;
rom[75670] = 12'hfff;
rom[75671] = 12'hfff;
rom[75672] = 12'hfff;
rom[75673] = 12'hfff;
rom[75674] = 12'hfff;
rom[75675] = 12'hfff;
rom[75676] = 12'hfff;
rom[75677] = 12'hfff;
rom[75678] = 12'hfff;
rom[75679] = 12'hfff;
rom[75680] = 12'hfff;
rom[75681] = 12'hfff;
rom[75682] = 12'hfff;
rom[75683] = 12'hfff;
rom[75684] = 12'hfff;
rom[75685] = 12'hfff;
rom[75686] = 12'hfff;
rom[75687] = 12'hfff;
rom[75688] = 12'hfff;
rom[75689] = 12'hfff;
rom[75690] = 12'hfff;
rom[75691] = 12'hfff;
rom[75692] = 12'hfff;
rom[75693] = 12'hfff;
rom[75694] = 12'hfff;
rom[75695] = 12'hfff;
rom[75696] = 12'hfff;
rom[75697] = 12'hfff;
rom[75698] = 12'hfff;
rom[75699] = 12'hfff;
rom[75700] = 12'hfff;
rom[75701] = 12'hfff;
rom[75702] = 12'hfff;
rom[75703] = 12'hfff;
rom[75704] = 12'hfff;
rom[75705] = 12'hfff;
rom[75706] = 12'hfff;
rom[75707] = 12'hfff;
rom[75708] = 12'hfff;
rom[75709] = 12'hfff;
rom[75710] = 12'hfff;
rom[75711] = 12'hfff;
rom[75712] = 12'hfff;
rom[75713] = 12'heee;
rom[75714] = 12'hddd;
rom[75715] = 12'hddd;
rom[75716] = 12'hccc;
rom[75717] = 12'hccc;
rom[75718] = 12'hbbb;
rom[75719] = 12'haaa;
rom[75720] = 12'haaa;
rom[75721] = 12'haaa;
rom[75722] = 12'h999;
rom[75723] = 12'h999;
rom[75724] = 12'h999;
rom[75725] = 12'h999;
rom[75726] = 12'h999;
rom[75727] = 12'h888;
rom[75728] = 12'h888;
rom[75729] = 12'h888;
rom[75730] = 12'h888;
rom[75731] = 12'h888;
rom[75732] = 12'h888;
rom[75733] = 12'h888;
rom[75734] = 12'h888;
rom[75735] = 12'h888;
rom[75736] = 12'h777;
rom[75737] = 12'h777;
rom[75738] = 12'h777;
rom[75739] = 12'h777;
rom[75740] = 12'h777;
rom[75741] = 12'h777;
rom[75742] = 12'h666;
rom[75743] = 12'h666;
rom[75744] = 12'h666;
rom[75745] = 12'h666;
rom[75746] = 12'h666;
rom[75747] = 12'h666;
rom[75748] = 12'h666;
rom[75749] = 12'h777;
rom[75750] = 12'h777;
rom[75751] = 12'h777;
rom[75752] = 12'h777;
rom[75753] = 12'h777;
rom[75754] = 12'h888;
rom[75755] = 12'h888;
rom[75756] = 12'h888;
rom[75757] = 12'h888;
rom[75758] = 12'h888;
rom[75759] = 12'h888;
rom[75760] = 12'h777;
rom[75761] = 12'h777;
rom[75762] = 12'h777;
rom[75763] = 12'h777;
rom[75764] = 12'h666;
rom[75765] = 12'h666;
rom[75766] = 12'h666;
rom[75767] = 12'h555;
rom[75768] = 12'h555;
rom[75769] = 12'h555;
rom[75770] = 12'h555;
rom[75771] = 12'h444;
rom[75772] = 12'h444;
rom[75773] = 12'h444;
rom[75774] = 12'h444;
rom[75775] = 12'h444;
rom[75776] = 12'h444;
rom[75777] = 12'h444;
rom[75778] = 12'h444;
rom[75779] = 12'h444;
rom[75780] = 12'h444;
rom[75781] = 12'h444;
rom[75782] = 12'h444;
rom[75783] = 12'h444;
rom[75784] = 12'h444;
rom[75785] = 12'h444;
rom[75786] = 12'h444;
rom[75787] = 12'h444;
rom[75788] = 12'h555;
rom[75789] = 12'h555;
rom[75790] = 12'h666;
rom[75791] = 12'h666;
rom[75792] = 12'h666;
rom[75793] = 12'h666;
rom[75794] = 12'h555;
rom[75795] = 12'h555;
rom[75796] = 12'h555;
rom[75797] = 12'h555;
rom[75798] = 12'h666;
rom[75799] = 12'h666;
rom[75800] = 12'h666;
rom[75801] = 12'h555;
rom[75802] = 12'h555;
rom[75803] = 12'h555;
rom[75804] = 12'h444;
rom[75805] = 12'h444;
rom[75806] = 12'h444;
rom[75807] = 12'h444;
rom[75808] = 12'h444;
rom[75809] = 12'h333;
rom[75810] = 12'h222;
rom[75811] = 12'h222;
rom[75812] = 12'h222;
rom[75813] = 12'h222;
rom[75814] = 12'h222;
rom[75815] = 12'h222;
rom[75816] = 12'h111;
rom[75817] = 12'h111;
rom[75818] = 12'h111;
rom[75819] = 12'h111;
rom[75820] = 12'h111;
rom[75821] = 12'h111;
rom[75822] = 12'h111;
rom[75823] = 12'h111;
rom[75824] = 12'h111;
rom[75825] = 12'h111;
rom[75826] = 12'h111;
rom[75827] = 12'h111;
rom[75828] = 12'h111;
rom[75829] = 12'h111;
rom[75830] = 12'h111;
rom[75831] = 12'h111;
rom[75832] = 12'h111;
rom[75833] = 12'h111;
rom[75834] = 12'h  0;
rom[75835] = 12'h  0;
rom[75836] = 12'h  0;
rom[75837] = 12'h  0;
rom[75838] = 12'h  0;
rom[75839] = 12'h  0;
rom[75840] = 12'h  0;
rom[75841] = 12'h  0;
rom[75842] = 12'h  0;
rom[75843] = 12'h  0;
rom[75844] = 12'h  0;
rom[75845] = 12'h  0;
rom[75846] = 12'h  0;
rom[75847] = 12'h  0;
rom[75848] = 12'h  0;
rom[75849] = 12'h  0;
rom[75850] = 12'h  0;
rom[75851] = 12'h  0;
rom[75852] = 12'h  0;
rom[75853] = 12'h  0;
rom[75854] = 12'h  0;
rom[75855] = 12'h  0;
rom[75856] = 12'h  0;
rom[75857] = 12'h  0;
rom[75858] = 12'h  0;
rom[75859] = 12'h  0;
rom[75860] = 12'h  0;
rom[75861] = 12'h  0;
rom[75862] = 12'h  0;
rom[75863] = 12'h  0;
rom[75864] = 12'h  0;
rom[75865] = 12'h  0;
rom[75866] = 12'h  0;
rom[75867] = 12'h  0;
rom[75868] = 12'h  0;
rom[75869] = 12'h111;
rom[75870] = 12'h111;
rom[75871] = 12'h111;
rom[75872] = 12'h111;
rom[75873] = 12'h111;
rom[75874] = 12'h222;
rom[75875] = 12'h333;
rom[75876] = 12'h444;
rom[75877] = 12'h444;
rom[75878] = 12'h666;
rom[75879] = 12'h777;
rom[75880] = 12'h777;
rom[75881] = 12'h555;
rom[75882] = 12'h333;
rom[75883] = 12'h222;
rom[75884] = 12'h222;
rom[75885] = 12'h222;
rom[75886] = 12'h222;
rom[75887] = 12'h222;
rom[75888] = 12'h222;
rom[75889] = 12'h222;
rom[75890] = 12'h222;
rom[75891] = 12'h222;
rom[75892] = 12'h222;
rom[75893] = 12'h222;
rom[75894] = 12'h222;
rom[75895] = 12'h222;
rom[75896] = 12'h333;
rom[75897] = 12'h333;
rom[75898] = 12'h333;
rom[75899] = 12'h333;
rom[75900] = 12'h333;
rom[75901] = 12'h444;
rom[75902] = 12'h444;
rom[75903] = 12'h444;
rom[75904] = 12'h444;
rom[75905] = 12'h444;
rom[75906] = 12'h555;
rom[75907] = 12'h555;
rom[75908] = 12'h555;
rom[75909] = 12'h666;
rom[75910] = 12'h666;
rom[75911] = 12'h777;
rom[75912] = 12'h777;
rom[75913] = 12'h888;
rom[75914] = 12'h999;
rom[75915] = 12'hbbb;
rom[75916] = 12'hbbb;
rom[75917] = 12'hccc;
rom[75918] = 12'hccc;
rom[75919] = 12'hddd;
rom[75920] = 12'heee;
rom[75921] = 12'heee;
rom[75922] = 12'hfff;
rom[75923] = 12'hfff;
rom[75924] = 12'hfff;
rom[75925] = 12'hfff;
rom[75926] = 12'hfff;
rom[75927] = 12'hfff;
rom[75928] = 12'hfff;
rom[75929] = 12'heee;
rom[75930] = 12'heee;
rom[75931] = 12'hddd;
rom[75932] = 12'hccc;
rom[75933] = 12'hbbb;
rom[75934] = 12'haaa;
rom[75935] = 12'haaa;
rom[75936] = 12'h999;
rom[75937] = 12'h999;
rom[75938] = 12'h888;
rom[75939] = 12'h888;
rom[75940] = 12'h888;
rom[75941] = 12'h888;
rom[75942] = 12'h777;
rom[75943] = 12'h777;
rom[75944] = 12'h666;
rom[75945] = 12'h666;
rom[75946] = 12'h666;
rom[75947] = 12'h666;
rom[75948] = 12'h666;
rom[75949] = 12'h666;
rom[75950] = 12'h666;
rom[75951] = 12'h777;
rom[75952] = 12'h777;
rom[75953] = 12'h666;
rom[75954] = 12'h666;
rom[75955] = 12'h666;
rom[75956] = 12'h666;
rom[75957] = 12'h555;
rom[75958] = 12'h555;
rom[75959] = 12'h555;
rom[75960] = 12'h555;
rom[75961] = 12'h555;
rom[75962] = 12'h444;
rom[75963] = 12'h444;
rom[75964] = 12'h444;
rom[75965] = 12'h444;
rom[75966] = 12'h444;
rom[75967] = 12'h444;
rom[75968] = 12'h444;
rom[75969] = 12'h444;
rom[75970] = 12'h444;
rom[75971] = 12'h444;
rom[75972] = 12'h444;
rom[75973] = 12'h444;
rom[75974] = 12'h444;
rom[75975] = 12'h444;
rom[75976] = 12'h444;
rom[75977] = 12'h444;
rom[75978] = 12'h444;
rom[75979] = 12'h444;
rom[75980] = 12'h444;
rom[75981] = 12'h444;
rom[75982] = 12'h444;
rom[75983] = 12'h444;
rom[75984] = 12'h444;
rom[75985] = 12'h444;
rom[75986] = 12'h444;
rom[75987] = 12'h444;
rom[75988] = 12'h333;
rom[75989] = 12'h444;
rom[75990] = 12'h444;
rom[75991] = 12'h444;
rom[75992] = 12'h444;
rom[75993] = 12'h444;
rom[75994] = 12'h444;
rom[75995] = 12'h555;
rom[75996] = 12'h555;
rom[75997] = 12'h444;
rom[75998] = 12'h444;
rom[75999] = 12'h444;
rom[76000] = 12'hfff;
rom[76001] = 12'hfff;
rom[76002] = 12'hfff;
rom[76003] = 12'hfff;
rom[76004] = 12'hfff;
rom[76005] = 12'hfff;
rom[76006] = 12'hfff;
rom[76007] = 12'hfff;
rom[76008] = 12'hfff;
rom[76009] = 12'hfff;
rom[76010] = 12'hfff;
rom[76011] = 12'hfff;
rom[76012] = 12'hfff;
rom[76013] = 12'hfff;
rom[76014] = 12'hfff;
rom[76015] = 12'hfff;
rom[76016] = 12'hfff;
rom[76017] = 12'hfff;
rom[76018] = 12'hfff;
rom[76019] = 12'hfff;
rom[76020] = 12'hfff;
rom[76021] = 12'hfff;
rom[76022] = 12'hfff;
rom[76023] = 12'hfff;
rom[76024] = 12'hfff;
rom[76025] = 12'hfff;
rom[76026] = 12'hfff;
rom[76027] = 12'hfff;
rom[76028] = 12'hfff;
rom[76029] = 12'hfff;
rom[76030] = 12'hfff;
rom[76031] = 12'hfff;
rom[76032] = 12'hfff;
rom[76033] = 12'hfff;
rom[76034] = 12'hfff;
rom[76035] = 12'hfff;
rom[76036] = 12'hfff;
rom[76037] = 12'hfff;
rom[76038] = 12'hfff;
rom[76039] = 12'hfff;
rom[76040] = 12'hfff;
rom[76041] = 12'hfff;
rom[76042] = 12'hfff;
rom[76043] = 12'hfff;
rom[76044] = 12'hfff;
rom[76045] = 12'hfff;
rom[76046] = 12'hfff;
rom[76047] = 12'hfff;
rom[76048] = 12'hfff;
rom[76049] = 12'hfff;
rom[76050] = 12'hfff;
rom[76051] = 12'hfff;
rom[76052] = 12'hfff;
rom[76053] = 12'hfff;
rom[76054] = 12'hfff;
rom[76055] = 12'hfff;
rom[76056] = 12'hfff;
rom[76057] = 12'hfff;
rom[76058] = 12'hfff;
rom[76059] = 12'hfff;
rom[76060] = 12'hfff;
rom[76061] = 12'hfff;
rom[76062] = 12'hfff;
rom[76063] = 12'hfff;
rom[76064] = 12'hfff;
rom[76065] = 12'hfff;
rom[76066] = 12'hfff;
rom[76067] = 12'hfff;
rom[76068] = 12'hfff;
rom[76069] = 12'hfff;
rom[76070] = 12'hfff;
rom[76071] = 12'hfff;
rom[76072] = 12'hfff;
rom[76073] = 12'hfff;
rom[76074] = 12'hfff;
rom[76075] = 12'hfff;
rom[76076] = 12'hfff;
rom[76077] = 12'hfff;
rom[76078] = 12'hfff;
rom[76079] = 12'hfff;
rom[76080] = 12'hfff;
rom[76081] = 12'hfff;
rom[76082] = 12'hfff;
rom[76083] = 12'hfff;
rom[76084] = 12'hfff;
rom[76085] = 12'hfff;
rom[76086] = 12'hfff;
rom[76087] = 12'hfff;
rom[76088] = 12'hfff;
rom[76089] = 12'hfff;
rom[76090] = 12'hfff;
rom[76091] = 12'hfff;
rom[76092] = 12'hfff;
rom[76093] = 12'hfff;
rom[76094] = 12'hfff;
rom[76095] = 12'hfff;
rom[76096] = 12'hfff;
rom[76097] = 12'hfff;
rom[76098] = 12'hfff;
rom[76099] = 12'hfff;
rom[76100] = 12'hfff;
rom[76101] = 12'hfff;
rom[76102] = 12'hfff;
rom[76103] = 12'hfff;
rom[76104] = 12'hfff;
rom[76105] = 12'hfff;
rom[76106] = 12'hfff;
rom[76107] = 12'hfff;
rom[76108] = 12'hfff;
rom[76109] = 12'hfff;
rom[76110] = 12'hfff;
rom[76111] = 12'hfff;
rom[76112] = 12'hfff;
rom[76113] = 12'heee;
rom[76114] = 12'heee;
rom[76115] = 12'hddd;
rom[76116] = 12'hddd;
rom[76117] = 12'hccc;
rom[76118] = 12'hbbb;
rom[76119] = 12'hbbb;
rom[76120] = 12'haaa;
rom[76121] = 12'haaa;
rom[76122] = 12'haaa;
rom[76123] = 12'haaa;
rom[76124] = 12'h999;
rom[76125] = 12'h999;
rom[76126] = 12'h888;
rom[76127] = 12'h888;
rom[76128] = 12'h888;
rom[76129] = 12'h888;
rom[76130] = 12'h888;
rom[76131] = 12'h777;
rom[76132] = 12'h777;
rom[76133] = 12'h777;
rom[76134] = 12'h888;
rom[76135] = 12'h888;
rom[76136] = 12'h777;
rom[76137] = 12'h888;
rom[76138] = 12'h888;
rom[76139] = 12'h888;
rom[76140] = 12'h777;
rom[76141] = 12'h777;
rom[76142] = 12'h777;
rom[76143] = 12'h777;
rom[76144] = 12'h666;
rom[76145] = 12'h666;
rom[76146] = 12'h666;
rom[76147] = 12'h666;
rom[76148] = 12'h666;
rom[76149] = 12'h666;
rom[76150] = 12'h777;
rom[76151] = 12'h777;
rom[76152] = 12'h777;
rom[76153] = 12'h777;
rom[76154] = 12'h777;
rom[76155] = 12'h888;
rom[76156] = 12'h888;
rom[76157] = 12'h888;
rom[76158] = 12'h888;
rom[76159] = 12'h888;
rom[76160] = 12'h777;
rom[76161] = 12'h777;
rom[76162] = 12'h777;
rom[76163] = 12'h777;
rom[76164] = 12'h777;
rom[76165] = 12'h777;
rom[76166] = 12'h777;
rom[76167] = 12'h666;
rom[76168] = 12'h666;
rom[76169] = 12'h666;
rom[76170] = 12'h666;
rom[76171] = 12'h555;
rom[76172] = 12'h555;
rom[76173] = 12'h555;
rom[76174] = 12'h555;
rom[76175] = 12'h555;
rom[76176] = 12'h555;
rom[76177] = 12'h555;
rom[76178] = 12'h555;
rom[76179] = 12'h555;
rom[76180] = 12'h555;
rom[76181] = 12'h555;
rom[76182] = 12'h555;
rom[76183] = 12'h555;
rom[76184] = 12'h444;
rom[76185] = 12'h444;
rom[76186] = 12'h444;
rom[76187] = 12'h444;
rom[76188] = 12'h555;
rom[76189] = 12'h555;
rom[76190] = 12'h555;
rom[76191] = 12'h666;
rom[76192] = 12'h666;
rom[76193] = 12'h666;
rom[76194] = 12'h666;
rom[76195] = 12'h666;
rom[76196] = 12'h555;
rom[76197] = 12'h555;
rom[76198] = 12'h666;
rom[76199] = 12'h666;
rom[76200] = 12'h777;
rom[76201] = 12'h666;
rom[76202] = 12'h555;
rom[76203] = 12'h555;
rom[76204] = 12'h555;
rom[76205] = 12'h444;
rom[76206] = 12'h444;
rom[76207] = 12'h444;
rom[76208] = 12'h444;
rom[76209] = 12'h333;
rom[76210] = 12'h222;
rom[76211] = 12'h222;
rom[76212] = 12'h333;
rom[76213] = 12'h222;
rom[76214] = 12'h222;
rom[76215] = 12'h222;
rom[76216] = 12'h222;
rom[76217] = 12'h222;
rom[76218] = 12'h222;
rom[76219] = 12'h222;
rom[76220] = 12'h222;
rom[76221] = 12'h111;
rom[76222] = 12'h111;
rom[76223] = 12'h111;
rom[76224] = 12'h111;
rom[76225] = 12'h111;
rom[76226] = 12'h111;
rom[76227] = 12'h111;
rom[76228] = 12'h222;
rom[76229] = 12'h222;
rom[76230] = 12'h111;
rom[76231] = 12'h111;
rom[76232] = 12'h111;
rom[76233] = 12'h111;
rom[76234] = 12'h  0;
rom[76235] = 12'h  0;
rom[76236] = 12'h  0;
rom[76237] = 12'h  0;
rom[76238] = 12'h  0;
rom[76239] = 12'h  0;
rom[76240] = 12'h  0;
rom[76241] = 12'h  0;
rom[76242] = 12'h  0;
rom[76243] = 12'h  0;
rom[76244] = 12'h  0;
rom[76245] = 12'h  0;
rom[76246] = 12'h  0;
rom[76247] = 12'h  0;
rom[76248] = 12'h  0;
rom[76249] = 12'h  0;
rom[76250] = 12'h  0;
rom[76251] = 12'h  0;
rom[76252] = 12'h  0;
rom[76253] = 12'h  0;
rom[76254] = 12'h  0;
rom[76255] = 12'h  0;
rom[76256] = 12'h  0;
rom[76257] = 12'h  0;
rom[76258] = 12'h  0;
rom[76259] = 12'h  0;
rom[76260] = 12'h  0;
rom[76261] = 12'h  0;
rom[76262] = 12'h  0;
rom[76263] = 12'h  0;
rom[76264] = 12'h  0;
rom[76265] = 12'h  0;
rom[76266] = 12'h  0;
rom[76267] = 12'h  0;
rom[76268] = 12'h  0;
rom[76269] = 12'h111;
rom[76270] = 12'h111;
rom[76271] = 12'h111;
rom[76272] = 12'h111;
rom[76273] = 12'h111;
rom[76274] = 12'h222;
rom[76275] = 12'h333;
rom[76276] = 12'h333;
rom[76277] = 12'h444;
rom[76278] = 12'h666;
rom[76279] = 12'h777;
rom[76280] = 12'h777;
rom[76281] = 12'h555;
rom[76282] = 12'h333;
rom[76283] = 12'h222;
rom[76284] = 12'h222;
rom[76285] = 12'h222;
rom[76286] = 12'h222;
rom[76287] = 12'h222;
rom[76288] = 12'h222;
rom[76289] = 12'h222;
rom[76290] = 12'h222;
rom[76291] = 12'h222;
rom[76292] = 12'h222;
rom[76293] = 12'h222;
rom[76294] = 12'h333;
rom[76295] = 12'h333;
rom[76296] = 12'h333;
rom[76297] = 12'h333;
rom[76298] = 12'h333;
rom[76299] = 12'h333;
rom[76300] = 12'h333;
rom[76301] = 12'h333;
rom[76302] = 12'h444;
rom[76303] = 12'h444;
rom[76304] = 12'h444;
rom[76305] = 12'h444;
rom[76306] = 12'h555;
rom[76307] = 12'h555;
rom[76308] = 12'h666;
rom[76309] = 12'h666;
rom[76310] = 12'h777;
rom[76311] = 12'h777;
rom[76312] = 12'h888;
rom[76313] = 12'h888;
rom[76314] = 12'haaa;
rom[76315] = 12'hbbb;
rom[76316] = 12'hccc;
rom[76317] = 12'hccc;
rom[76318] = 12'hddd;
rom[76319] = 12'heee;
rom[76320] = 12'hfff;
rom[76321] = 12'hfff;
rom[76322] = 12'hfff;
rom[76323] = 12'hfff;
rom[76324] = 12'hfff;
rom[76325] = 12'hfff;
rom[76326] = 12'hfff;
rom[76327] = 12'hfff;
rom[76328] = 12'heee;
rom[76329] = 12'hddd;
rom[76330] = 12'hccc;
rom[76331] = 12'hbbb;
rom[76332] = 12'hbbb;
rom[76333] = 12'haaa;
rom[76334] = 12'haaa;
rom[76335] = 12'h999;
rom[76336] = 12'h888;
rom[76337] = 12'h888;
rom[76338] = 12'h888;
rom[76339] = 12'h777;
rom[76340] = 12'h777;
rom[76341] = 12'h777;
rom[76342] = 12'h777;
rom[76343] = 12'h777;
rom[76344] = 12'h666;
rom[76345] = 12'h666;
rom[76346] = 12'h666;
rom[76347] = 12'h555;
rom[76348] = 12'h555;
rom[76349] = 12'h666;
rom[76350] = 12'h666;
rom[76351] = 12'h666;
rom[76352] = 12'h666;
rom[76353] = 12'h666;
rom[76354] = 12'h666;
rom[76355] = 12'h666;
rom[76356] = 12'h666;
rom[76357] = 12'h555;
rom[76358] = 12'h555;
rom[76359] = 12'h555;
rom[76360] = 12'h555;
rom[76361] = 12'h444;
rom[76362] = 12'h444;
rom[76363] = 12'h444;
rom[76364] = 12'h444;
rom[76365] = 12'h444;
rom[76366] = 12'h444;
rom[76367] = 12'h444;
rom[76368] = 12'h444;
rom[76369] = 12'h444;
rom[76370] = 12'h444;
rom[76371] = 12'h444;
rom[76372] = 12'h444;
rom[76373] = 12'h444;
rom[76374] = 12'h444;
rom[76375] = 12'h444;
rom[76376] = 12'h333;
rom[76377] = 12'h333;
rom[76378] = 12'h333;
rom[76379] = 12'h333;
rom[76380] = 12'h333;
rom[76381] = 12'h333;
rom[76382] = 12'h333;
rom[76383] = 12'h333;
rom[76384] = 12'h333;
rom[76385] = 12'h333;
rom[76386] = 12'h333;
rom[76387] = 12'h333;
rom[76388] = 12'h333;
rom[76389] = 12'h333;
rom[76390] = 12'h444;
rom[76391] = 12'h444;
rom[76392] = 12'h444;
rom[76393] = 12'h444;
rom[76394] = 12'h444;
rom[76395] = 12'h444;
rom[76396] = 12'h444;
rom[76397] = 12'h444;
rom[76398] = 12'h444;
rom[76399] = 12'h444;
rom[76400] = 12'hfff;
rom[76401] = 12'hfff;
rom[76402] = 12'hfff;
rom[76403] = 12'hfff;
rom[76404] = 12'hfff;
rom[76405] = 12'hfff;
rom[76406] = 12'hfff;
rom[76407] = 12'hfff;
rom[76408] = 12'hfff;
rom[76409] = 12'hfff;
rom[76410] = 12'hfff;
rom[76411] = 12'hfff;
rom[76412] = 12'hfff;
rom[76413] = 12'hfff;
rom[76414] = 12'hfff;
rom[76415] = 12'hfff;
rom[76416] = 12'hfff;
rom[76417] = 12'hfff;
rom[76418] = 12'hfff;
rom[76419] = 12'hfff;
rom[76420] = 12'hfff;
rom[76421] = 12'hfff;
rom[76422] = 12'hfff;
rom[76423] = 12'hfff;
rom[76424] = 12'hfff;
rom[76425] = 12'hfff;
rom[76426] = 12'hfff;
rom[76427] = 12'hfff;
rom[76428] = 12'hfff;
rom[76429] = 12'hfff;
rom[76430] = 12'hfff;
rom[76431] = 12'hfff;
rom[76432] = 12'hfff;
rom[76433] = 12'hfff;
rom[76434] = 12'hfff;
rom[76435] = 12'hfff;
rom[76436] = 12'hfff;
rom[76437] = 12'hfff;
rom[76438] = 12'hfff;
rom[76439] = 12'hfff;
rom[76440] = 12'hfff;
rom[76441] = 12'hfff;
rom[76442] = 12'hfff;
rom[76443] = 12'hfff;
rom[76444] = 12'hfff;
rom[76445] = 12'hfff;
rom[76446] = 12'hfff;
rom[76447] = 12'hfff;
rom[76448] = 12'hfff;
rom[76449] = 12'hfff;
rom[76450] = 12'hfff;
rom[76451] = 12'hfff;
rom[76452] = 12'hfff;
rom[76453] = 12'hfff;
rom[76454] = 12'hfff;
rom[76455] = 12'hfff;
rom[76456] = 12'hfff;
rom[76457] = 12'hfff;
rom[76458] = 12'hfff;
rom[76459] = 12'hfff;
rom[76460] = 12'hfff;
rom[76461] = 12'hfff;
rom[76462] = 12'hfff;
rom[76463] = 12'hfff;
rom[76464] = 12'hfff;
rom[76465] = 12'hfff;
rom[76466] = 12'hfff;
rom[76467] = 12'hfff;
rom[76468] = 12'hfff;
rom[76469] = 12'hfff;
rom[76470] = 12'hfff;
rom[76471] = 12'hfff;
rom[76472] = 12'hfff;
rom[76473] = 12'hfff;
rom[76474] = 12'hfff;
rom[76475] = 12'hfff;
rom[76476] = 12'hfff;
rom[76477] = 12'hfff;
rom[76478] = 12'hfff;
rom[76479] = 12'hfff;
rom[76480] = 12'hfff;
rom[76481] = 12'hfff;
rom[76482] = 12'hfff;
rom[76483] = 12'hfff;
rom[76484] = 12'hfff;
rom[76485] = 12'hfff;
rom[76486] = 12'hfff;
rom[76487] = 12'hfff;
rom[76488] = 12'hfff;
rom[76489] = 12'hfff;
rom[76490] = 12'hfff;
rom[76491] = 12'hfff;
rom[76492] = 12'hfff;
rom[76493] = 12'hfff;
rom[76494] = 12'hfff;
rom[76495] = 12'hfff;
rom[76496] = 12'hfff;
rom[76497] = 12'hfff;
rom[76498] = 12'hfff;
rom[76499] = 12'hfff;
rom[76500] = 12'hfff;
rom[76501] = 12'hfff;
rom[76502] = 12'hfff;
rom[76503] = 12'hfff;
rom[76504] = 12'hfff;
rom[76505] = 12'hfff;
rom[76506] = 12'hfff;
rom[76507] = 12'hfff;
rom[76508] = 12'hfff;
rom[76509] = 12'hfff;
rom[76510] = 12'hfff;
rom[76511] = 12'hfff;
rom[76512] = 12'hfff;
rom[76513] = 12'hfff;
rom[76514] = 12'heee;
rom[76515] = 12'hddd;
rom[76516] = 12'hddd;
rom[76517] = 12'hccc;
rom[76518] = 12'hccc;
rom[76519] = 12'hbbb;
rom[76520] = 12'hbbb;
rom[76521] = 12'hbbb;
rom[76522] = 12'haaa;
rom[76523] = 12'haaa;
rom[76524] = 12'haaa;
rom[76525] = 12'h999;
rom[76526] = 12'h999;
rom[76527] = 12'h999;
rom[76528] = 12'h888;
rom[76529] = 12'h888;
rom[76530] = 12'h777;
rom[76531] = 12'h777;
rom[76532] = 12'h666;
rom[76533] = 12'h666;
rom[76534] = 12'h777;
rom[76535] = 12'h777;
rom[76536] = 12'h777;
rom[76537] = 12'h777;
rom[76538] = 12'h777;
rom[76539] = 12'h777;
rom[76540] = 12'h777;
rom[76541] = 12'h777;
rom[76542] = 12'h777;
rom[76543] = 12'h777;
rom[76544] = 12'h777;
rom[76545] = 12'h777;
rom[76546] = 12'h777;
rom[76547] = 12'h777;
rom[76548] = 12'h777;
rom[76549] = 12'h777;
rom[76550] = 12'h777;
rom[76551] = 12'h777;
rom[76552] = 12'h777;
rom[76553] = 12'h777;
rom[76554] = 12'h777;
rom[76555] = 12'h777;
rom[76556] = 12'h777;
rom[76557] = 12'h777;
rom[76558] = 12'h777;
rom[76559] = 12'h666;
rom[76560] = 12'h777;
rom[76561] = 12'h777;
rom[76562] = 12'h777;
rom[76563] = 12'h777;
rom[76564] = 12'h777;
rom[76565] = 12'h777;
rom[76566] = 12'h777;
rom[76567] = 12'h777;
rom[76568] = 12'h777;
rom[76569] = 12'h777;
rom[76570] = 12'h777;
rom[76571] = 12'h666;
rom[76572] = 12'h666;
rom[76573] = 12'h666;
rom[76574] = 12'h555;
rom[76575] = 12'h555;
rom[76576] = 12'h555;
rom[76577] = 12'h555;
rom[76578] = 12'h555;
rom[76579] = 12'h555;
rom[76580] = 12'h555;
rom[76581] = 12'h555;
rom[76582] = 12'h555;
rom[76583] = 12'h555;
rom[76584] = 12'h555;
rom[76585] = 12'h555;
rom[76586] = 12'h555;
rom[76587] = 12'h555;
rom[76588] = 12'h555;
rom[76589] = 12'h555;
rom[76590] = 12'h555;
rom[76591] = 12'h555;
rom[76592] = 12'h666;
rom[76593] = 12'h777;
rom[76594] = 12'h777;
rom[76595] = 12'h777;
rom[76596] = 12'h666;
rom[76597] = 12'h666;
rom[76598] = 12'h666;
rom[76599] = 12'h777;
rom[76600] = 12'h777;
rom[76601] = 12'h666;
rom[76602] = 12'h666;
rom[76603] = 12'h555;
rom[76604] = 12'h555;
rom[76605] = 12'h444;
rom[76606] = 12'h444;
rom[76607] = 12'h444;
rom[76608] = 12'h444;
rom[76609] = 12'h333;
rom[76610] = 12'h222;
rom[76611] = 12'h222;
rom[76612] = 12'h333;
rom[76613] = 12'h333;
rom[76614] = 12'h222;
rom[76615] = 12'h222;
rom[76616] = 12'h222;
rom[76617] = 12'h222;
rom[76618] = 12'h222;
rom[76619] = 12'h222;
rom[76620] = 12'h222;
rom[76621] = 12'h222;
rom[76622] = 12'h222;
rom[76623] = 12'h222;
rom[76624] = 12'h111;
rom[76625] = 12'h111;
rom[76626] = 12'h111;
rom[76627] = 12'h222;
rom[76628] = 12'h222;
rom[76629] = 12'h222;
rom[76630] = 12'h111;
rom[76631] = 12'h111;
rom[76632] = 12'h111;
rom[76633] = 12'h111;
rom[76634] = 12'h111;
rom[76635] = 12'h  0;
rom[76636] = 12'h  0;
rom[76637] = 12'h  0;
rom[76638] = 12'h  0;
rom[76639] = 12'h  0;
rom[76640] = 12'h  0;
rom[76641] = 12'h  0;
rom[76642] = 12'h  0;
rom[76643] = 12'h  0;
rom[76644] = 12'h  0;
rom[76645] = 12'h  0;
rom[76646] = 12'h  0;
rom[76647] = 12'h  0;
rom[76648] = 12'h  0;
rom[76649] = 12'h  0;
rom[76650] = 12'h  0;
rom[76651] = 12'h  0;
rom[76652] = 12'h  0;
rom[76653] = 12'h  0;
rom[76654] = 12'h  0;
rom[76655] = 12'h  0;
rom[76656] = 12'h  0;
rom[76657] = 12'h  0;
rom[76658] = 12'h  0;
rom[76659] = 12'h  0;
rom[76660] = 12'h  0;
rom[76661] = 12'h  0;
rom[76662] = 12'h  0;
rom[76663] = 12'h  0;
rom[76664] = 12'h  0;
rom[76665] = 12'h  0;
rom[76666] = 12'h  0;
rom[76667] = 12'h  0;
rom[76668] = 12'h  0;
rom[76669] = 12'h111;
rom[76670] = 12'h111;
rom[76671] = 12'h111;
rom[76672] = 12'h111;
rom[76673] = 12'h111;
rom[76674] = 12'h222;
rom[76675] = 12'h333;
rom[76676] = 12'h333;
rom[76677] = 12'h444;
rom[76678] = 12'h666;
rom[76679] = 12'h777;
rom[76680] = 12'h777;
rom[76681] = 12'h555;
rom[76682] = 12'h333;
rom[76683] = 12'h222;
rom[76684] = 12'h222;
rom[76685] = 12'h222;
rom[76686] = 12'h222;
rom[76687] = 12'h222;
rom[76688] = 12'h222;
rom[76689] = 12'h222;
rom[76690] = 12'h222;
rom[76691] = 12'h222;
rom[76692] = 12'h222;
rom[76693] = 12'h333;
rom[76694] = 12'h333;
rom[76695] = 12'h333;
rom[76696] = 12'h333;
rom[76697] = 12'h333;
rom[76698] = 12'h333;
rom[76699] = 12'h333;
rom[76700] = 12'h333;
rom[76701] = 12'h333;
rom[76702] = 12'h444;
rom[76703] = 12'h444;
rom[76704] = 12'h444;
rom[76705] = 12'h555;
rom[76706] = 12'h555;
rom[76707] = 12'h666;
rom[76708] = 12'h666;
rom[76709] = 12'h777;
rom[76710] = 12'h777;
rom[76711] = 12'h777;
rom[76712] = 12'h888;
rom[76713] = 12'h999;
rom[76714] = 12'haaa;
rom[76715] = 12'hbbb;
rom[76716] = 12'hccc;
rom[76717] = 12'hccc;
rom[76718] = 12'hddd;
rom[76719] = 12'heee;
rom[76720] = 12'hfff;
rom[76721] = 12'hfff;
rom[76722] = 12'hfff;
rom[76723] = 12'hfff;
rom[76724] = 12'hfff;
rom[76725] = 12'hfff;
rom[76726] = 12'hfff;
rom[76727] = 12'hfff;
rom[76728] = 12'heee;
rom[76729] = 12'hccc;
rom[76730] = 12'hbbb;
rom[76731] = 12'haaa;
rom[76732] = 12'haaa;
rom[76733] = 12'haaa;
rom[76734] = 12'h999;
rom[76735] = 12'h999;
rom[76736] = 12'h888;
rom[76737] = 12'h777;
rom[76738] = 12'h777;
rom[76739] = 12'h777;
rom[76740] = 12'h777;
rom[76741] = 12'h777;
rom[76742] = 12'h777;
rom[76743] = 12'h666;
rom[76744] = 12'h666;
rom[76745] = 12'h666;
rom[76746] = 12'h666;
rom[76747] = 12'h555;
rom[76748] = 12'h555;
rom[76749] = 12'h555;
rom[76750] = 12'h555;
rom[76751] = 12'h555;
rom[76752] = 12'h555;
rom[76753] = 12'h555;
rom[76754] = 12'h555;
rom[76755] = 12'h555;
rom[76756] = 12'h555;
rom[76757] = 12'h555;
rom[76758] = 12'h555;
rom[76759] = 12'h444;
rom[76760] = 12'h444;
rom[76761] = 12'h444;
rom[76762] = 12'h444;
rom[76763] = 12'h444;
rom[76764] = 12'h444;
rom[76765] = 12'h444;
rom[76766] = 12'h444;
rom[76767] = 12'h444;
rom[76768] = 12'h444;
rom[76769] = 12'h444;
rom[76770] = 12'h444;
rom[76771] = 12'h444;
rom[76772] = 12'h444;
rom[76773] = 12'h444;
rom[76774] = 12'h444;
rom[76775] = 12'h444;
rom[76776] = 12'h333;
rom[76777] = 12'h333;
rom[76778] = 12'h333;
rom[76779] = 12'h333;
rom[76780] = 12'h333;
rom[76781] = 12'h333;
rom[76782] = 12'h333;
rom[76783] = 12'h333;
rom[76784] = 12'h333;
rom[76785] = 12'h333;
rom[76786] = 12'h333;
rom[76787] = 12'h333;
rom[76788] = 12'h333;
rom[76789] = 12'h333;
rom[76790] = 12'h333;
rom[76791] = 12'h444;
rom[76792] = 12'h444;
rom[76793] = 12'h333;
rom[76794] = 12'h444;
rom[76795] = 12'h444;
rom[76796] = 12'h444;
rom[76797] = 12'h444;
rom[76798] = 12'h444;
rom[76799] = 12'h444;
rom[76800] = 12'hfff;
rom[76801] = 12'hfff;
rom[76802] = 12'hfff;
rom[76803] = 12'hfff;
rom[76804] = 12'hfff;
rom[76805] = 12'hfff;
rom[76806] = 12'hfff;
rom[76807] = 12'hfff;
rom[76808] = 12'hfff;
rom[76809] = 12'hfff;
rom[76810] = 12'hfff;
rom[76811] = 12'hfff;
rom[76812] = 12'hfff;
rom[76813] = 12'hfff;
rom[76814] = 12'hfff;
rom[76815] = 12'hfff;
rom[76816] = 12'hfff;
rom[76817] = 12'hfff;
rom[76818] = 12'hfff;
rom[76819] = 12'hfff;
rom[76820] = 12'hfff;
rom[76821] = 12'hfff;
rom[76822] = 12'hfff;
rom[76823] = 12'hfff;
rom[76824] = 12'hfff;
rom[76825] = 12'hfff;
rom[76826] = 12'hfff;
rom[76827] = 12'hfff;
rom[76828] = 12'hfff;
rom[76829] = 12'hfff;
rom[76830] = 12'hfff;
rom[76831] = 12'hfff;
rom[76832] = 12'hfff;
rom[76833] = 12'hfff;
rom[76834] = 12'hfff;
rom[76835] = 12'hfff;
rom[76836] = 12'hfff;
rom[76837] = 12'hfff;
rom[76838] = 12'hfff;
rom[76839] = 12'hfff;
rom[76840] = 12'hfff;
rom[76841] = 12'hfff;
rom[76842] = 12'hfff;
rom[76843] = 12'hfff;
rom[76844] = 12'hfff;
rom[76845] = 12'hfff;
rom[76846] = 12'hfff;
rom[76847] = 12'hfff;
rom[76848] = 12'hfff;
rom[76849] = 12'hfff;
rom[76850] = 12'hfff;
rom[76851] = 12'hfff;
rom[76852] = 12'hfff;
rom[76853] = 12'hfff;
rom[76854] = 12'hfff;
rom[76855] = 12'hfff;
rom[76856] = 12'hfff;
rom[76857] = 12'hfff;
rom[76858] = 12'hfff;
rom[76859] = 12'hfff;
rom[76860] = 12'hfff;
rom[76861] = 12'hfff;
rom[76862] = 12'hfff;
rom[76863] = 12'hfff;
rom[76864] = 12'hfff;
rom[76865] = 12'hfff;
rom[76866] = 12'hfff;
rom[76867] = 12'hfff;
rom[76868] = 12'hfff;
rom[76869] = 12'hfff;
rom[76870] = 12'hfff;
rom[76871] = 12'hfff;
rom[76872] = 12'hfff;
rom[76873] = 12'hfff;
rom[76874] = 12'hfff;
rom[76875] = 12'hfff;
rom[76876] = 12'hfff;
rom[76877] = 12'hfff;
rom[76878] = 12'hfff;
rom[76879] = 12'hfff;
rom[76880] = 12'hfff;
rom[76881] = 12'hfff;
rom[76882] = 12'hfff;
rom[76883] = 12'hfff;
rom[76884] = 12'hfff;
rom[76885] = 12'hfff;
rom[76886] = 12'hfff;
rom[76887] = 12'hfff;
rom[76888] = 12'hfff;
rom[76889] = 12'hfff;
rom[76890] = 12'hfff;
rom[76891] = 12'hfff;
rom[76892] = 12'hfff;
rom[76893] = 12'hfff;
rom[76894] = 12'hfff;
rom[76895] = 12'hfff;
rom[76896] = 12'hfff;
rom[76897] = 12'hfff;
rom[76898] = 12'hfff;
rom[76899] = 12'hfff;
rom[76900] = 12'hfff;
rom[76901] = 12'hfff;
rom[76902] = 12'hfff;
rom[76903] = 12'hfff;
rom[76904] = 12'hfff;
rom[76905] = 12'hfff;
rom[76906] = 12'hfff;
rom[76907] = 12'hfff;
rom[76908] = 12'hfff;
rom[76909] = 12'hfff;
rom[76910] = 12'hfff;
rom[76911] = 12'hfff;
rom[76912] = 12'hfff;
rom[76913] = 12'hfff;
rom[76914] = 12'heee;
rom[76915] = 12'heee;
rom[76916] = 12'hddd;
rom[76917] = 12'hddd;
rom[76918] = 12'hccc;
rom[76919] = 12'hccc;
rom[76920] = 12'hbbb;
rom[76921] = 12'hbbb;
rom[76922] = 12'hbbb;
rom[76923] = 12'haaa;
rom[76924] = 12'haaa;
rom[76925] = 12'haaa;
rom[76926] = 12'h999;
rom[76927] = 12'h999;
rom[76928] = 12'h888;
rom[76929] = 12'h777;
rom[76930] = 12'h777;
rom[76931] = 12'h777;
rom[76932] = 12'h777;
rom[76933] = 12'h777;
rom[76934] = 12'h777;
rom[76935] = 12'h777;
rom[76936] = 12'h777;
rom[76937] = 12'h777;
rom[76938] = 12'h777;
rom[76939] = 12'h777;
rom[76940] = 12'h777;
rom[76941] = 12'h777;
rom[76942] = 12'h777;
rom[76943] = 12'h777;
rom[76944] = 12'h777;
rom[76945] = 12'h777;
rom[76946] = 12'h777;
rom[76947] = 12'h777;
rom[76948] = 12'h777;
rom[76949] = 12'h777;
rom[76950] = 12'h777;
rom[76951] = 12'h777;
rom[76952] = 12'h777;
rom[76953] = 12'h777;
rom[76954] = 12'h777;
rom[76955] = 12'h777;
rom[76956] = 12'h666;
rom[76957] = 12'h666;
rom[76958] = 12'h666;
rom[76959] = 12'h666;
rom[76960] = 12'h666;
rom[76961] = 12'h666;
rom[76962] = 12'h666;
rom[76963] = 12'h666;
rom[76964] = 12'h666;
rom[76965] = 12'h666;
rom[76966] = 12'h666;
rom[76967] = 12'h666;
rom[76968] = 12'h666;
rom[76969] = 12'h666;
rom[76970] = 12'h666;
rom[76971] = 12'h666;
rom[76972] = 12'h666;
rom[76973] = 12'h666;
rom[76974] = 12'h666;
rom[76975] = 12'h666;
rom[76976] = 12'h555;
rom[76977] = 12'h555;
rom[76978] = 12'h555;
rom[76979] = 12'h444;
rom[76980] = 12'h444;
rom[76981] = 12'h444;
rom[76982] = 12'h555;
rom[76983] = 12'h555;
rom[76984] = 12'h555;
rom[76985] = 12'h555;
rom[76986] = 12'h555;
rom[76987] = 12'h666;
rom[76988] = 12'h666;
rom[76989] = 12'h666;
rom[76990] = 12'h666;
rom[76991] = 12'h555;
rom[76992] = 12'h555;
rom[76993] = 12'h666;
rom[76994] = 12'h666;
rom[76995] = 12'h777;
rom[76996] = 12'h777;
rom[76997] = 12'h666;
rom[76998] = 12'h666;
rom[76999] = 12'h666;
rom[77000] = 12'h777;
rom[77001] = 12'h777;
rom[77002] = 12'h777;
rom[77003] = 12'h777;
rom[77004] = 12'h555;
rom[77005] = 12'h444;
rom[77006] = 12'h444;
rom[77007] = 12'h444;
rom[77008] = 12'h444;
rom[77009] = 12'h333;
rom[77010] = 12'h333;
rom[77011] = 12'h222;
rom[77012] = 12'h333;
rom[77013] = 12'h333;
rom[77014] = 12'h222;
rom[77015] = 12'h222;
rom[77016] = 12'h222;
rom[77017] = 12'h222;
rom[77018] = 12'h222;
rom[77019] = 12'h222;
rom[77020] = 12'h222;
rom[77021] = 12'h222;
rom[77022] = 12'h222;
rom[77023] = 12'h222;
rom[77024] = 12'h222;
rom[77025] = 12'h222;
rom[77026] = 12'h222;
rom[77027] = 12'h222;
rom[77028] = 12'h222;
rom[77029] = 12'h111;
rom[77030] = 12'h111;
rom[77031] = 12'h111;
rom[77032] = 12'h111;
rom[77033] = 12'h111;
rom[77034] = 12'h111;
rom[77035] = 12'h  0;
rom[77036] = 12'h  0;
rom[77037] = 12'h  0;
rom[77038] = 12'h  0;
rom[77039] = 12'h  0;
rom[77040] = 12'h  0;
rom[77041] = 12'h  0;
rom[77042] = 12'h  0;
rom[77043] = 12'h  0;
rom[77044] = 12'h  0;
rom[77045] = 12'h  0;
rom[77046] = 12'h  0;
rom[77047] = 12'h  0;
rom[77048] = 12'h  0;
rom[77049] = 12'h  0;
rom[77050] = 12'h  0;
rom[77051] = 12'h  0;
rom[77052] = 12'h  0;
rom[77053] = 12'h  0;
rom[77054] = 12'h  0;
rom[77055] = 12'h  0;
rom[77056] = 12'h  0;
rom[77057] = 12'h  0;
rom[77058] = 12'h  0;
rom[77059] = 12'h  0;
rom[77060] = 12'h  0;
rom[77061] = 12'h  0;
rom[77062] = 12'h  0;
rom[77063] = 12'h  0;
rom[77064] = 12'h  0;
rom[77065] = 12'h  0;
rom[77066] = 12'h  0;
rom[77067] = 12'h  0;
rom[77068] = 12'h  0;
rom[77069] = 12'h  0;
rom[77070] = 12'h111;
rom[77071] = 12'h111;
rom[77072] = 12'h111;
rom[77073] = 12'h222;
rom[77074] = 12'h222;
rom[77075] = 12'h333;
rom[77076] = 12'h333;
rom[77077] = 12'h444;
rom[77078] = 12'h666;
rom[77079] = 12'h888;
rom[77080] = 12'h888;
rom[77081] = 12'h666;
rom[77082] = 12'h333;
rom[77083] = 12'h333;
rom[77084] = 12'h333;
rom[77085] = 12'h222;
rom[77086] = 12'h222;
rom[77087] = 12'h222;
rom[77088] = 12'h333;
rom[77089] = 12'h333;
rom[77090] = 12'h333;
rom[77091] = 12'h333;
rom[77092] = 12'h333;
rom[77093] = 12'h333;
rom[77094] = 12'h333;
rom[77095] = 12'h333;
rom[77096] = 12'h333;
rom[77097] = 12'h333;
rom[77098] = 12'h333;
rom[77099] = 12'h333;
rom[77100] = 12'h333;
rom[77101] = 12'h333;
rom[77102] = 12'h444;
rom[77103] = 12'h444;
rom[77104] = 12'h444;
rom[77105] = 12'h555;
rom[77106] = 12'h555;
rom[77107] = 12'h666;
rom[77108] = 12'h666;
rom[77109] = 12'h777;
rom[77110] = 12'h777;
rom[77111] = 12'h777;
rom[77112] = 12'h888;
rom[77113] = 12'h999;
rom[77114] = 12'haaa;
rom[77115] = 12'hbbb;
rom[77116] = 12'hccc;
rom[77117] = 12'hddd;
rom[77118] = 12'heee;
rom[77119] = 12'hfff;
rom[77120] = 12'hfff;
rom[77121] = 12'hfff;
rom[77122] = 12'hfff;
rom[77123] = 12'hfff;
rom[77124] = 12'hfff;
rom[77125] = 12'hfff;
rom[77126] = 12'heee;
rom[77127] = 12'hddd;
rom[77128] = 12'hccc;
rom[77129] = 12'hbbb;
rom[77130] = 12'haaa;
rom[77131] = 12'haaa;
rom[77132] = 12'h999;
rom[77133] = 12'h999;
rom[77134] = 12'h888;
rom[77135] = 12'h888;
rom[77136] = 12'h777;
rom[77137] = 12'h777;
rom[77138] = 12'h777;
rom[77139] = 12'h777;
rom[77140] = 12'h777;
rom[77141] = 12'h777;
rom[77142] = 12'h777;
rom[77143] = 12'h666;
rom[77144] = 12'h666;
rom[77145] = 12'h666;
rom[77146] = 12'h555;
rom[77147] = 12'h555;
rom[77148] = 12'h555;
rom[77149] = 12'h555;
rom[77150] = 12'h444;
rom[77151] = 12'h444;
rom[77152] = 12'h555;
rom[77153] = 12'h555;
rom[77154] = 12'h555;
rom[77155] = 12'h555;
rom[77156] = 12'h555;
rom[77157] = 12'h555;
rom[77158] = 12'h555;
rom[77159] = 12'h555;
rom[77160] = 12'h555;
rom[77161] = 12'h444;
rom[77162] = 12'h444;
rom[77163] = 12'h444;
rom[77164] = 12'h444;
rom[77165] = 12'h444;
rom[77166] = 12'h444;
rom[77167] = 12'h444;
rom[77168] = 12'h444;
rom[77169] = 12'h444;
rom[77170] = 12'h333;
rom[77171] = 12'h333;
rom[77172] = 12'h333;
rom[77173] = 12'h333;
rom[77174] = 12'h333;
rom[77175] = 12'h333;
rom[77176] = 12'h333;
rom[77177] = 12'h333;
rom[77178] = 12'h333;
rom[77179] = 12'h333;
rom[77180] = 12'h333;
rom[77181] = 12'h333;
rom[77182] = 12'h333;
rom[77183] = 12'h333;
rom[77184] = 12'h333;
rom[77185] = 12'h333;
rom[77186] = 12'h333;
rom[77187] = 12'h333;
rom[77188] = 12'h333;
rom[77189] = 12'h333;
rom[77190] = 12'h333;
rom[77191] = 12'h333;
rom[77192] = 12'h333;
rom[77193] = 12'h333;
rom[77194] = 12'h333;
rom[77195] = 12'h444;
rom[77196] = 12'h444;
rom[77197] = 12'h444;
rom[77198] = 12'h444;
rom[77199] = 12'h444;
rom[77200] = 12'hfff;
rom[77201] = 12'hfff;
rom[77202] = 12'hfff;
rom[77203] = 12'hfff;
rom[77204] = 12'hfff;
rom[77205] = 12'hfff;
rom[77206] = 12'hfff;
rom[77207] = 12'hfff;
rom[77208] = 12'hfff;
rom[77209] = 12'hfff;
rom[77210] = 12'hfff;
rom[77211] = 12'hfff;
rom[77212] = 12'hfff;
rom[77213] = 12'hfff;
rom[77214] = 12'hfff;
rom[77215] = 12'hfff;
rom[77216] = 12'hfff;
rom[77217] = 12'hfff;
rom[77218] = 12'hfff;
rom[77219] = 12'hfff;
rom[77220] = 12'hfff;
rom[77221] = 12'hfff;
rom[77222] = 12'hfff;
rom[77223] = 12'hfff;
rom[77224] = 12'hfff;
rom[77225] = 12'hfff;
rom[77226] = 12'hfff;
rom[77227] = 12'hfff;
rom[77228] = 12'hfff;
rom[77229] = 12'hfff;
rom[77230] = 12'hfff;
rom[77231] = 12'hfff;
rom[77232] = 12'hfff;
rom[77233] = 12'hfff;
rom[77234] = 12'hfff;
rom[77235] = 12'hfff;
rom[77236] = 12'hfff;
rom[77237] = 12'hfff;
rom[77238] = 12'hfff;
rom[77239] = 12'hfff;
rom[77240] = 12'hfff;
rom[77241] = 12'hfff;
rom[77242] = 12'hfff;
rom[77243] = 12'hfff;
rom[77244] = 12'hfff;
rom[77245] = 12'hfff;
rom[77246] = 12'hfff;
rom[77247] = 12'hfff;
rom[77248] = 12'hfff;
rom[77249] = 12'hfff;
rom[77250] = 12'hfff;
rom[77251] = 12'hfff;
rom[77252] = 12'hfff;
rom[77253] = 12'hfff;
rom[77254] = 12'hfff;
rom[77255] = 12'hfff;
rom[77256] = 12'hfff;
rom[77257] = 12'hfff;
rom[77258] = 12'hfff;
rom[77259] = 12'hfff;
rom[77260] = 12'hfff;
rom[77261] = 12'hfff;
rom[77262] = 12'hfff;
rom[77263] = 12'hfff;
rom[77264] = 12'hfff;
rom[77265] = 12'hfff;
rom[77266] = 12'hfff;
rom[77267] = 12'hfff;
rom[77268] = 12'hfff;
rom[77269] = 12'hfff;
rom[77270] = 12'hfff;
rom[77271] = 12'hfff;
rom[77272] = 12'hfff;
rom[77273] = 12'hfff;
rom[77274] = 12'hfff;
rom[77275] = 12'hfff;
rom[77276] = 12'hfff;
rom[77277] = 12'hfff;
rom[77278] = 12'hfff;
rom[77279] = 12'hfff;
rom[77280] = 12'hfff;
rom[77281] = 12'hfff;
rom[77282] = 12'hfff;
rom[77283] = 12'hfff;
rom[77284] = 12'hfff;
rom[77285] = 12'hfff;
rom[77286] = 12'hfff;
rom[77287] = 12'hfff;
rom[77288] = 12'hfff;
rom[77289] = 12'hfff;
rom[77290] = 12'hfff;
rom[77291] = 12'hfff;
rom[77292] = 12'hfff;
rom[77293] = 12'hfff;
rom[77294] = 12'hfff;
rom[77295] = 12'hfff;
rom[77296] = 12'hfff;
rom[77297] = 12'hfff;
rom[77298] = 12'hfff;
rom[77299] = 12'hfff;
rom[77300] = 12'hfff;
rom[77301] = 12'hfff;
rom[77302] = 12'hfff;
rom[77303] = 12'hfff;
rom[77304] = 12'hfff;
rom[77305] = 12'hfff;
rom[77306] = 12'hfff;
rom[77307] = 12'hfff;
rom[77308] = 12'hfff;
rom[77309] = 12'hfff;
rom[77310] = 12'hfff;
rom[77311] = 12'hfff;
rom[77312] = 12'hfff;
rom[77313] = 12'hfff;
rom[77314] = 12'hfff;
rom[77315] = 12'heee;
rom[77316] = 12'heee;
rom[77317] = 12'hddd;
rom[77318] = 12'hccc;
rom[77319] = 12'hccc;
rom[77320] = 12'hccc;
rom[77321] = 12'hbbb;
rom[77322] = 12'hbbb;
rom[77323] = 12'hbbb;
rom[77324] = 12'haaa;
rom[77325] = 12'haaa;
rom[77326] = 12'h999;
rom[77327] = 12'h999;
rom[77328] = 12'h999;
rom[77329] = 12'h888;
rom[77330] = 12'h888;
rom[77331] = 12'h777;
rom[77332] = 12'h777;
rom[77333] = 12'h777;
rom[77334] = 12'h777;
rom[77335] = 12'h777;
rom[77336] = 12'h777;
rom[77337] = 12'h777;
rom[77338] = 12'h777;
rom[77339] = 12'h777;
rom[77340] = 12'h777;
rom[77341] = 12'h777;
rom[77342] = 12'h777;
rom[77343] = 12'h777;
rom[77344] = 12'h777;
rom[77345] = 12'h777;
rom[77346] = 12'h777;
rom[77347] = 12'h777;
rom[77348] = 12'h777;
rom[77349] = 12'h777;
rom[77350] = 12'h777;
rom[77351] = 12'h777;
rom[77352] = 12'h777;
rom[77353] = 12'h777;
rom[77354] = 12'h666;
rom[77355] = 12'h666;
rom[77356] = 12'h666;
rom[77357] = 12'h666;
rom[77358] = 12'h666;
rom[77359] = 12'h666;
rom[77360] = 12'h666;
rom[77361] = 12'h666;
rom[77362] = 12'h666;
rom[77363] = 12'h666;
rom[77364] = 12'h666;
rom[77365] = 12'h666;
rom[77366] = 12'h666;
rom[77367] = 12'h666;
rom[77368] = 12'h666;
rom[77369] = 12'h666;
rom[77370] = 12'h666;
rom[77371] = 12'h666;
rom[77372] = 12'h666;
rom[77373] = 12'h666;
rom[77374] = 12'h666;
rom[77375] = 12'h666;
rom[77376] = 12'h555;
rom[77377] = 12'h555;
rom[77378] = 12'h555;
rom[77379] = 12'h555;
rom[77380] = 12'h555;
rom[77381] = 12'h555;
rom[77382] = 12'h555;
rom[77383] = 12'h555;
rom[77384] = 12'h555;
rom[77385] = 12'h555;
rom[77386] = 12'h555;
rom[77387] = 12'h555;
rom[77388] = 12'h555;
rom[77389] = 12'h555;
rom[77390] = 12'h555;
rom[77391] = 12'h555;
rom[77392] = 12'h555;
rom[77393] = 12'h666;
rom[77394] = 12'h666;
rom[77395] = 12'h777;
rom[77396] = 12'h777;
rom[77397] = 12'h777;
rom[77398] = 12'h777;
rom[77399] = 12'h777;
rom[77400] = 12'h777;
rom[77401] = 12'h777;
rom[77402] = 12'h888;
rom[77403] = 12'h777;
rom[77404] = 12'h666;
rom[77405] = 12'h555;
rom[77406] = 12'h444;
rom[77407] = 12'h444;
rom[77408] = 12'h444;
rom[77409] = 12'h444;
rom[77410] = 12'h333;
rom[77411] = 12'h333;
rom[77412] = 12'h333;
rom[77413] = 12'h333;
rom[77414] = 12'h333;
rom[77415] = 12'h222;
rom[77416] = 12'h222;
rom[77417] = 12'h222;
rom[77418] = 12'h222;
rom[77419] = 12'h222;
rom[77420] = 12'h222;
rom[77421] = 12'h222;
rom[77422] = 12'h222;
rom[77423] = 12'h222;
rom[77424] = 12'h222;
rom[77425] = 12'h222;
rom[77426] = 12'h222;
rom[77427] = 12'h222;
rom[77428] = 12'h222;
rom[77429] = 12'h222;
rom[77430] = 12'h111;
rom[77431] = 12'h111;
rom[77432] = 12'h111;
rom[77433] = 12'h111;
rom[77434] = 12'h111;
rom[77435] = 12'h  0;
rom[77436] = 12'h  0;
rom[77437] = 12'h  0;
rom[77438] = 12'h  0;
rom[77439] = 12'h  0;
rom[77440] = 12'h  0;
rom[77441] = 12'h  0;
rom[77442] = 12'h  0;
rom[77443] = 12'h  0;
rom[77444] = 12'h  0;
rom[77445] = 12'h  0;
rom[77446] = 12'h  0;
rom[77447] = 12'h  0;
rom[77448] = 12'h  0;
rom[77449] = 12'h  0;
rom[77450] = 12'h  0;
rom[77451] = 12'h  0;
rom[77452] = 12'h  0;
rom[77453] = 12'h  0;
rom[77454] = 12'h  0;
rom[77455] = 12'h  0;
rom[77456] = 12'h  0;
rom[77457] = 12'h  0;
rom[77458] = 12'h  0;
rom[77459] = 12'h  0;
rom[77460] = 12'h  0;
rom[77461] = 12'h  0;
rom[77462] = 12'h  0;
rom[77463] = 12'h  0;
rom[77464] = 12'h  0;
rom[77465] = 12'h  0;
rom[77466] = 12'h  0;
rom[77467] = 12'h  0;
rom[77468] = 12'h  0;
rom[77469] = 12'h  0;
rom[77470] = 12'h111;
rom[77471] = 12'h111;
rom[77472] = 12'h111;
rom[77473] = 12'h222;
rom[77474] = 12'h222;
rom[77475] = 12'h333;
rom[77476] = 12'h333;
rom[77477] = 12'h444;
rom[77478] = 12'h666;
rom[77479] = 12'h888;
rom[77480] = 12'h888;
rom[77481] = 12'h666;
rom[77482] = 12'h444;
rom[77483] = 12'h333;
rom[77484] = 12'h333;
rom[77485] = 12'h222;
rom[77486] = 12'h222;
rom[77487] = 12'h333;
rom[77488] = 12'h333;
rom[77489] = 12'h333;
rom[77490] = 12'h333;
rom[77491] = 12'h333;
rom[77492] = 12'h333;
rom[77493] = 12'h333;
rom[77494] = 12'h333;
rom[77495] = 12'h333;
rom[77496] = 12'h333;
rom[77497] = 12'h333;
rom[77498] = 12'h333;
rom[77499] = 12'h444;
rom[77500] = 12'h444;
rom[77501] = 12'h444;
rom[77502] = 12'h444;
rom[77503] = 12'h444;
rom[77504] = 12'h555;
rom[77505] = 12'h555;
rom[77506] = 12'h666;
rom[77507] = 12'h666;
rom[77508] = 12'h666;
rom[77509] = 12'h777;
rom[77510] = 12'h888;
rom[77511] = 12'h888;
rom[77512] = 12'h999;
rom[77513] = 12'haaa;
rom[77514] = 12'hbbb;
rom[77515] = 12'hccc;
rom[77516] = 12'hddd;
rom[77517] = 12'heee;
rom[77518] = 12'hfff;
rom[77519] = 12'hfff;
rom[77520] = 12'hfff;
rom[77521] = 12'hfff;
rom[77522] = 12'hfff;
rom[77523] = 12'hfff;
rom[77524] = 12'hfff;
rom[77525] = 12'heee;
rom[77526] = 12'hddd;
rom[77527] = 12'hccc;
rom[77528] = 12'hbbb;
rom[77529] = 12'haaa;
rom[77530] = 12'haaa;
rom[77531] = 12'h999;
rom[77532] = 12'h999;
rom[77533] = 12'h888;
rom[77534] = 12'h888;
rom[77535] = 12'h777;
rom[77536] = 12'h777;
rom[77537] = 12'h777;
rom[77538] = 12'h777;
rom[77539] = 12'h777;
rom[77540] = 12'h666;
rom[77541] = 12'h666;
rom[77542] = 12'h666;
rom[77543] = 12'h666;
rom[77544] = 12'h666;
rom[77545] = 12'h555;
rom[77546] = 12'h555;
rom[77547] = 12'h555;
rom[77548] = 12'h555;
rom[77549] = 12'h555;
rom[77550] = 12'h444;
rom[77551] = 12'h444;
rom[77552] = 12'h444;
rom[77553] = 12'h444;
rom[77554] = 12'h555;
rom[77555] = 12'h555;
rom[77556] = 12'h555;
rom[77557] = 12'h555;
rom[77558] = 12'h555;
rom[77559] = 12'h555;
rom[77560] = 12'h444;
rom[77561] = 12'h444;
rom[77562] = 12'h444;
rom[77563] = 12'h444;
rom[77564] = 12'h444;
rom[77565] = 12'h444;
rom[77566] = 12'h444;
rom[77567] = 12'h444;
rom[77568] = 12'h444;
rom[77569] = 12'h444;
rom[77570] = 12'h333;
rom[77571] = 12'h333;
rom[77572] = 12'h333;
rom[77573] = 12'h333;
rom[77574] = 12'h333;
rom[77575] = 12'h333;
rom[77576] = 12'h333;
rom[77577] = 12'h333;
rom[77578] = 12'h333;
rom[77579] = 12'h333;
rom[77580] = 12'h333;
rom[77581] = 12'h333;
rom[77582] = 12'h333;
rom[77583] = 12'h333;
rom[77584] = 12'h333;
rom[77585] = 12'h333;
rom[77586] = 12'h333;
rom[77587] = 12'h333;
rom[77588] = 12'h333;
rom[77589] = 12'h333;
rom[77590] = 12'h333;
rom[77591] = 12'h333;
rom[77592] = 12'h333;
rom[77593] = 12'h333;
rom[77594] = 12'h333;
rom[77595] = 12'h333;
rom[77596] = 12'h444;
rom[77597] = 12'h444;
rom[77598] = 12'h444;
rom[77599] = 12'h444;
rom[77600] = 12'hfff;
rom[77601] = 12'hfff;
rom[77602] = 12'hfff;
rom[77603] = 12'hfff;
rom[77604] = 12'hfff;
rom[77605] = 12'hfff;
rom[77606] = 12'hfff;
rom[77607] = 12'hfff;
rom[77608] = 12'hfff;
rom[77609] = 12'hfff;
rom[77610] = 12'hfff;
rom[77611] = 12'hfff;
rom[77612] = 12'hfff;
rom[77613] = 12'hfff;
rom[77614] = 12'hfff;
rom[77615] = 12'hfff;
rom[77616] = 12'hfff;
rom[77617] = 12'hfff;
rom[77618] = 12'hfff;
rom[77619] = 12'hfff;
rom[77620] = 12'hfff;
rom[77621] = 12'hfff;
rom[77622] = 12'hfff;
rom[77623] = 12'hfff;
rom[77624] = 12'hfff;
rom[77625] = 12'hfff;
rom[77626] = 12'hfff;
rom[77627] = 12'hfff;
rom[77628] = 12'hfff;
rom[77629] = 12'hfff;
rom[77630] = 12'hfff;
rom[77631] = 12'hfff;
rom[77632] = 12'hfff;
rom[77633] = 12'hfff;
rom[77634] = 12'hfff;
rom[77635] = 12'hfff;
rom[77636] = 12'hfff;
rom[77637] = 12'hfff;
rom[77638] = 12'hfff;
rom[77639] = 12'hfff;
rom[77640] = 12'hfff;
rom[77641] = 12'hfff;
rom[77642] = 12'hfff;
rom[77643] = 12'hfff;
rom[77644] = 12'hfff;
rom[77645] = 12'hfff;
rom[77646] = 12'hfff;
rom[77647] = 12'hfff;
rom[77648] = 12'hfff;
rom[77649] = 12'hfff;
rom[77650] = 12'hfff;
rom[77651] = 12'hfff;
rom[77652] = 12'hfff;
rom[77653] = 12'hfff;
rom[77654] = 12'hfff;
rom[77655] = 12'hfff;
rom[77656] = 12'hfff;
rom[77657] = 12'hfff;
rom[77658] = 12'hfff;
rom[77659] = 12'hfff;
rom[77660] = 12'hfff;
rom[77661] = 12'hfff;
rom[77662] = 12'hfff;
rom[77663] = 12'hfff;
rom[77664] = 12'hfff;
rom[77665] = 12'hfff;
rom[77666] = 12'hfff;
rom[77667] = 12'hfff;
rom[77668] = 12'hfff;
rom[77669] = 12'hfff;
rom[77670] = 12'hfff;
rom[77671] = 12'hfff;
rom[77672] = 12'hfff;
rom[77673] = 12'hfff;
rom[77674] = 12'hfff;
rom[77675] = 12'hfff;
rom[77676] = 12'hfff;
rom[77677] = 12'hfff;
rom[77678] = 12'hfff;
rom[77679] = 12'hfff;
rom[77680] = 12'hfff;
rom[77681] = 12'hfff;
rom[77682] = 12'hfff;
rom[77683] = 12'hfff;
rom[77684] = 12'hfff;
rom[77685] = 12'hfff;
rom[77686] = 12'hfff;
rom[77687] = 12'hfff;
rom[77688] = 12'hfff;
rom[77689] = 12'hfff;
rom[77690] = 12'hfff;
rom[77691] = 12'hfff;
rom[77692] = 12'hfff;
rom[77693] = 12'hfff;
rom[77694] = 12'hfff;
rom[77695] = 12'hfff;
rom[77696] = 12'hfff;
rom[77697] = 12'hfff;
rom[77698] = 12'hfff;
rom[77699] = 12'hfff;
rom[77700] = 12'hfff;
rom[77701] = 12'hfff;
rom[77702] = 12'hfff;
rom[77703] = 12'hfff;
rom[77704] = 12'hfff;
rom[77705] = 12'hfff;
rom[77706] = 12'hfff;
rom[77707] = 12'hfff;
rom[77708] = 12'hfff;
rom[77709] = 12'hfff;
rom[77710] = 12'hfff;
rom[77711] = 12'hfff;
rom[77712] = 12'hfff;
rom[77713] = 12'hfff;
rom[77714] = 12'hfff;
rom[77715] = 12'hfff;
rom[77716] = 12'heee;
rom[77717] = 12'heee;
rom[77718] = 12'hddd;
rom[77719] = 12'hddd;
rom[77720] = 12'hccc;
rom[77721] = 12'hccc;
rom[77722] = 12'hbbb;
rom[77723] = 12'hbbb;
rom[77724] = 12'hbbb;
rom[77725] = 12'haaa;
rom[77726] = 12'haaa;
rom[77727] = 12'h999;
rom[77728] = 12'h999;
rom[77729] = 12'h999;
rom[77730] = 12'h888;
rom[77731] = 12'h888;
rom[77732] = 12'h777;
rom[77733] = 12'h777;
rom[77734] = 12'h777;
rom[77735] = 12'h777;
rom[77736] = 12'h777;
rom[77737] = 12'h777;
rom[77738] = 12'h777;
rom[77739] = 12'h777;
rom[77740] = 12'h777;
rom[77741] = 12'h888;
rom[77742] = 12'h888;
rom[77743] = 12'h888;
rom[77744] = 12'h888;
rom[77745] = 12'h888;
rom[77746] = 12'h888;
rom[77747] = 12'h888;
rom[77748] = 12'h888;
rom[77749] = 12'h777;
rom[77750] = 12'h777;
rom[77751] = 12'h777;
rom[77752] = 12'h777;
rom[77753] = 12'h666;
rom[77754] = 12'h666;
rom[77755] = 12'h666;
rom[77756] = 12'h666;
rom[77757] = 12'h666;
rom[77758] = 12'h666;
rom[77759] = 12'h666;
rom[77760] = 12'h666;
rom[77761] = 12'h666;
rom[77762] = 12'h666;
rom[77763] = 12'h666;
rom[77764] = 12'h666;
rom[77765] = 12'h666;
rom[77766] = 12'h555;
rom[77767] = 12'h555;
rom[77768] = 12'h555;
rom[77769] = 12'h555;
rom[77770] = 12'h555;
rom[77771] = 12'h555;
rom[77772] = 12'h555;
rom[77773] = 12'h555;
rom[77774] = 12'h555;
rom[77775] = 12'h555;
rom[77776] = 12'h555;
rom[77777] = 12'h555;
rom[77778] = 12'h555;
rom[77779] = 12'h555;
rom[77780] = 12'h555;
rom[77781] = 12'h555;
rom[77782] = 12'h555;
rom[77783] = 12'h555;
rom[77784] = 12'h555;
rom[77785] = 12'h444;
rom[77786] = 12'h444;
rom[77787] = 12'h444;
rom[77788] = 12'h444;
rom[77789] = 12'h555;
rom[77790] = 12'h555;
rom[77791] = 12'h555;
rom[77792] = 12'h666;
rom[77793] = 12'h666;
rom[77794] = 12'h666;
rom[77795] = 12'h777;
rom[77796] = 12'h777;
rom[77797] = 12'h777;
rom[77798] = 12'h777;
rom[77799] = 12'h777;
rom[77800] = 12'h777;
rom[77801] = 12'h888;
rom[77802] = 12'h888;
rom[77803] = 12'h777;
rom[77804] = 12'h777;
rom[77805] = 12'h666;
rom[77806] = 12'h555;
rom[77807] = 12'h555;
rom[77808] = 12'h444;
rom[77809] = 12'h444;
rom[77810] = 12'h444;
rom[77811] = 12'h333;
rom[77812] = 12'h333;
rom[77813] = 12'h333;
rom[77814] = 12'h333;
rom[77815] = 12'h333;
rom[77816] = 12'h333;
rom[77817] = 12'h333;
rom[77818] = 12'h222;
rom[77819] = 12'h222;
rom[77820] = 12'h222;
rom[77821] = 12'h222;
rom[77822] = 12'h222;
rom[77823] = 12'h222;
rom[77824] = 12'h222;
rom[77825] = 12'h222;
rom[77826] = 12'h222;
rom[77827] = 12'h222;
rom[77828] = 12'h222;
rom[77829] = 12'h222;
rom[77830] = 12'h111;
rom[77831] = 12'h111;
rom[77832] = 12'h111;
rom[77833] = 12'h111;
rom[77834] = 12'h111;
rom[77835] = 12'h  0;
rom[77836] = 12'h  0;
rom[77837] = 12'h  0;
rom[77838] = 12'h  0;
rom[77839] = 12'h  0;
rom[77840] = 12'h  0;
rom[77841] = 12'h  0;
rom[77842] = 12'h  0;
rom[77843] = 12'h  0;
rom[77844] = 12'h  0;
rom[77845] = 12'h  0;
rom[77846] = 12'h  0;
rom[77847] = 12'h  0;
rom[77848] = 12'h  0;
rom[77849] = 12'h  0;
rom[77850] = 12'h  0;
rom[77851] = 12'h  0;
rom[77852] = 12'h  0;
rom[77853] = 12'h  0;
rom[77854] = 12'h  0;
rom[77855] = 12'h  0;
rom[77856] = 12'h  0;
rom[77857] = 12'h  0;
rom[77858] = 12'h  0;
rom[77859] = 12'h  0;
rom[77860] = 12'h  0;
rom[77861] = 12'h  0;
rom[77862] = 12'h  0;
rom[77863] = 12'h  0;
rom[77864] = 12'h  0;
rom[77865] = 12'h  0;
rom[77866] = 12'h  0;
rom[77867] = 12'h  0;
rom[77868] = 12'h  0;
rom[77869] = 12'h  0;
rom[77870] = 12'h111;
rom[77871] = 12'h111;
rom[77872] = 12'h111;
rom[77873] = 12'h222;
rom[77874] = 12'h222;
rom[77875] = 12'h333;
rom[77876] = 12'h333;
rom[77877] = 12'h444;
rom[77878] = 12'h666;
rom[77879] = 12'h888;
rom[77880] = 12'h888;
rom[77881] = 12'h777;
rom[77882] = 12'h444;
rom[77883] = 12'h333;
rom[77884] = 12'h333;
rom[77885] = 12'h333;
rom[77886] = 12'h222;
rom[77887] = 12'h333;
rom[77888] = 12'h333;
rom[77889] = 12'h333;
rom[77890] = 12'h333;
rom[77891] = 12'h333;
rom[77892] = 12'h333;
rom[77893] = 12'h333;
rom[77894] = 12'h333;
rom[77895] = 12'h333;
rom[77896] = 12'h333;
rom[77897] = 12'h444;
rom[77898] = 12'h444;
rom[77899] = 12'h444;
rom[77900] = 12'h444;
rom[77901] = 12'h444;
rom[77902] = 12'h555;
rom[77903] = 12'h555;
rom[77904] = 12'h555;
rom[77905] = 12'h555;
rom[77906] = 12'h666;
rom[77907] = 12'h666;
rom[77908] = 12'h777;
rom[77909] = 12'h777;
rom[77910] = 12'h888;
rom[77911] = 12'h999;
rom[77912] = 12'h999;
rom[77913] = 12'haaa;
rom[77914] = 12'hbbb;
rom[77915] = 12'hccc;
rom[77916] = 12'hddd;
rom[77917] = 12'heee;
rom[77918] = 12'hfff;
rom[77919] = 12'hfff;
rom[77920] = 12'hfff;
rom[77921] = 12'hfff;
rom[77922] = 12'hfff;
rom[77923] = 12'heee;
rom[77924] = 12'hddd;
rom[77925] = 12'hddd;
rom[77926] = 12'hccc;
rom[77927] = 12'hbbb;
rom[77928] = 12'haaa;
rom[77929] = 12'haaa;
rom[77930] = 12'h999;
rom[77931] = 12'h999;
rom[77932] = 12'h888;
rom[77933] = 12'h888;
rom[77934] = 12'h777;
rom[77935] = 12'h777;
rom[77936] = 12'h666;
rom[77937] = 12'h666;
rom[77938] = 12'h666;
rom[77939] = 12'h666;
rom[77940] = 12'h666;
rom[77941] = 12'h666;
rom[77942] = 12'h555;
rom[77943] = 12'h555;
rom[77944] = 12'h555;
rom[77945] = 12'h555;
rom[77946] = 12'h555;
rom[77947] = 12'h555;
rom[77948] = 12'h555;
rom[77949] = 12'h444;
rom[77950] = 12'h444;
rom[77951] = 12'h444;
rom[77952] = 12'h444;
rom[77953] = 12'h444;
rom[77954] = 12'h444;
rom[77955] = 12'h444;
rom[77956] = 12'h444;
rom[77957] = 12'h444;
rom[77958] = 12'h444;
rom[77959] = 12'h444;
rom[77960] = 12'h444;
rom[77961] = 12'h444;
rom[77962] = 12'h444;
rom[77963] = 12'h444;
rom[77964] = 12'h444;
rom[77965] = 12'h444;
rom[77966] = 12'h444;
rom[77967] = 12'h444;
rom[77968] = 12'h444;
rom[77969] = 12'h333;
rom[77970] = 12'h333;
rom[77971] = 12'h333;
rom[77972] = 12'h333;
rom[77973] = 12'h333;
rom[77974] = 12'h333;
rom[77975] = 12'h333;
rom[77976] = 12'h333;
rom[77977] = 12'h333;
rom[77978] = 12'h333;
rom[77979] = 12'h333;
rom[77980] = 12'h333;
rom[77981] = 12'h333;
rom[77982] = 12'h333;
rom[77983] = 12'h333;
rom[77984] = 12'h333;
rom[77985] = 12'h333;
rom[77986] = 12'h333;
rom[77987] = 12'h333;
rom[77988] = 12'h333;
rom[77989] = 12'h333;
rom[77990] = 12'h333;
rom[77991] = 12'h333;
rom[77992] = 12'h333;
rom[77993] = 12'h333;
rom[77994] = 12'h333;
rom[77995] = 12'h333;
rom[77996] = 12'h333;
rom[77997] = 12'h333;
rom[77998] = 12'h444;
rom[77999] = 12'h444;
rom[78000] = 12'hfff;
rom[78001] = 12'hfff;
rom[78002] = 12'hfff;
rom[78003] = 12'hfff;
rom[78004] = 12'hfff;
rom[78005] = 12'hfff;
rom[78006] = 12'hfff;
rom[78007] = 12'hfff;
rom[78008] = 12'hfff;
rom[78009] = 12'hfff;
rom[78010] = 12'hfff;
rom[78011] = 12'hfff;
rom[78012] = 12'hfff;
rom[78013] = 12'hfff;
rom[78014] = 12'hfff;
rom[78015] = 12'hfff;
rom[78016] = 12'hfff;
rom[78017] = 12'hfff;
rom[78018] = 12'hfff;
rom[78019] = 12'hfff;
rom[78020] = 12'hfff;
rom[78021] = 12'hfff;
rom[78022] = 12'hfff;
rom[78023] = 12'hfff;
rom[78024] = 12'hfff;
rom[78025] = 12'hfff;
rom[78026] = 12'hfff;
rom[78027] = 12'hfff;
rom[78028] = 12'hfff;
rom[78029] = 12'hfff;
rom[78030] = 12'hfff;
rom[78031] = 12'hfff;
rom[78032] = 12'hfff;
rom[78033] = 12'hfff;
rom[78034] = 12'hfff;
rom[78035] = 12'hfff;
rom[78036] = 12'hfff;
rom[78037] = 12'hfff;
rom[78038] = 12'hfff;
rom[78039] = 12'hfff;
rom[78040] = 12'hfff;
rom[78041] = 12'hfff;
rom[78042] = 12'hfff;
rom[78043] = 12'hfff;
rom[78044] = 12'hfff;
rom[78045] = 12'hfff;
rom[78046] = 12'hfff;
rom[78047] = 12'hfff;
rom[78048] = 12'hfff;
rom[78049] = 12'hfff;
rom[78050] = 12'hfff;
rom[78051] = 12'hfff;
rom[78052] = 12'hfff;
rom[78053] = 12'hfff;
rom[78054] = 12'hfff;
rom[78055] = 12'hfff;
rom[78056] = 12'hfff;
rom[78057] = 12'hfff;
rom[78058] = 12'hfff;
rom[78059] = 12'hfff;
rom[78060] = 12'hfff;
rom[78061] = 12'hfff;
rom[78062] = 12'hfff;
rom[78063] = 12'hfff;
rom[78064] = 12'hfff;
rom[78065] = 12'hfff;
rom[78066] = 12'hfff;
rom[78067] = 12'hfff;
rom[78068] = 12'hfff;
rom[78069] = 12'hfff;
rom[78070] = 12'hfff;
rom[78071] = 12'hfff;
rom[78072] = 12'hfff;
rom[78073] = 12'hfff;
rom[78074] = 12'hfff;
rom[78075] = 12'hfff;
rom[78076] = 12'hfff;
rom[78077] = 12'hfff;
rom[78078] = 12'hfff;
rom[78079] = 12'hfff;
rom[78080] = 12'hfff;
rom[78081] = 12'hfff;
rom[78082] = 12'hfff;
rom[78083] = 12'hfff;
rom[78084] = 12'hfff;
rom[78085] = 12'hfff;
rom[78086] = 12'hfff;
rom[78087] = 12'hfff;
rom[78088] = 12'hfff;
rom[78089] = 12'hfff;
rom[78090] = 12'hfff;
rom[78091] = 12'hfff;
rom[78092] = 12'hfff;
rom[78093] = 12'hfff;
rom[78094] = 12'hfff;
rom[78095] = 12'hfff;
rom[78096] = 12'hfff;
rom[78097] = 12'hfff;
rom[78098] = 12'hfff;
rom[78099] = 12'hfff;
rom[78100] = 12'hfff;
rom[78101] = 12'hfff;
rom[78102] = 12'hfff;
rom[78103] = 12'hfff;
rom[78104] = 12'hfff;
rom[78105] = 12'hfff;
rom[78106] = 12'hfff;
rom[78107] = 12'hfff;
rom[78108] = 12'hfff;
rom[78109] = 12'hfff;
rom[78110] = 12'hfff;
rom[78111] = 12'hfff;
rom[78112] = 12'hfff;
rom[78113] = 12'hfff;
rom[78114] = 12'hfff;
rom[78115] = 12'hfff;
rom[78116] = 12'hfff;
rom[78117] = 12'heee;
rom[78118] = 12'heee;
rom[78119] = 12'hddd;
rom[78120] = 12'hddd;
rom[78121] = 12'hccc;
rom[78122] = 12'hccc;
rom[78123] = 12'hccc;
rom[78124] = 12'hbbb;
rom[78125] = 12'hbbb;
rom[78126] = 12'hbbb;
rom[78127] = 12'haaa;
rom[78128] = 12'h999;
rom[78129] = 12'h999;
rom[78130] = 12'h888;
rom[78131] = 12'h888;
rom[78132] = 12'h888;
rom[78133] = 12'h888;
rom[78134] = 12'h888;
rom[78135] = 12'h888;
rom[78136] = 12'h888;
rom[78137] = 12'h888;
rom[78138] = 12'h888;
rom[78139] = 12'h888;
rom[78140] = 12'h888;
rom[78141] = 12'h888;
rom[78142] = 12'h888;
rom[78143] = 12'h888;
rom[78144] = 12'h888;
rom[78145] = 12'h888;
rom[78146] = 12'h888;
rom[78147] = 12'h888;
rom[78148] = 12'h888;
rom[78149] = 12'h777;
rom[78150] = 12'h777;
rom[78151] = 12'h777;
rom[78152] = 12'h777;
rom[78153] = 12'h666;
rom[78154] = 12'h666;
rom[78155] = 12'h666;
rom[78156] = 12'h666;
rom[78157] = 12'h666;
rom[78158] = 12'h666;
rom[78159] = 12'h666;
rom[78160] = 12'h555;
rom[78161] = 12'h666;
rom[78162] = 12'h666;
rom[78163] = 12'h666;
rom[78164] = 12'h666;
rom[78165] = 12'h666;
rom[78166] = 12'h666;
rom[78167] = 12'h555;
rom[78168] = 12'h555;
rom[78169] = 12'h555;
rom[78170] = 12'h555;
rom[78171] = 12'h555;
rom[78172] = 12'h555;
rom[78173] = 12'h555;
rom[78174] = 12'h555;
rom[78175] = 12'h555;
rom[78176] = 12'h555;
rom[78177] = 12'h555;
rom[78178] = 12'h555;
rom[78179] = 12'h555;
rom[78180] = 12'h555;
rom[78181] = 12'h555;
rom[78182] = 12'h555;
rom[78183] = 12'h444;
rom[78184] = 12'h444;
rom[78185] = 12'h444;
rom[78186] = 12'h444;
rom[78187] = 12'h444;
rom[78188] = 12'h444;
rom[78189] = 12'h555;
rom[78190] = 12'h555;
rom[78191] = 12'h555;
rom[78192] = 12'h555;
rom[78193] = 12'h555;
rom[78194] = 12'h555;
rom[78195] = 12'h666;
rom[78196] = 12'h777;
rom[78197] = 12'h777;
rom[78198] = 12'h777;
rom[78199] = 12'h777;
rom[78200] = 12'h888;
rom[78201] = 12'h888;
rom[78202] = 12'h888;
rom[78203] = 12'h888;
rom[78204] = 12'h777;
rom[78205] = 12'h666;
rom[78206] = 12'h555;
rom[78207] = 12'h555;
rom[78208] = 12'h444;
rom[78209] = 12'h444;
rom[78210] = 12'h444;
rom[78211] = 12'h444;
rom[78212] = 12'h333;
rom[78213] = 12'h333;
rom[78214] = 12'h333;
rom[78215] = 12'h333;
rom[78216] = 12'h333;
rom[78217] = 12'h333;
rom[78218] = 12'h333;
rom[78219] = 12'h333;
rom[78220] = 12'h333;
rom[78221] = 12'h333;
rom[78222] = 12'h222;
rom[78223] = 12'h222;
rom[78224] = 12'h222;
rom[78225] = 12'h222;
rom[78226] = 12'h222;
rom[78227] = 12'h222;
rom[78228] = 12'h222;
rom[78229] = 12'h222;
rom[78230] = 12'h111;
rom[78231] = 12'h111;
rom[78232] = 12'h111;
rom[78233] = 12'h111;
rom[78234] = 12'h111;
rom[78235] = 12'h  0;
rom[78236] = 12'h  0;
rom[78237] = 12'h  0;
rom[78238] = 12'h  0;
rom[78239] = 12'h  0;
rom[78240] = 12'h  0;
rom[78241] = 12'h  0;
rom[78242] = 12'h  0;
rom[78243] = 12'h  0;
rom[78244] = 12'h  0;
rom[78245] = 12'h  0;
rom[78246] = 12'h  0;
rom[78247] = 12'h  0;
rom[78248] = 12'h  0;
rom[78249] = 12'h  0;
rom[78250] = 12'h  0;
rom[78251] = 12'h  0;
rom[78252] = 12'h  0;
rom[78253] = 12'h  0;
rom[78254] = 12'h  0;
rom[78255] = 12'h  0;
rom[78256] = 12'h  0;
rom[78257] = 12'h  0;
rom[78258] = 12'h  0;
rom[78259] = 12'h  0;
rom[78260] = 12'h  0;
rom[78261] = 12'h  0;
rom[78262] = 12'h  0;
rom[78263] = 12'h  0;
rom[78264] = 12'h  0;
rom[78265] = 12'h  0;
rom[78266] = 12'h  0;
rom[78267] = 12'h  0;
rom[78268] = 12'h  0;
rom[78269] = 12'h111;
rom[78270] = 12'h111;
rom[78271] = 12'h111;
rom[78272] = 12'h111;
rom[78273] = 12'h111;
rom[78274] = 12'h222;
rom[78275] = 12'h333;
rom[78276] = 12'h333;
rom[78277] = 12'h444;
rom[78278] = 12'h666;
rom[78279] = 12'h888;
rom[78280] = 12'h888;
rom[78281] = 12'h777;
rom[78282] = 12'h555;
rom[78283] = 12'h333;
rom[78284] = 12'h333;
rom[78285] = 12'h333;
rom[78286] = 12'h222;
rom[78287] = 12'h333;
rom[78288] = 12'h333;
rom[78289] = 12'h333;
rom[78290] = 12'h333;
rom[78291] = 12'h333;
rom[78292] = 12'h333;
rom[78293] = 12'h333;
rom[78294] = 12'h333;
rom[78295] = 12'h333;
rom[78296] = 12'h444;
rom[78297] = 12'h444;
rom[78298] = 12'h444;
rom[78299] = 12'h444;
rom[78300] = 12'h555;
rom[78301] = 12'h555;
rom[78302] = 12'h555;
rom[78303] = 12'h555;
rom[78304] = 12'h666;
rom[78305] = 12'h666;
rom[78306] = 12'h666;
rom[78307] = 12'h777;
rom[78308] = 12'h777;
rom[78309] = 12'h888;
rom[78310] = 12'h999;
rom[78311] = 12'h999;
rom[78312] = 12'h999;
rom[78313] = 12'haaa;
rom[78314] = 12'hccc;
rom[78315] = 12'hddd;
rom[78316] = 12'heee;
rom[78317] = 12'hfff;
rom[78318] = 12'hfff;
rom[78319] = 12'hfff;
rom[78320] = 12'hfff;
rom[78321] = 12'hfff;
rom[78322] = 12'heee;
rom[78323] = 12'hddd;
rom[78324] = 12'hccc;
rom[78325] = 12'hbbb;
rom[78326] = 12'hbbb;
rom[78327] = 12'haaa;
rom[78328] = 12'haaa;
rom[78329] = 12'h999;
rom[78330] = 12'h999;
rom[78331] = 12'h888;
rom[78332] = 12'h888;
rom[78333] = 12'h888;
rom[78334] = 12'h777;
rom[78335] = 12'h777;
rom[78336] = 12'h666;
rom[78337] = 12'h666;
rom[78338] = 12'h666;
rom[78339] = 12'h666;
rom[78340] = 12'h666;
rom[78341] = 12'h555;
rom[78342] = 12'h555;
rom[78343] = 12'h555;
rom[78344] = 12'h555;
rom[78345] = 12'h555;
rom[78346] = 12'h555;
rom[78347] = 12'h555;
rom[78348] = 12'h444;
rom[78349] = 12'h444;
rom[78350] = 12'h444;
rom[78351] = 12'h444;
rom[78352] = 12'h444;
rom[78353] = 12'h444;
rom[78354] = 12'h444;
rom[78355] = 12'h444;
rom[78356] = 12'h444;
rom[78357] = 12'h444;
rom[78358] = 12'h444;
rom[78359] = 12'h444;
rom[78360] = 12'h444;
rom[78361] = 12'h444;
rom[78362] = 12'h444;
rom[78363] = 12'h444;
rom[78364] = 12'h444;
rom[78365] = 12'h444;
rom[78366] = 12'h444;
rom[78367] = 12'h444;
rom[78368] = 12'h333;
rom[78369] = 12'h333;
rom[78370] = 12'h333;
rom[78371] = 12'h333;
rom[78372] = 12'h333;
rom[78373] = 12'h333;
rom[78374] = 12'h333;
rom[78375] = 12'h333;
rom[78376] = 12'h333;
rom[78377] = 12'h333;
rom[78378] = 12'h333;
rom[78379] = 12'h333;
rom[78380] = 12'h333;
rom[78381] = 12'h333;
rom[78382] = 12'h333;
rom[78383] = 12'h333;
rom[78384] = 12'h333;
rom[78385] = 12'h333;
rom[78386] = 12'h333;
rom[78387] = 12'h333;
rom[78388] = 12'h333;
rom[78389] = 12'h333;
rom[78390] = 12'h333;
rom[78391] = 12'h333;
rom[78392] = 12'h333;
rom[78393] = 12'h333;
rom[78394] = 12'h333;
rom[78395] = 12'h333;
rom[78396] = 12'h333;
rom[78397] = 12'h333;
rom[78398] = 12'h333;
rom[78399] = 12'h333;
rom[78400] = 12'hfff;
rom[78401] = 12'hfff;
rom[78402] = 12'hfff;
rom[78403] = 12'hfff;
rom[78404] = 12'hfff;
rom[78405] = 12'hfff;
rom[78406] = 12'hfff;
rom[78407] = 12'hfff;
rom[78408] = 12'hfff;
rom[78409] = 12'hfff;
rom[78410] = 12'hfff;
rom[78411] = 12'hfff;
rom[78412] = 12'hfff;
rom[78413] = 12'hfff;
rom[78414] = 12'hfff;
rom[78415] = 12'hfff;
rom[78416] = 12'hfff;
rom[78417] = 12'hfff;
rom[78418] = 12'hfff;
rom[78419] = 12'hfff;
rom[78420] = 12'hfff;
rom[78421] = 12'hfff;
rom[78422] = 12'hfff;
rom[78423] = 12'hfff;
rom[78424] = 12'hfff;
rom[78425] = 12'hfff;
rom[78426] = 12'hfff;
rom[78427] = 12'hfff;
rom[78428] = 12'hfff;
rom[78429] = 12'hfff;
rom[78430] = 12'hfff;
rom[78431] = 12'hfff;
rom[78432] = 12'hfff;
rom[78433] = 12'hfff;
rom[78434] = 12'hfff;
rom[78435] = 12'hfff;
rom[78436] = 12'hfff;
rom[78437] = 12'hfff;
rom[78438] = 12'hfff;
rom[78439] = 12'hfff;
rom[78440] = 12'hfff;
rom[78441] = 12'hfff;
rom[78442] = 12'hfff;
rom[78443] = 12'hfff;
rom[78444] = 12'hfff;
rom[78445] = 12'hfff;
rom[78446] = 12'hfff;
rom[78447] = 12'hfff;
rom[78448] = 12'hfff;
rom[78449] = 12'hfff;
rom[78450] = 12'hfff;
rom[78451] = 12'hfff;
rom[78452] = 12'hfff;
rom[78453] = 12'hfff;
rom[78454] = 12'hfff;
rom[78455] = 12'hfff;
rom[78456] = 12'hfff;
rom[78457] = 12'hfff;
rom[78458] = 12'hfff;
rom[78459] = 12'hfff;
rom[78460] = 12'hfff;
rom[78461] = 12'hfff;
rom[78462] = 12'hfff;
rom[78463] = 12'hfff;
rom[78464] = 12'hfff;
rom[78465] = 12'hfff;
rom[78466] = 12'hfff;
rom[78467] = 12'hfff;
rom[78468] = 12'hfff;
rom[78469] = 12'hfff;
rom[78470] = 12'hfff;
rom[78471] = 12'hfff;
rom[78472] = 12'hfff;
rom[78473] = 12'hfff;
rom[78474] = 12'hfff;
rom[78475] = 12'hfff;
rom[78476] = 12'hfff;
rom[78477] = 12'hfff;
rom[78478] = 12'hfff;
rom[78479] = 12'hfff;
rom[78480] = 12'hfff;
rom[78481] = 12'hfff;
rom[78482] = 12'hfff;
rom[78483] = 12'hfff;
rom[78484] = 12'hfff;
rom[78485] = 12'hfff;
rom[78486] = 12'hfff;
rom[78487] = 12'hfff;
rom[78488] = 12'hfff;
rom[78489] = 12'hfff;
rom[78490] = 12'hfff;
rom[78491] = 12'hfff;
rom[78492] = 12'hfff;
rom[78493] = 12'hfff;
rom[78494] = 12'hfff;
rom[78495] = 12'hfff;
rom[78496] = 12'hfff;
rom[78497] = 12'hfff;
rom[78498] = 12'hfff;
rom[78499] = 12'hfff;
rom[78500] = 12'hfff;
rom[78501] = 12'hfff;
rom[78502] = 12'hfff;
rom[78503] = 12'hfff;
rom[78504] = 12'hfff;
rom[78505] = 12'hfff;
rom[78506] = 12'hfff;
rom[78507] = 12'hfff;
rom[78508] = 12'hfff;
rom[78509] = 12'hfff;
rom[78510] = 12'hfff;
rom[78511] = 12'hfff;
rom[78512] = 12'hfff;
rom[78513] = 12'hfff;
rom[78514] = 12'hfff;
rom[78515] = 12'hfff;
rom[78516] = 12'hfff;
rom[78517] = 12'hfff;
rom[78518] = 12'heee;
rom[78519] = 12'heee;
rom[78520] = 12'hddd;
rom[78521] = 12'hddd;
rom[78522] = 12'hddd;
rom[78523] = 12'hccc;
rom[78524] = 12'hccc;
rom[78525] = 12'hccc;
rom[78526] = 12'hbbb;
rom[78527] = 12'hbbb;
rom[78528] = 12'haaa;
rom[78529] = 12'haaa;
rom[78530] = 12'haaa;
rom[78531] = 12'haaa;
rom[78532] = 12'h999;
rom[78533] = 12'h999;
rom[78534] = 12'h999;
rom[78535] = 12'h999;
rom[78536] = 12'h999;
rom[78537] = 12'h999;
rom[78538] = 12'h999;
rom[78539] = 12'h999;
rom[78540] = 12'h999;
rom[78541] = 12'h999;
rom[78542] = 12'h999;
rom[78543] = 12'h999;
rom[78544] = 12'h888;
rom[78545] = 12'h888;
rom[78546] = 12'h888;
rom[78547] = 12'h888;
rom[78548] = 12'h888;
rom[78549] = 12'h777;
rom[78550] = 12'h777;
rom[78551] = 12'h777;
rom[78552] = 12'h666;
rom[78553] = 12'h666;
rom[78554] = 12'h666;
rom[78555] = 12'h666;
rom[78556] = 12'h666;
rom[78557] = 12'h666;
rom[78558] = 12'h555;
rom[78559] = 12'h555;
rom[78560] = 12'h555;
rom[78561] = 12'h555;
rom[78562] = 12'h555;
rom[78563] = 12'h555;
rom[78564] = 12'h666;
rom[78565] = 12'h666;
rom[78566] = 12'h555;
rom[78567] = 12'h555;
rom[78568] = 12'h555;
rom[78569] = 12'h555;
rom[78570] = 12'h555;
rom[78571] = 12'h555;
rom[78572] = 12'h444;
rom[78573] = 12'h444;
rom[78574] = 12'h444;
rom[78575] = 12'h444;
rom[78576] = 12'h444;
rom[78577] = 12'h444;
rom[78578] = 12'h444;
rom[78579] = 12'h444;
rom[78580] = 12'h444;
rom[78581] = 12'h444;
rom[78582] = 12'h444;
rom[78583] = 12'h444;
rom[78584] = 12'h444;
rom[78585] = 12'h444;
rom[78586] = 12'h555;
rom[78587] = 12'h555;
rom[78588] = 12'h555;
rom[78589] = 12'h555;
rom[78590] = 12'h555;
rom[78591] = 12'h555;
rom[78592] = 12'h555;
rom[78593] = 12'h555;
rom[78594] = 12'h555;
rom[78595] = 12'h666;
rom[78596] = 12'h666;
rom[78597] = 12'h777;
rom[78598] = 12'h777;
rom[78599] = 12'h777;
rom[78600] = 12'h888;
rom[78601] = 12'h888;
rom[78602] = 12'h888;
rom[78603] = 12'h888;
rom[78604] = 12'h888;
rom[78605] = 12'h777;
rom[78606] = 12'h666;
rom[78607] = 12'h555;
rom[78608] = 12'h444;
rom[78609] = 12'h444;
rom[78610] = 12'h444;
rom[78611] = 12'h444;
rom[78612] = 12'h333;
rom[78613] = 12'h333;
rom[78614] = 12'h333;
rom[78615] = 12'h333;
rom[78616] = 12'h333;
rom[78617] = 12'h333;
rom[78618] = 12'h333;
rom[78619] = 12'h333;
rom[78620] = 12'h333;
rom[78621] = 12'h333;
rom[78622] = 12'h333;
rom[78623] = 12'h222;
rom[78624] = 12'h222;
rom[78625] = 12'h222;
rom[78626] = 12'h222;
rom[78627] = 12'h222;
rom[78628] = 12'h222;
rom[78629] = 12'h222;
rom[78630] = 12'h111;
rom[78631] = 12'h111;
rom[78632] = 12'h111;
rom[78633] = 12'h111;
rom[78634] = 12'h111;
rom[78635] = 12'h  0;
rom[78636] = 12'h  0;
rom[78637] = 12'h  0;
rom[78638] = 12'h  0;
rom[78639] = 12'h  0;
rom[78640] = 12'h  0;
rom[78641] = 12'h  0;
rom[78642] = 12'h  0;
rom[78643] = 12'h  0;
rom[78644] = 12'h  0;
rom[78645] = 12'h  0;
rom[78646] = 12'h  0;
rom[78647] = 12'h  0;
rom[78648] = 12'h  0;
rom[78649] = 12'h  0;
rom[78650] = 12'h  0;
rom[78651] = 12'h  0;
rom[78652] = 12'h  0;
rom[78653] = 12'h  0;
rom[78654] = 12'h  0;
rom[78655] = 12'h  0;
rom[78656] = 12'h  0;
rom[78657] = 12'h  0;
rom[78658] = 12'h  0;
rom[78659] = 12'h  0;
rom[78660] = 12'h  0;
rom[78661] = 12'h  0;
rom[78662] = 12'h  0;
rom[78663] = 12'h  0;
rom[78664] = 12'h  0;
rom[78665] = 12'h  0;
rom[78666] = 12'h  0;
rom[78667] = 12'h  0;
rom[78668] = 12'h  0;
rom[78669] = 12'h111;
rom[78670] = 12'h111;
rom[78671] = 12'h111;
rom[78672] = 12'h111;
rom[78673] = 12'h111;
rom[78674] = 12'h222;
rom[78675] = 12'h333;
rom[78676] = 12'h333;
rom[78677] = 12'h444;
rom[78678] = 12'h666;
rom[78679] = 12'h777;
rom[78680] = 12'h888;
rom[78681] = 12'h777;
rom[78682] = 12'h555;
rom[78683] = 12'h444;
rom[78684] = 12'h333;
rom[78685] = 12'h333;
rom[78686] = 12'h222;
rom[78687] = 12'h333;
rom[78688] = 12'h333;
rom[78689] = 12'h333;
rom[78690] = 12'h333;
rom[78691] = 12'h333;
rom[78692] = 12'h333;
rom[78693] = 12'h333;
rom[78694] = 12'h444;
rom[78695] = 12'h444;
rom[78696] = 12'h444;
rom[78697] = 12'h444;
rom[78698] = 12'h444;
rom[78699] = 12'h555;
rom[78700] = 12'h555;
rom[78701] = 12'h555;
rom[78702] = 12'h555;
rom[78703] = 12'h666;
rom[78704] = 12'h666;
rom[78705] = 12'h777;
rom[78706] = 12'h777;
rom[78707] = 12'h888;
rom[78708] = 12'h888;
rom[78709] = 12'h888;
rom[78710] = 12'h999;
rom[78711] = 12'h999;
rom[78712] = 12'haaa;
rom[78713] = 12'hbbb;
rom[78714] = 12'hccc;
rom[78715] = 12'hddd;
rom[78716] = 12'heee;
rom[78717] = 12'hfff;
rom[78718] = 12'hfff;
rom[78719] = 12'hfff;
rom[78720] = 12'hfff;
rom[78721] = 12'heee;
rom[78722] = 12'hddd;
rom[78723] = 12'hccc;
rom[78724] = 12'hbbb;
rom[78725] = 12'hbbb;
rom[78726] = 12'haaa;
rom[78727] = 12'haaa;
rom[78728] = 12'h999;
rom[78729] = 12'h999;
rom[78730] = 12'h888;
rom[78731] = 12'h888;
rom[78732] = 12'h888;
rom[78733] = 12'h888;
rom[78734] = 12'h777;
rom[78735] = 12'h777;
rom[78736] = 12'h666;
rom[78737] = 12'h666;
rom[78738] = 12'h666;
rom[78739] = 12'h666;
rom[78740] = 12'h555;
rom[78741] = 12'h555;
rom[78742] = 12'h555;
rom[78743] = 12'h555;
rom[78744] = 12'h555;
rom[78745] = 12'h555;
rom[78746] = 12'h444;
rom[78747] = 12'h444;
rom[78748] = 12'h444;
rom[78749] = 12'h444;
rom[78750] = 12'h444;
rom[78751] = 12'h444;
rom[78752] = 12'h333;
rom[78753] = 12'h333;
rom[78754] = 12'h333;
rom[78755] = 12'h333;
rom[78756] = 12'h444;
rom[78757] = 12'h444;
rom[78758] = 12'h444;
rom[78759] = 12'h444;
rom[78760] = 12'h444;
rom[78761] = 12'h444;
rom[78762] = 12'h444;
rom[78763] = 12'h444;
rom[78764] = 12'h444;
rom[78765] = 12'h444;
rom[78766] = 12'h444;
rom[78767] = 12'h444;
rom[78768] = 12'h333;
rom[78769] = 12'h333;
rom[78770] = 12'h333;
rom[78771] = 12'h333;
rom[78772] = 12'h333;
rom[78773] = 12'h333;
rom[78774] = 12'h333;
rom[78775] = 12'h333;
rom[78776] = 12'h333;
rom[78777] = 12'h333;
rom[78778] = 12'h333;
rom[78779] = 12'h333;
rom[78780] = 12'h333;
rom[78781] = 12'h333;
rom[78782] = 12'h333;
rom[78783] = 12'h333;
rom[78784] = 12'h333;
rom[78785] = 12'h333;
rom[78786] = 12'h333;
rom[78787] = 12'h333;
rom[78788] = 12'h333;
rom[78789] = 12'h333;
rom[78790] = 12'h333;
rom[78791] = 12'h333;
rom[78792] = 12'h333;
rom[78793] = 12'h333;
rom[78794] = 12'h333;
rom[78795] = 12'h333;
rom[78796] = 12'h333;
rom[78797] = 12'h333;
rom[78798] = 12'h333;
rom[78799] = 12'h333;
rom[78800] = 12'hfff;
rom[78801] = 12'hfff;
rom[78802] = 12'hfff;
rom[78803] = 12'hfff;
rom[78804] = 12'hfff;
rom[78805] = 12'hfff;
rom[78806] = 12'hfff;
rom[78807] = 12'hfff;
rom[78808] = 12'hfff;
rom[78809] = 12'hfff;
rom[78810] = 12'hfff;
rom[78811] = 12'hfff;
rom[78812] = 12'hfff;
rom[78813] = 12'hfff;
rom[78814] = 12'hfff;
rom[78815] = 12'hfff;
rom[78816] = 12'hfff;
rom[78817] = 12'hfff;
rom[78818] = 12'hfff;
rom[78819] = 12'hfff;
rom[78820] = 12'hfff;
rom[78821] = 12'hfff;
rom[78822] = 12'hfff;
rom[78823] = 12'hfff;
rom[78824] = 12'hfff;
rom[78825] = 12'hfff;
rom[78826] = 12'hfff;
rom[78827] = 12'hfff;
rom[78828] = 12'hfff;
rom[78829] = 12'hfff;
rom[78830] = 12'hfff;
rom[78831] = 12'hfff;
rom[78832] = 12'hfff;
rom[78833] = 12'hfff;
rom[78834] = 12'hfff;
rom[78835] = 12'hfff;
rom[78836] = 12'hfff;
rom[78837] = 12'hfff;
rom[78838] = 12'hfff;
rom[78839] = 12'hfff;
rom[78840] = 12'hfff;
rom[78841] = 12'hfff;
rom[78842] = 12'hfff;
rom[78843] = 12'hfff;
rom[78844] = 12'hfff;
rom[78845] = 12'hfff;
rom[78846] = 12'hfff;
rom[78847] = 12'hfff;
rom[78848] = 12'hfff;
rom[78849] = 12'hfff;
rom[78850] = 12'hfff;
rom[78851] = 12'hfff;
rom[78852] = 12'hfff;
rom[78853] = 12'hfff;
rom[78854] = 12'hfff;
rom[78855] = 12'hfff;
rom[78856] = 12'hfff;
rom[78857] = 12'hfff;
rom[78858] = 12'hfff;
rom[78859] = 12'hfff;
rom[78860] = 12'hfff;
rom[78861] = 12'hfff;
rom[78862] = 12'hfff;
rom[78863] = 12'hfff;
rom[78864] = 12'hfff;
rom[78865] = 12'hfff;
rom[78866] = 12'hfff;
rom[78867] = 12'hfff;
rom[78868] = 12'hfff;
rom[78869] = 12'hfff;
rom[78870] = 12'hfff;
rom[78871] = 12'hfff;
rom[78872] = 12'hfff;
rom[78873] = 12'hfff;
rom[78874] = 12'hfff;
rom[78875] = 12'hfff;
rom[78876] = 12'hfff;
rom[78877] = 12'hfff;
rom[78878] = 12'hfff;
rom[78879] = 12'hfff;
rom[78880] = 12'hfff;
rom[78881] = 12'hfff;
rom[78882] = 12'hfff;
rom[78883] = 12'hfff;
rom[78884] = 12'hfff;
rom[78885] = 12'hfff;
rom[78886] = 12'hfff;
rom[78887] = 12'hfff;
rom[78888] = 12'hfff;
rom[78889] = 12'hfff;
rom[78890] = 12'hfff;
rom[78891] = 12'hfff;
rom[78892] = 12'hfff;
rom[78893] = 12'hfff;
rom[78894] = 12'hfff;
rom[78895] = 12'hfff;
rom[78896] = 12'hfff;
rom[78897] = 12'hfff;
rom[78898] = 12'hfff;
rom[78899] = 12'hfff;
rom[78900] = 12'hfff;
rom[78901] = 12'hfff;
rom[78902] = 12'hfff;
rom[78903] = 12'hfff;
rom[78904] = 12'hfff;
rom[78905] = 12'hfff;
rom[78906] = 12'hfff;
rom[78907] = 12'hfff;
rom[78908] = 12'hfff;
rom[78909] = 12'hfff;
rom[78910] = 12'hfff;
rom[78911] = 12'hfff;
rom[78912] = 12'hfff;
rom[78913] = 12'hfff;
rom[78914] = 12'hfff;
rom[78915] = 12'hfff;
rom[78916] = 12'hfff;
rom[78917] = 12'hfff;
rom[78918] = 12'hfff;
rom[78919] = 12'hfff;
rom[78920] = 12'heee;
rom[78921] = 12'heee;
rom[78922] = 12'hddd;
rom[78923] = 12'hddd;
rom[78924] = 12'hddd;
rom[78925] = 12'hccc;
rom[78926] = 12'hccc;
rom[78927] = 12'hccc;
rom[78928] = 12'hccc;
rom[78929] = 12'hbbb;
rom[78930] = 12'hbbb;
rom[78931] = 12'hbbb;
rom[78932] = 12'haaa;
rom[78933] = 12'haaa;
rom[78934] = 12'haaa;
rom[78935] = 12'haaa;
rom[78936] = 12'haaa;
rom[78937] = 12'haaa;
rom[78938] = 12'h999;
rom[78939] = 12'h999;
rom[78940] = 12'h999;
rom[78941] = 12'h999;
rom[78942] = 12'h999;
rom[78943] = 12'h999;
rom[78944] = 12'h888;
rom[78945] = 12'h888;
rom[78946] = 12'h888;
rom[78947] = 12'h777;
rom[78948] = 12'h777;
rom[78949] = 12'h777;
rom[78950] = 12'h777;
rom[78951] = 12'h666;
rom[78952] = 12'h666;
rom[78953] = 12'h555;
rom[78954] = 12'h555;
rom[78955] = 12'h555;
rom[78956] = 12'h555;
rom[78957] = 12'h555;
rom[78958] = 12'h555;
rom[78959] = 12'h555;
rom[78960] = 12'h444;
rom[78961] = 12'h555;
rom[78962] = 12'h555;
rom[78963] = 12'h555;
rom[78964] = 12'h555;
rom[78965] = 12'h555;
rom[78966] = 12'h555;
rom[78967] = 12'h555;
rom[78968] = 12'h555;
rom[78969] = 12'h555;
rom[78970] = 12'h555;
rom[78971] = 12'h555;
rom[78972] = 12'h555;
rom[78973] = 12'h444;
rom[78974] = 12'h444;
rom[78975] = 12'h444;
rom[78976] = 12'h444;
rom[78977] = 12'h444;
rom[78978] = 12'h444;
rom[78979] = 12'h444;
rom[78980] = 12'h444;
rom[78981] = 12'h444;
rom[78982] = 12'h444;
rom[78983] = 12'h444;
rom[78984] = 12'h444;
rom[78985] = 12'h444;
rom[78986] = 12'h555;
rom[78987] = 12'h555;
rom[78988] = 12'h555;
rom[78989] = 12'h555;
rom[78990] = 12'h555;
rom[78991] = 12'h555;
rom[78992] = 12'h555;
rom[78993] = 12'h555;
rom[78994] = 12'h555;
rom[78995] = 12'h666;
rom[78996] = 12'h666;
rom[78997] = 12'h777;
rom[78998] = 12'h777;
rom[78999] = 12'h888;
rom[79000] = 12'h888;
rom[79001] = 12'h888;
rom[79002] = 12'h999;
rom[79003] = 12'h999;
rom[79004] = 12'h888;
rom[79005] = 12'h888;
rom[79006] = 12'h777;
rom[79007] = 12'h555;
rom[79008] = 12'h555;
rom[79009] = 12'h555;
rom[79010] = 12'h444;
rom[79011] = 12'h444;
rom[79012] = 12'h333;
rom[79013] = 12'h333;
rom[79014] = 12'h333;
rom[79015] = 12'h333;
rom[79016] = 12'h333;
rom[79017] = 12'h333;
rom[79018] = 12'h333;
rom[79019] = 12'h333;
rom[79020] = 12'h333;
rom[79021] = 12'h333;
rom[79022] = 12'h333;
rom[79023] = 12'h333;
rom[79024] = 12'h333;
rom[79025] = 12'h333;
rom[79026] = 12'h222;
rom[79027] = 12'h222;
rom[79028] = 12'h222;
rom[79029] = 12'h222;
rom[79030] = 12'h111;
rom[79031] = 12'h111;
rom[79032] = 12'h111;
rom[79033] = 12'h111;
rom[79034] = 12'h111;
rom[79035] = 12'h  0;
rom[79036] = 12'h  0;
rom[79037] = 12'h  0;
rom[79038] = 12'h  0;
rom[79039] = 12'h  0;
rom[79040] = 12'h  0;
rom[79041] = 12'h  0;
rom[79042] = 12'h  0;
rom[79043] = 12'h  0;
rom[79044] = 12'h  0;
rom[79045] = 12'h  0;
rom[79046] = 12'h  0;
rom[79047] = 12'h  0;
rom[79048] = 12'h  0;
rom[79049] = 12'h  0;
rom[79050] = 12'h  0;
rom[79051] = 12'h  0;
rom[79052] = 12'h  0;
rom[79053] = 12'h  0;
rom[79054] = 12'h  0;
rom[79055] = 12'h  0;
rom[79056] = 12'h  0;
rom[79057] = 12'h  0;
rom[79058] = 12'h  0;
rom[79059] = 12'h  0;
rom[79060] = 12'h  0;
rom[79061] = 12'h  0;
rom[79062] = 12'h  0;
rom[79063] = 12'h  0;
rom[79064] = 12'h  0;
rom[79065] = 12'h  0;
rom[79066] = 12'h  0;
rom[79067] = 12'h  0;
rom[79068] = 12'h  0;
rom[79069] = 12'h111;
rom[79070] = 12'h111;
rom[79071] = 12'h111;
rom[79072] = 12'h111;
rom[79073] = 12'h111;
rom[79074] = 12'h222;
rom[79075] = 12'h333;
rom[79076] = 12'h333;
rom[79077] = 12'h444;
rom[79078] = 12'h555;
rom[79079] = 12'h777;
rom[79080] = 12'h999;
rom[79081] = 12'h888;
rom[79082] = 12'h555;
rom[79083] = 12'h444;
rom[79084] = 12'h444;
rom[79085] = 12'h333;
rom[79086] = 12'h333;
rom[79087] = 12'h333;
rom[79088] = 12'h333;
rom[79089] = 12'h333;
rom[79090] = 12'h333;
rom[79091] = 12'h333;
rom[79092] = 12'h333;
rom[79093] = 12'h444;
rom[79094] = 12'h444;
rom[79095] = 12'h444;
rom[79096] = 12'h444;
rom[79097] = 12'h444;
rom[79098] = 12'h555;
rom[79099] = 12'h555;
rom[79100] = 12'h555;
rom[79101] = 12'h555;
rom[79102] = 12'h666;
rom[79103] = 12'h666;
rom[79104] = 12'h666;
rom[79105] = 12'h777;
rom[79106] = 12'h888;
rom[79107] = 12'h888;
rom[79108] = 12'h888;
rom[79109] = 12'h999;
rom[79110] = 12'h999;
rom[79111] = 12'h999;
rom[79112] = 12'haaa;
rom[79113] = 12'hbbb;
rom[79114] = 12'hddd;
rom[79115] = 12'heee;
rom[79116] = 12'hfff;
rom[79117] = 12'hfff;
rom[79118] = 12'hfff;
rom[79119] = 12'heee;
rom[79120] = 12'hddd;
rom[79121] = 12'hddd;
rom[79122] = 12'hccc;
rom[79123] = 12'hbbb;
rom[79124] = 12'hbbb;
rom[79125] = 12'haaa;
rom[79126] = 12'haaa;
rom[79127] = 12'h999;
rom[79128] = 12'h999;
rom[79129] = 12'h888;
rom[79130] = 12'h888;
rom[79131] = 12'h888;
rom[79132] = 12'h777;
rom[79133] = 12'h777;
rom[79134] = 12'h777;
rom[79135] = 12'h666;
rom[79136] = 12'h666;
rom[79137] = 12'h666;
rom[79138] = 12'h555;
rom[79139] = 12'h555;
rom[79140] = 12'h555;
rom[79141] = 12'h555;
rom[79142] = 12'h444;
rom[79143] = 12'h444;
rom[79144] = 12'h444;
rom[79145] = 12'h444;
rom[79146] = 12'h444;
rom[79147] = 12'h444;
rom[79148] = 12'h444;
rom[79149] = 12'h444;
rom[79150] = 12'h444;
rom[79151] = 12'h444;
rom[79152] = 12'h333;
rom[79153] = 12'h333;
rom[79154] = 12'h333;
rom[79155] = 12'h333;
rom[79156] = 12'h333;
rom[79157] = 12'h333;
rom[79158] = 12'h444;
rom[79159] = 12'h444;
rom[79160] = 12'h444;
rom[79161] = 12'h444;
rom[79162] = 12'h444;
rom[79163] = 12'h444;
rom[79164] = 12'h444;
rom[79165] = 12'h444;
rom[79166] = 12'h444;
rom[79167] = 12'h444;
rom[79168] = 12'h333;
rom[79169] = 12'h333;
rom[79170] = 12'h333;
rom[79171] = 12'h333;
rom[79172] = 12'h333;
rom[79173] = 12'h333;
rom[79174] = 12'h333;
rom[79175] = 12'h333;
rom[79176] = 12'h333;
rom[79177] = 12'h333;
rom[79178] = 12'h333;
rom[79179] = 12'h333;
rom[79180] = 12'h333;
rom[79181] = 12'h333;
rom[79182] = 12'h333;
rom[79183] = 12'h333;
rom[79184] = 12'h333;
rom[79185] = 12'h222;
rom[79186] = 12'h222;
rom[79187] = 12'h222;
rom[79188] = 12'h222;
rom[79189] = 12'h222;
rom[79190] = 12'h222;
rom[79191] = 12'h333;
rom[79192] = 12'h333;
rom[79193] = 12'h333;
rom[79194] = 12'h333;
rom[79195] = 12'h333;
rom[79196] = 12'h333;
rom[79197] = 12'h333;
rom[79198] = 12'h333;
rom[79199] = 12'h333;
rom[79200] = 12'hfff;
rom[79201] = 12'hfff;
rom[79202] = 12'hfff;
rom[79203] = 12'hfff;
rom[79204] = 12'hfff;
rom[79205] = 12'hfff;
rom[79206] = 12'hfff;
rom[79207] = 12'hfff;
rom[79208] = 12'hfff;
rom[79209] = 12'hfff;
rom[79210] = 12'hfff;
rom[79211] = 12'hfff;
rom[79212] = 12'hfff;
rom[79213] = 12'hfff;
rom[79214] = 12'hfff;
rom[79215] = 12'hfff;
rom[79216] = 12'hfff;
rom[79217] = 12'hfff;
rom[79218] = 12'hfff;
rom[79219] = 12'hfff;
rom[79220] = 12'hfff;
rom[79221] = 12'hfff;
rom[79222] = 12'hfff;
rom[79223] = 12'hfff;
rom[79224] = 12'hfff;
rom[79225] = 12'hfff;
rom[79226] = 12'hfff;
rom[79227] = 12'hfff;
rom[79228] = 12'hfff;
rom[79229] = 12'hfff;
rom[79230] = 12'hfff;
rom[79231] = 12'hfff;
rom[79232] = 12'hfff;
rom[79233] = 12'hfff;
rom[79234] = 12'hfff;
rom[79235] = 12'hfff;
rom[79236] = 12'hfff;
rom[79237] = 12'hfff;
rom[79238] = 12'hfff;
rom[79239] = 12'hfff;
rom[79240] = 12'hfff;
rom[79241] = 12'hfff;
rom[79242] = 12'hfff;
rom[79243] = 12'hfff;
rom[79244] = 12'hfff;
rom[79245] = 12'hfff;
rom[79246] = 12'hfff;
rom[79247] = 12'hfff;
rom[79248] = 12'hfff;
rom[79249] = 12'hfff;
rom[79250] = 12'hfff;
rom[79251] = 12'hfff;
rom[79252] = 12'hfff;
rom[79253] = 12'hfff;
rom[79254] = 12'hfff;
rom[79255] = 12'hfff;
rom[79256] = 12'hfff;
rom[79257] = 12'hfff;
rom[79258] = 12'hfff;
rom[79259] = 12'hfff;
rom[79260] = 12'hfff;
rom[79261] = 12'hfff;
rom[79262] = 12'hfff;
rom[79263] = 12'hfff;
rom[79264] = 12'hfff;
rom[79265] = 12'hfff;
rom[79266] = 12'hfff;
rom[79267] = 12'hfff;
rom[79268] = 12'hfff;
rom[79269] = 12'hfff;
rom[79270] = 12'hfff;
rom[79271] = 12'hfff;
rom[79272] = 12'hfff;
rom[79273] = 12'hfff;
rom[79274] = 12'hfff;
rom[79275] = 12'hfff;
rom[79276] = 12'hfff;
rom[79277] = 12'hfff;
rom[79278] = 12'hfff;
rom[79279] = 12'hfff;
rom[79280] = 12'hfff;
rom[79281] = 12'hfff;
rom[79282] = 12'hfff;
rom[79283] = 12'hfff;
rom[79284] = 12'hfff;
rom[79285] = 12'hfff;
rom[79286] = 12'hfff;
rom[79287] = 12'hfff;
rom[79288] = 12'hfff;
rom[79289] = 12'hfff;
rom[79290] = 12'hfff;
rom[79291] = 12'hfff;
rom[79292] = 12'hfff;
rom[79293] = 12'hfff;
rom[79294] = 12'hfff;
rom[79295] = 12'hfff;
rom[79296] = 12'hfff;
rom[79297] = 12'hfff;
rom[79298] = 12'hfff;
rom[79299] = 12'hfff;
rom[79300] = 12'hfff;
rom[79301] = 12'hfff;
rom[79302] = 12'hfff;
rom[79303] = 12'hfff;
rom[79304] = 12'hfff;
rom[79305] = 12'hfff;
rom[79306] = 12'hfff;
rom[79307] = 12'hfff;
rom[79308] = 12'hfff;
rom[79309] = 12'hfff;
rom[79310] = 12'hfff;
rom[79311] = 12'hfff;
rom[79312] = 12'hfff;
rom[79313] = 12'hfff;
rom[79314] = 12'hfff;
rom[79315] = 12'hfff;
rom[79316] = 12'hfff;
rom[79317] = 12'hfff;
rom[79318] = 12'hfff;
rom[79319] = 12'hfff;
rom[79320] = 12'hfff;
rom[79321] = 12'heee;
rom[79322] = 12'heee;
rom[79323] = 12'heee;
rom[79324] = 12'hddd;
rom[79325] = 12'hddd;
rom[79326] = 12'hccc;
rom[79327] = 12'hccc;
rom[79328] = 12'hccc;
rom[79329] = 12'hbbb;
rom[79330] = 12'hbbb;
rom[79331] = 12'hbbb;
rom[79332] = 12'haaa;
rom[79333] = 12'haaa;
rom[79334] = 12'haaa;
rom[79335] = 12'haaa;
rom[79336] = 12'haaa;
rom[79337] = 12'haaa;
rom[79338] = 12'haaa;
rom[79339] = 12'haaa;
rom[79340] = 12'h999;
rom[79341] = 12'h999;
rom[79342] = 12'h999;
rom[79343] = 12'h999;
rom[79344] = 12'h888;
rom[79345] = 12'h888;
rom[79346] = 12'h777;
rom[79347] = 12'h777;
rom[79348] = 12'h777;
rom[79349] = 12'h666;
rom[79350] = 12'h666;
rom[79351] = 12'h666;
rom[79352] = 12'h555;
rom[79353] = 12'h555;
rom[79354] = 12'h444;
rom[79355] = 12'h444;
rom[79356] = 12'h444;
rom[79357] = 12'h444;
rom[79358] = 12'h555;
rom[79359] = 12'h555;
rom[79360] = 12'h444;
rom[79361] = 12'h444;
rom[79362] = 12'h444;
rom[79363] = 12'h444;
rom[79364] = 12'h444;
rom[79365] = 12'h444;
rom[79366] = 12'h444;
rom[79367] = 12'h444;
rom[79368] = 12'h555;
rom[79369] = 12'h555;
rom[79370] = 12'h555;
rom[79371] = 12'h555;
rom[79372] = 12'h555;
rom[79373] = 12'h555;
rom[79374] = 12'h444;
rom[79375] = 12'h444;
rom[79376] = 12'h444;
rom[79377] = 12'h444;
rom[79378] = 12'h444;
rom[79379] = 12'h444;
rom[79380] = 12'h444;
rom[79381] = 12'h444;
rom[79382] = 12'h444;
rom[79383] = 12'h444;
rom[79384] = 12'h444;
rom[79385] = 12'h444;
rom[79386] = 12'h444;
rom[79387] = 12'h444;
rom[79388] = 12'h555;
rom[79389] = 12'h555;
rom[79390] = 12'h555;
rom[79391] = 12'h555;
rom[79392] = 12'h555;
rom[79393] = 12'h555;
rom[79394] = 12'h555;
rom[79395] = 12'h666;
rom[79396] = 12'h666;
rom[79397] = 12'h666;
rom[79398] = 12'h777;
rom[79399] = 12'h777;
rom[79400] = 12'h888;
rom[79401] = 12'h999;
rom[79402] = 12'h999;
rom[79403] = 12'h999;
rom[79404] = 12'h999;
rom[79405] = 12'h999;
rom[79406] = 12'h888;
rom[79407] = 12'h666;
rom[79408] = 12'h666;
rom[79409] = 12'h555;
rom[79410] = 12'h555;
rom[79411] = 12'h444;
rom[79412] = 12'h444;
rom[79413] = 12'h444;
rom[79414] = 12'h444;
rom[79415] = 12'h333;
rom[79416] = 12'h333;
rom[79417] = 12'h333;
rom[79418] = 12'h333;
rom[79419] = 12'h333;
rom[79420] = 12'h333;
rom[79421] = 12'h333;
rom[79422] = 12'h333;
rom[79423] = 12'h333;
rom[79424] = 12'h333;
rom[79425] = 12'h333;
rom[79426] = 12'h222;
rom[79427] = 12'h222;
rom[79428] = 12'h222;
rom[79429] = 12'h111;
rom[79430] = 12'h111;
rom[79431] = 12'h111;
rom[79432] = 12'h111;
rom[79433] = 12'h111;
rom[79434] = 12'h111;
rom[79435] = 12'h  0;
rom[79436] = 12'h  0;
rom[79437] = 12'h  0;
rom[79438] = 12'h  0;
rom[79439] = 12'h  0;
rom[79440] = 12'h  0;
rom[79441] = 12'h  0;
rom[79442] = 12'h  0;
rom[79443] = 12'h  0;
rom[79444] = 12'h  0;
rom[79445] = 12'h  0;
rom[79446] = 12'h  0;
rom[79447] = 12'h  0;
rom[79448] = 12'h  0;
rom[79449] = 12'h  0;
rom[79450] = 12'h  0;
rom[79451] = 12'h  0;
rom[79452] = 12'h  0;
rom[79453] = 12'h  0;
rom[79454] = 12'h  0;
rom[79455] = 12'h  0;
rom[79456] = 12'h  0;
rom[79457] = 12'h  0;
rom[79458] = 12'h  0;
rom[79459] = 12'h  0;
rom[79460] = 12'h  0;
rom[79461] = 12'h  0;
rom[79462] = 12'h  0;
rom[79463] = 12'h  0;
rom[79464] = 12'h  0;
rom[79465] = 12'h  0;
rom[79466] = 12'h  0;
rom[79467] = 12'h  0;
rom[79468] = 12'h  0;
rom[79469] = 12'h111;
rom[79470] = 12'h111;
rom[79471] = 12'h111;
rom[79472] = 12'h111;
rom[79473] = 12'h111;
rom[79474] = 12'h222;
rom[79475] = 12'h333;
rom[79476] = 12'h333;
rom[79477] = 12'h333;
rom[79478] = 12'h555;
rom[79479] = 12'h777;
rom[79480] = 12'h999;
rom[79481] = 12'h888;
rom[79482] = 12'h666;
rom[79483] = 12'h444;
rom[79484] = 12'h444;
rom[79485] = 12'h444;
rom[79486] = 12'h333;
rom[79487] = 12'h333;
rom[79488] = 12'h333;
rom[79489] = 12'h333;
rom[79490] = 12'h333;
rom[79491] = 12'h333;
rom[79492] = 12'h444;
rom[79493] = 12'h444;
rom[79494] = 12'h444;
rom[79495] = 12'h444;
rom[79496] = 12'h444;
rom[79497] = 12'h444;
rom[79498] = 12'h555;
rom[79499] = 12'h555;
rom[79500] = 12'h555;
rom[79501] = 12'h666;
rom[79502] = 12'h666;
rom[79503] = 12'h666;
rom[79504] = 12'h777;
rom[79505] = 12'h777;
rom[79506] = 12'h888;
rom[79507] = 12'h888;
rom[79508] = 12'h888;
rom[79509] = 12'h999;
rom[79510] = 12'h999;
rom[79511] = 12'haaa;
rom[79512] = 12'hbbb;
rom[79513] = 12'hccc;
rom[79514] = 12'hddd;
rom[79515] = 12'heee;
rom[79516] = 12'hfff;
rom[79517] = 12'hfff;
rom[79518] = 12'heee;
rom[79519] = 12'hddd;
rom[79520] = 12'hccc;
rom[79521] = 12'hbbb;
rom[79522] = 12'hbbb;
rom[79523] = 12'haaa;
rom[79524] = 12'haaa;
rom[79525] = 12'haaa;
rom[79526] = 12'h999;
rom[79527] = 12'h999;
rom[79528] = 12'h888;
rom[79529] = 12'h888;
rom[79530] = 12'h777;
rom[79531] = 12'h777;
rom[79532] = 12'h777;
rom[79533] = 12'h777;
rom[79534] = 12'h666;
rom[79535] = 12'h666;
rom[79536] = 12'h666;
rom[79537] = 12'h555;
rom[79538] = 12'h555;
rom[79539] = 12'h555;
rom[79540] = 12'h444;
rom[79541] = 12'h444;
rom[79542] = 12'h444;
rom[79543] = 12'h444;
rom[79544] = 12'h444;
rom[79545] = 12'h444;
rom[79546] = 12'h444;
rom[79547] = 12'h444;
rom[79548] = 12'h444;
rom[79549] = 12'h444;
rom[79550] = 12'h444;
rom[79551] = 12'h333;
rom[79552] = 12'h444;
rom[79553] = 12'h333;
rom[79554] = 12'h333;
rom[79555] = 12'h333;
rom[79556] = 12'h333;
rom[79557] = 12'h333;
rom[79558] = 12'h444;
rom[79559] = 12'h444;
rom[79560] = 12'h444;
rom[79561] = 12'h444;
rom[79562] = 12'h444;
rom[79563] = 12'h444;
rom[79564] = 12'h444;
rom[79565] = 12'h444;
rom[79566] = 12'h444;
rom[79567] = 12'h333;
rom[79568] = 12'h333;
rom[79569] = 12'h333;
rom[79570] = 12'h333;
rom[79571] = 12'h333;
rom[79572] = 12'h333;
rom[79573] = 12'h333;
rom[79574] = 12'h333;
rom[79575] = 12'h333;
rom[79576] = 12'h333;
rom[79577] = 12'h333;
rom[79578] = 12'h333;
rom[79579] = 12'h333;
rom[79580] = 12'h333;
rom[79581] = 12'h333;
rom[79582] = 12'h333;
rom[79583] = 12'h333;
rom[79584] = 12'h222;
rom[79585] = 12'h222;
rom[79586] = 12'h222;
rom[79587] = 12'h222;
rom[79588] = 12'h222;
rom[79589] = 12'h222;
rom[79590] = 12'h222;
rom[79591] = 12'h222;
rom[79592] = 12'h222;
rom[79593] = 12'h222;
rom[79594] = 12'h222;
rom[79595] = 12'h333;
rom[79596] = 12'h333;
rom[79597] = 12'h333;
rom[79598] = 12'h333;
rom[79599] = 12'h333;
rom[79600] = 12'hfff;
rom[79601] = 12'hfff;
rom[79602] = 12'hfff;
rom[79603] = 12'hfff;
rom[79604] = 12'hfff;
rom[79605] = 12'hfff;
rom[79606] = 12'hfff;
rom[79607] = 12'hfff;
rom[79608] = 12'hfff;
rom[79609] = 12'hfff;
rom[79610] = 12'hfff;
rom[79611] = 12'hfff;
rom[79612] = 12'hfff;
rom[79613] = 12'hfff;
rom[79614] = 12'hfff;
rom[79615] = 12'hfff;
rom[79616] = 12'hfff;
rom[79617] = 12'hfff;
rom[79618] = 12'hfff;
rom[79619] = 12'hfff;
rom[79620] = 12'hfff;
rom[79621] = 12'hfff;
rom[79622] = 12'hfff;
rom[79623] = 12'hfff;
rom[79624] = 12'hfff;
rom[79625] = 12'hfff;
rom[79626] = 12'hfff;
rom[79627] = 12'hfff;
rom[79628] = 12'hfff;
rom[79629] = 12'hfff;
rom[79630] = 12'hfff;
rom[79631] = 12'hfff;
rom[79632] = 12'hfff;
rom[79633] = 12'hfff;
rom[79634] = 12'hfff;
rom[79635] = 12'hfff;
rom[79636] = 12'hfff;
rom[79637] = 12'hfff;
rom[79638] = 12'hfff;
rom[79639] = 12'hfff;
rom[79640] = 12'hfff;
rom[79641] = 12'hfff;
rom[79642] = 12'hfff;
rom[79643] = 12'hfff;
rom[79644] = 12'hfff;
rom[79645] = 12'hfff;
rom[79646] = 12'hfff;
rom[79647] = 12'hfff;
rom[79648] = 12'hfff;
rom[79649] = 12'hfff;
rom[79650] = 12'hfff;
rom[79651] = 12'hfff;
rom[79652] = 12'hfff;
rom[79653] = 12'hfff;
rom[79654] = 12'hfff;
rom[79655] = 12'hfff;
rom[79656] = 12'hfff;
rom[79657] = 12'hfff;
rom[79658] = 12'hfff;
rom[79659] = 12'hfff;
rom[79660] = 12'hfff;
rom[79661] = 12'hfff;
rom[79662] = 12'hfff;
rom[79663] = 12'hfff;
rom[79664] = 12'hfff;
rom[79665] = 12'hfff;
rom[79666] = 12'hfff;
rom[79667] = 12'hfff;
rom[79668] = 12'hfff;
rom[79669] = 12'hfff;
rom[79670] = 12'hfff;
rom[79671] = 12'hfff;
rom[79672] = 12'hfff;
rom[79673] = 12'hfff;
rom[79674] = 12'hfff;
rom[79675] = 12'hfff;
rom[79676] = 12'hfff;
rom[79677] = 12'hfff;
rom[79678] = 12'hfff;
rom[79679] = 12'hfff;
rom[79680] = 12'hfff;
rom[79681] = 12'hfff;
rom[79682] = 12'hfff;
rom[79683] = 12'hfff;
rom[79684] = 12'hfff;
rom[79685] = 12'hfff;
rom[79686] = 12'hfff;
rom[79687] = 12'hfff;
rom[79688] = 12'hfff;
rom[79689] = 12'hfff;
rom[79690] = 12'hfff;
rom[79691] = 12'hfff;
rom[79692] = 12'hfff;
rom[79693] = 12'hfff;
rom[79694] = 12'hfff;
rom[79695] = 12'hfff;
rom[79696] = 12'hfff;
rom[79697] = 12'hfff;
rom[79698] = 12'hfff;
rom[79699] = 12'hfff;
rom[79700] = 12'hfff;
rom[79701] = 12'hfff;
rom[79702] = 12'hfff;
rom[79703] = 12'hfff;
rom[79704] = 12'hfff;
rom[79705] = 12'hfff;
rom[79706] = 12'hfff;
rom[79707] = 12'hfff;
rom[79708] = 12'hfff;
rom[79709] = 12'hfff;
rom[79710] = 12'hfff;
rom[79711] = 12'hfff;
rom[79712] = 12'hfff;
rom[79713] = 12'hfff;
rom[79714] = 12'hfff;
rom[79715] = 12'hfff;
rom[79716] = 12'hfff;
rom[79717] = 12'hfff;
rom[79718] = 12'hfff;
rom[79719] = 12'hfff;
rom[79720] = 12'hfff;
rom[79721] = 12'hfff;
rom[79722] = 12'heee;
rom[79723] = 12'heee;
rom[79724] = 12'hddd;
rom[79725] = 12'hddd;
rom[79726] = 12'hccc;
rom[79727] = 12'hccc;
rom[79728] = 12'hbbb;
rom[79729] = 12'hbbb;
rom[79730] = 12'hbbb;
rom[79731] = 12'hbbb;
rom[79732] = 12'haaa;
rom[79733] = 12'haaa;
rom[79734] = 12'haaa;
rom[79735] = 12'haaa;
rom[79736] = 12'h999;
rom[79737] = 12'h999;
rom[79738] = 12'haaa;
rom[79739] = 12'haaa;
rom[79740] = 12'h999;
rom[79741] = 12'h999;
rom[79742] = 12'h999;
rom[79743] = 12'h999;
rom[79744] = 12'h888;
rom[79745] = 12'h888;
rom[79746] = 12'h777;
rom[79747] = 12'h777;
rom[79748] = 12'h666;
rom[79749] = 12'h666;
rom[79750] = 12'h555;
rom[79751] = 12'h555;
rom[79752] = 12'h555;
rom[79753] = 12'h444;
rom[79754] = 12'h444;
rom[79755] = 12'h444;
rom[79756] = 12'h444;
rom[79757] = 12'h444;
rom[79758] = 12'h555;
rom[79759] = 12'h555;
rom[79760] = 12'h444;
rom[79761] = 12'h444;
rom[79762] = 12'h444;
rom[79763] = 12'h444;
rom[79764] = 12'h444;
rom[79765] = 12'h444;
rom[79766] = 12'h444;
rom[79767] = 12'h444;
rom[79768] = 12'h444;
rom[79769] = 12'h444;
rom[79770] = 12'h444;
rom[79771] = 12'h555;
rom[79772] = 12'h555;
rom[79773] = 12'h555;
rom[79774] = 12'h555;
rom[79775] = 12'h555;
rom[79776] = 12'h444;
rom[79777] = 12'h444;
rom[79778] = 12'h444;
rom[79779] = 12'h444;
rom[79780] = 12'h444;
rom[79781] = 12'h444;
rom[79782] = 12'h444;
rom[79783] = 12'h444;
rom[79784] = 12'h444;
rom[79785] = 12'h444;
rom[79786] = 12'h444;
rom[79787] = 12'h444;
rom[79788] = 12'h444;
rom[79789] = 12'h444;
rom[79790] = 12'h555;
rom[79791] = 12'h555;
rom[79792] = 12'h555;
rom[79793] = 12'h555;
rom[79794] = 12'h555;
rom[79795] = 12'h555;
rom[79796] = 12'h555;
rom[79797] = 12'h666;
rom[79798] = 12'h666;
rom[79799] = 12'h777;
rom[79800] = 12'h888;
rom[79801] = 12'h999;
rom[79802] = 12'h999;
rom[79803] = 12'h999;
rom[79804] = 12'h999;
rom[79805] = 12'h999;
rom[79806] = 12'h888;
rom[79807] = 12'h777;
rom[79808] = 12'h666;
rom[79809] = 12'h666;
rom[79810] = 12'h555;
rom[79811] = 12'h555;
rom[79812] = 12'h555;
rom[79813] = 12'h444;
rom[79814] = 12'h444;
rom[79815] = 12'h444;
rom[79816] = 12'h444;
rom[79817] = 12'h444;
rom[79818] = 12'h333;
rom[79819] = 12'h333;
rom[79820] = 12'h333;
rom[79821] = 12'h333;
rom[79822] = 12'h333;
rom[79823] = 12'h333;
rom[79824] = 12'h333;
rom[79825] = 12'h333;
rom[79826] = 12'h222;
rom[79827] = 12'h222;
rom[79828] = 12'h222;
rom[79829] = 12'h111;
rom[79830] = 12'h111;
rom[79831] = 12'h111;
rom[79832] = 12'h111;
rom[79833] = 12'h111;
rom[79834] = 12'h111;
rom[79835] = 12'h  0;
rom[79836] = 12'h  0;
rom[79837] = 12'h  0;
rom[79838] = 12'h  0;
rom[79839] = 12'h  0;
rom[79840] = 12'h  0;
rom[79841] = 12'h  0;
rom[79842] = 12'h  0;
rom[79843] = 12'h  0;
rom[79844] = 12'h  0;
rom[79845] = 12'h  0;
rom[79846] = 12'h  0;
rom[79847] = 12'h  0;
rom[79848] = 12'h  0;
rom[79849] = 12'h  0;
rom[79850] = 12'h  0;
rom[79851] = 12'h  0;
rom[79852] = 12'h  0;
rom[79853] = 12'h  0;
rom[79854] = 12'h  0;
rom[79855] = 12'h  0;
rom[79856] = 12'h  0;
rom[79857] = 12'h  0;
rom[79858] = 12'h  0;
rom[79859] = 12'h  0;
rom[79860] = 12'h  0;
rom[79861] = 12'h  0;
rom[79862] = 12'h  0;
rom[79863] = 12'h  0;
rom[79864] = 12'h  0;
rom[79865] = 12'h  0;
rom[79866] = 12'h  0;
rom[79867] = 12'h  0;
rom[79868] = 12'h  0;
rom[79869] = 12'h111;
rom[79870] = 12'h111;
rom[79871] = 12'h111;
rom[79872] = 12'h111;
rom[79873] = 12'h111;
rom[79874] = 12'h222;
rom[79875] = 12'h222;
rom[79876] = 12'h333;
rom[79877] = 12'h333;
rom[79878] = 12'h555;
rom[79879] = 12'h666;
rom[79880] = 12'h999;
rom[79881] = 12'h888;
rom[79882] = 12'h666;
rom[79883] = 12'h444;
rom[79884] = 12'h444;
rom[79885] = 12'h444;
rom[79886] = 12'h333;
rom[79887] = 12'h444;
rom[79888] = 12'h333;
rom[79889] = 12'h333;
rom[79890] = 12'h333;
rom[79891] = 12'h444;
rom[79892] = 12'h444;
rom[79893] = 12'h444;
rom[79894] = 12'h444;
rom[79895] = 12'h444;
rom[79896] = 12'h444;
rom[79897] = 12'h555;
rom[79898] = 12'h555;
rom[79899] = 12'h555;
rom[79900] = 12'h666;
rom[79901] = 12'h666;
rom[79902] = 12'h666;
rom[79903] = 12'h666;
rom[79904] = 12'h777;
rom[79905] = 12'h777;
rom[79906] = 12'h777;
rom[79907] = 12'h888;
rom[79908] = 12'h888;
rom[79909] = 12'h999;
rom[79910] = 12'haaa;
rom[79911] = 12'haaa;
rom[79912] = 12'hccc;
rom[79913] = 12'hddd;
rom[79914] = 12'hddd;
rom[79915] = 12'heee;
rom[79916] = 12'heee;
rom[79917] = 12'heee;
rom[79918] = 12'hddd;
rom[79919] = 12'hccc;
rom[79920] = 12'hbbb;
rom[79921] = 12'hbbb;
rom[79922] = 12'haaa;
rom[79923] = 12'haaa;
rom[79924] = 12'haaa;
rom[79925] = 12'h999;
rom[79926] = 12'h999;
rom[79927] = 12'h999;
rom[79928] = 12'h888;
rom[79929] = 12'h888;
rom[79930] = 12'h777;
rom[79931] = 12'h777;
rom[79932] = 12'h777;
rom[79933] = 12'h777;
rom[79934] = 12'h666;
rom[79935] = 12'h666;
rom[79936] = 12'h666;
rom[79937] = 12'h555;
rom[79938] = 12'h555;
rom[79939] = 12'h555;
rom[79940] = 12'h444;
rom[79941] = 12'h444;
rom[79942] = 12'h444;
rom[79943] = 12'h444;
rom[79944] = 12'h333;
rom[79945] = 12'h333;
rom[79946] = 12'h333;
rom[79947] = 12'h333;
rom[79948] = 12'h333;
rom[79949] = 12'h333;
rom[79950] = 12'h333;
rom[79951] = 12'h333;
rom[79952] = 12'h444;
rom[79953] = 12'h444;
rom[79954] = 12'h333;
rom[79955] = 12'h333;
rom[79956] = 12'h333;
rom[79957] = 12'h333;
rom[79958] = 12'h333;
rom[79959] = 12'h444;
rom[79960] = 12'h444;
rom[79961] = 12'h333;
rom[79962] = 12'h333;
rom[79963] = 12'h444;
rom[79964] = 12'h444;
rom[79965] = 12'h444;
rom[79966] = 12'h444;
rom[79967] = 12'h333;
rom[79968] = 12'h333;
rom[79969] = 12'h333;
rom[79970] = 12'h333;
rom[79971] = 12'h333;
rom[79972] = 12'h333;
rom[79973] = 12'h333;
rom[79974] = 12'h333;
rom[79975] = 12'h333;
rom[79976] = 12'h333;
rom[79977] = 12'h333;
rom[79978] = 12'h333;
rom[79979] = 12'h333;
rom[79980] = 12'h333;
rom[79981] = 12'h333;
rom[79982] = 12'h333;
rom[79983] = 12'h333;
rom[79984] = 12'h222;
rom[79985] = 12'h222;
rom[79986] = 12'h222;
rom[79987] = 12'h222;
rom[79988] = 12'h222;
rom[79989] = 12'h222;
rom[79990] = 12'h222;
rom[79991] = 12'h222;
rom[79992] = 12'h222;
rom[79993] = 12'h222;
rom[79994] = 12'h222;
rom[79995] = 12'h222;
rom[79996] = 12'h222;
rom[79997] = 12'h222;
rom[79998] = 12'h333;
rom[79999] = 12'h333;
rom[80000] = 12'hfff;
rom[80001] = 12'hfff;
rom[80002] = 12'hfff;
rom[80003] = 12'hfff;
rom[80004] = 12'hfff;
rom[80005] = 12'hfff;
rom[80006] = 12'hfff;
rom[80007] = 12'hfff;
rom[80008] = 12'hfff;
rom[80009] = 12'hfff;
rom[80010] = 12'hfff;
rom[80011] = 12'hfff;
rom[80012] = 12'hfff;
rom[80013] = 12'hfff;
rom[80014] = 12'hfff;
rom[80015] = 12'hfff;
rom[80016] = 12'hfff;
rom[80017] = 12'hfff;
rom[80018] = 12'hfff;
rom[80019] = 12'hfff;
rom[80020] = 12'hfff;
rom[80021] = 12'hfff;
rom[80022] = 12'hfff;
rom[80023] = 12'hfff;
rom[80024] = 12'hfff;
rom[80025] = 12'hfff;
rom[80026] = 12'hfff;
rom[80027] = 12'hfff;
rom[80028] = 12'hfff;
rom[80029] = 12'hfff;
rom[80030] = 12'hfff;
rom[80031] = 12'hfff;
rom[80032] = 12'hfff;
rom[80033] = 12'hfff;
rom[80034] = 12'hfff;
rom[80035] = 12'hfff;
rom[80036] = 12'hfff;
rom[80037] = 12'hfff;
rom[80038] = 12'hfff;
rom[80039] = 12'hfff;
rom[80040] = 12'hfff;
rom[80041] = 12'hfff;
rom[80042] = 12'hfff;
rom[80043] = 12'hfff;
rom[80044] = 12'hfff;
rom[80045] = 12'hfff;
rom[80046] = 12'hfff;
rom[80047] = 12'hfff;
rom[80048] = 12'hfff;
rom[80049] = 12'hfff;
rom[80050] = 12'hfff;
rom[80051] = 12'hfff;
rom[80052] = 12'hfff;
rom[80053] = 12'hfff;
rom[80054] = 12'hfff;
rom[80055] = 12'hfff;
rom[80056] = 12'hfff;
rom[80057] = 12'hfff;
rom[80058] = 12'hfff;
rom[80059] = 12'hfff;
rom[80060] = 12'hfff;
rom[80061] = 12'hfff;
rom[80062] = 12'hfff;
rom[80063] = 12'hfff;
rom[80064] = 12'hfff;
rom[80065] = 12'hfff;
rom[80066] = 12'hfff;
rom[80067] = 12'hfff;
rom[80068] = 12'hfff;
rom[80069] = 12'hfff;
rom[80070] = 12'hfff;
rom[80071] = 12'hfff;
rom[80072] = 12'hfff;
rom[80073] = 12'hfff;
rom[80074] = 12'hfff;
rom[80075] = 12'hfff;
rom[80076] = 12'hfff;
rom[80077] = 12'hfff;
rom[80078] = 12'hfff;
rom[80079] = 12'hfff;
rom[80080] = 12'hfff;
rom[80081] = 12'hfff;
rom[80082] = 12'hfff;
rom[80083] = 12'hfff;
rom[80084] = 12'hfff;
rom[80085] = 12'hfff;
rom[80086] = 12'hfff;
rom[80087] = 12'hfff;
rom[80088] = 12'hfff;
rom[80089] = 12'hfff;
rom[80090] = 12'hfff;
rom[80091] = 12'hfff;
rom[80092] = 12'hfff;
rom[80093] = 12'hfff;
rom[80094] = 12'hfff;
rom[80095] = 12'hfff;
rom[80096] = 12'hfff;
rom[80097] = 12'hfff;
rom[80098] = 12'hfff;
rom[80099] = 12'hfff;
rom[80100] = 12'hfff;
rom[80101] = 12'hfff;
rom[80102] = 12'hfff;
rom[80103] = 12'hfff;
rom[80104] = 12'hfff;
rom[80105] = 12'hfff;
rom[80106] = 12'hfff;
rom[80107] = 12'hfff;
rom[80108] = 12'hfff;
rom[80109] = 12'hfff;
rom[80110] = 12'hfff;
rom[80111] = 12'hfff;
rom[80112] = 12'hfff;
rom[80113] = 12'hfff;
rom[80114] = 12'hfff;
rom[80115] = 12'hfff;
rom[80116] = 12'hfff;
rom[80117] = 12'hfff;
rom[80118] = 12'hfff;
rom[80119] = 12'hfff;
rom[80120] = 12'hfff;
rom[80121] = 12'hfff;
rom[80122] = 12'hfff;
rom[80123] = 12'hfff;
rom[80124] = 12'heee;
rom[80125] = 12'heee;
rom[80126] = 12'hddd;
rom[80127] = 12'hddd;
rom[80128] = 12'hccc;
rom[80129] = 12'hccc;
rom[80130] = 12'hbbb;
rom[80131] = 12'hbbb;
rom[80132] = 12'hbbb;
rom[80133] = 12'hbbb;
rom[80134] = 12'hbbb;
rom[80135] = 12'hbbb;
rom[80136] = 12'hbbb;
rom[80137] = 12'hbbb;
rom[80138] = 12'haaa;
rom[80139] = 12'haaa;
rom[80140] = 12'h999;
rom[80141] = 12'h999;
rom[80142] = 12'h999;
rom[80143] = 12'h888;
rom[80144] = 12'h888;
rom[80145] = 12'h777;
rom[80146] = 12'h777;
rom[80147] = 12'h777;
rom[80148] = 12'h666;
rom[80149] = 12'h666;
rom[80150] = 12'h666;
rom[80151] = 12'h555;
rom[80152] = 12'h555;
rom[80153] = 12'h555;
rom[80154] = 12'h444;
rom[80155] = 12'h444;
rom[80156] = 12'h444;
rom[80157] = 12'h555;
rom[80158] = 12'h444;
rom[80159] = 12'h444;
rom[80160] = 12'h555;
rom[80161] = 12'h555;
rom[80162] = 12'h444;
rom[80163] = 12'h444;
rom[80164] = 12'h444;
rom[80165] = 12'h444;
rom[80166] = 12'h444;
rom[80167] = 12'h444;
rom[80168] = 12'h444;
rom[80169] = 12'h444;
rom[80170] = 12'h444;
rom[80171] = 12'h444;
rom[80172] = 12'h444;
rom[80173] = 12'h444;
rom[80174] = 12'h444;
rom[80175] = 12'h444;
rom[80176] = 12'h444;
rom[80177] = 12'h444;
rom[80178] = 12'h444;
rom[80179] = 12'h444;
rom[80180] = 12'h444;
rom[80181] = 12'h444;
rom[80182] = 12'h444;
rom[80183] = 12'h444;
rom[80184] = 12'h444;
rom[80185] = 12'h444;
rom[80186] = 12'h444;
rom[80187] = 12'h444;
rom[80188] = 12'h444;
rom[80189] = 12'h444;
rom[80190] = 12'h444;
rom[80191] = 12'h444;
rom[80192] = 12'h444;
rom[80193] = 12'h444;
rom[80194] = 12'h444;
rom[80195] = 12'h444;
rom[80196] = 12'h444;
rom[80197] = 12'h555;
rom[80198] = 12'h555;
rom[80199] = 12'h666;
rom[80200] = 12'h777;
rom[80201] = 12'h888;
rom[80202] = 12'h888;
rom[80203] = 12'h999;
rom[80204] = 12'haaa;
rom[80205] = 12'haaa;
rom[80206] = 12'h999;
rom[80207] = 12'h888;
rom[80208] = 12'h888;
rom[80209] = 12'h666;
rom[80210] = 12'h555;
rom[80211] = 12'h555;
rom[80212] = 12'h555;
rom[80213] = 12'h555;
rom[80214] = 12'h444;
rom[80215] = 12'h555;
rom[80216] = 12'h444;
rom[80217] = 12'h444;
rom[80218] = 12'h444;
rom[80219] = 12'h444;
rom[80220] = 12'h333;
rom[80221] = 12'h333;
rom[80222] = 12'h333;
rom[80223] = 12'h333;
rom[80224] = 12'h333;
rom[80225] = 12'h222;
rom[80226] = 12'h222;
rom[80227] = 12'h222;
rom[80228] = 12'h222;
rom[80229] = 12'h222;
rom[80230] = 12'h111;
rom[80231] = 12'h111;
rom[80232] = 12'h111;
rom[80233] = 12'h111;
rom[80234] = 12'h111;
rom[80235] = 12'h  0;
rom[80236] = 12'h  0;
rom[80237] = 12'h  0;
rom[80238] = 12'h  0;
rom[80239] = 12'h  0;
rom[80240] = 12'h  0;
rom[80241] = 12'h  0;
rom[80242] = 12'h  0;
rom[80243] = 12'h  0;
rom[80244] = 12'h  0;
rom[80245] = 12'h  0;
rom[80246] = 12'h  0;
rom[80247] = 12'h  0;
rom[80248] = 12'h  0;
rom[80249] = 12'h  0;
rom[80250] = 12'h  0;
rom[80251] = 12'h  0;
rom[80252] = 12'h  0;
rom[80253] = 12'h  0;
rom[80254] = 12'h  0;
rom[80255] = 12'h  0;
rom[80256] = 12'h  0;
rom[80257] = 12'h  0;
rom[80258] = 12'h  0;
rom[80259] = 12'h  0;
rom[80260] = 12'h  0;
rom[80261] = 12'h  0;
rom[80262] = 12'h  0;
rom[80263] = 12'h  0;
rom[80264] = 12'h  0;
rom[80265] = 12'h  0;
rom[80266] = 12'h  0;
rom[80267] = 12'h  0;
rom[80268] = 12'h  0;
rom[80269] = 12'h111;
rom[80270] = 12'h111;
rom[80271] = 12'h111;
rom[80272] = 12'h111;
rom[80273] = 12'h111;
rom[80274] = 12'h222;
rom[80275] = 12'h222;
rom[80276] = 12'h333;
rom[80277] = 12'h333;
rom[80278] = 12'h555;
rom[80279] = 12'h666;
rom[80280] = 12'h999;
rom[80281] = 12'h999;
rom[80282] = 12'h777;
rom[80283] = 12'h555;
rom[80284] = 12'h444;
rom[80285] = 12'h444;
rom[80286] = 12'h444;
rom[80287] = 12'h444;
rom[80288] = 12'h444;
rom[80289] = 12'h444;
rom[80290] = 12'h444;
rom[80291] = 12'h444;
rom[80292] = 12'h444;
rom[80293] = 12'h444;
rom[80294] = 12'h444;
rom[80295] = 12'h444;
rom[80296] = 12'h555;
rom[80297] = 12'h555;
rom[80298] = 12'h555;
rom[80299] = 12'h555;
rom[80300] = 12'h666;
rom[80301] = 12'h666;
rom[80302] = 12'h666;
rom[80303] = 12'h666;
rom[80304] = 12'h777;
rom[80305] = 12'h777;
rom[80306] = 12'h777;
rom[80307] = 12'h888;
rom[80308] = 12'h888;
rom[80309] = 12'h999;
rom[80310] = 12'haaa;
rom[80311] = 12'hbbb;
rom[80312] = 12'hccc;
rom[80313] = 12'hddd;
rom[80314] = 12'heee;
rom[80315] = 12'hddd;
rom[80316] = 12'hddd;
rom[80317] = 12'hccc;
rom[80318] = 12'hbbb;
rom[80319] = 12'haaa;
rom[80320] = 12'haaa;
rom[80321] = 12'haaa;
rom[80322] = 12'haaa;
rom[80323] = 12'h999;
rom[80324] = 12'h999;
rom[80325] = 12'h999;
rom[80326] = 12'h999;
rom[80327] = 12'h888;
rom[80328] = 12'h888;
rom[80329] = 12'h777;
rom[80330] = 12'h777;
rom[80331] = 12'h777;
rom[80332] = 12'h777;
rom[80333] = 12'h666;
rom[80334] = 12'h666;
rom[80335] = 12'h666;
rom[80336] = 12'h666;
rom[80337] = 12'h555;
rom[80338] = 12'h555;
rom[80339] = 12'h555;
rom[80340] = 12'h444;
rom[80341] = 12'h444;
rom[80342] = 12'h444;
rom[80343] = 12'h444;
rom[80344] = 12'h333;
rom[80345] = 12'h333;
rom[80346] = 12'h333;
rom[80347] = 12'h333;
rom[80348] = 12'h333;
rom[80349] = 12'h333;
rom[80350] = 12'h333;
rom[80351] = 12'h333;
rom[80352] = 12'h333;
rom[80353] = 12'h333;
rom[80354] = 12'h333;
rom[80355] = 12'h333;
rom[80356] = 12'h333;
rom[80357] = 12'h333;
rom[80358] = 12'h333;
rom[80359] = 12'h333;
rom[80360] = 12'h444;
rom[80361] = 12'h333;
rom[80362] = 12'h333;
rom[80363] = 12'h333;
rom[80364] = 12'h333;
rom[80365] = 12'h444;
rom[80366] = 12'h444;
rom[80367] = 12'h333;
rom[80368] = 12'h333;
rom[80369] = 12'h333;
rom[80370] = 12'h333;
rom[80371] = 12'h333;
rom[80372] = 12'h333;
rom[80373] = 12'h333;
rom[80374] = 12'h333;
rom[80375] = 12'h333;
rom[80376] = 12'h333;
rom[80377] = 12'h333;
rom[80378] = 12'h333;
rom[80379] = 12'h333;
rom[80380] = 12'h222;
rom[80381] = 12'h222;
rom[80382] = 12'h222;
rom[80383] = 12'h222;
rom[80384] = 12'h222;
rom[80385] = 12'h222;
rom[80386] = 12'h222;
rom[80387] = 12'h222;
rom[80388] = 12'h222;
rom[80389] = 12'h222;
rom[80390] = 12'h222;
rom[80391] = 12'h222;
rom[80392] = 12'h222;
rom[80393] = 12'h222;
rom[80394] = 12'h222;
rom[80395] = 12'h222;
rom[80396] = 12'h222;
rom[80397] = 12'h222;
rom[80398] = 12'h222;
rom[80399] = 12'h222;
rom[80400] = 12'hfff;
rom[80401] = 12'hfff;
rom[80402] = 12'hfff;
rom[80403] = 12'hfff;
rom[80404] = 12'hfff;
rom[80405] = 12'hfff;
rom[80406] = 12'hfff;
rom[80407] = 12'hfff;
rom[80408] = 12'hfff;
rom[80409] = 12'hfff;
rom[80410] = 12'hfff;
rom[80411] = 12'hfff;
rom[80412] = 12'hfff;
rom[80413] = 12'hfff;
rom[80414] = 12'hfff;
rom[80415] = 12'hfff;
rom[80416] = 12'hfff;
rom[80417] = 12'hfff;
rom[80418] = 12'hfff;
rom[80419] = 12'hfff;
rom[80420] = 12'hfff;
rom[80421] = 12'hfff;
rom[80422] = 12'hfff;
rom[80423] = 12'hfff;
rom[80424] = 12'hfff;
rom[80425] = 12'hfff;
rom[80426] = 12'hfff;
rom[80427] = 12'hfff;
rom[80428] = 12'hfff;
rom[80429] = 12'hfff;
rom[80430] = 12'hfff;
rom[80431] = 12'hfff;
rom[80432] = 12'hfff;
rom[80433] = 12'hfff;
rom[80434] = 12'hfff;
rom[80435] = 12'hfff;
rom[80436] = 12'hfff;
rom[80437] = 12'hfff;
rom[80438] = 12'hfff;
rom[80439] = 12'hfff;
rom[80440] = 12'hfff;
rom[80441] = 12'hfff;
rom[80442] = 12'hfff;
rom[80443] = 12'hfff;
rom[80444] = 12'hfff;
rom[80445] = 12'hfff;
rom[80446] = 12'hfff;
rom[80447] = 12'hfff;
rom[80448] = 12'hfff;
rom[80449] = 12'hfff;
rom[80450] = 12'hfff;
rom[80451] = 12'hfff;
rom[80452] = 12'hfff;
rom[80453] = 12'hfff;
rom[80454] = 12'hfff;
rom[80455] = 12'hfff;
rom[80456] = 12'hfff;
rom[80457] = 12'hfff;
rom[80458] = 12'hfff;
rom[80459] = 12'hfff;
rom[80460] = 12'hfff;
rom[80461] = 12'hfff;
rom[80462] = 12'hfff;
rom[80463] = 12'hfff;
rom[80464] = 12'hfff;
rom[80465] = 12'hfff;
rom[80466] = 12'hfff;
rom[80467] = 12'hfff;
rom[80468] = 12'hfff;
rom[80469] = 12'hfff;
rom[80470] = 12'hfff;
rom[80471] = 12'hfff;
rom[80472] = 12'hfff;
rom[80473] = 12'hfff;
rom[80474] = 12'hfff;
rom[80475] = 12'hfff;
rom[80476] = 12'hfff;
rom[80477] = 12'hfff;
rom[80478] = 12'hfff;
rom[80479] = 12'hfff;
rom[80480] = 12'hfff;
rom[80481] = 12'hfff;
rom[80482] = 12'hfff;
rom[80483] = 12'hfff;
rom[80484] = 12'hfff;
rom[80485] = 12'hfff;
rom[80486] = 12'hfff;
rom[80487] = 12'hfff;
rom[80488] = 12'hfff;
rom[80489] = 12'hfff;
rom[80490] = 12'hfff;
rom[80491] = 12'hfff;
rom[80492] = 12'hfff;
rom[80493] = 12'hfff;
rom[80494] = 12'hfff;
rom[80495] = 12'hfff;
rom[80496] = 12'hfff;
rom[80497] = 12'hfff;
rom[80498] = 12'hfff;
rom[80499] = 12'hfff;
rom[80500] = 12'hfff;
rom[80501] = 12'hfff;
rom[80502] = 12'hfff;
rom[80503] = 12'hfff;
rom[80504] = 12'hfff;
rom[80505] = 12'hfff;
rom[80506] = 12'hfff;
rom[80507] = 12'hfff;
rom[80508] = 12'hfff;
rom[80509] = 12'hfff;
rom[80510] = 12'hfff;
rom[80511] = 12'hfff;
rom[80512] = 12'hfff;
rom[80513] = 12'hfff;
rom[80514] = 12'hfff;
rom[80515] = 12'hfff;
rom[80516] = 12'hfff;
rom[80517] = 12'hfff;
rom[80518] = 12'hfff;
rom[80519] = 12'hfff;
rom[80520] = 12'hfff;
rom[80521] = 12'hfff;
rom[80522] = 12'hfff;
rom[80523] = 12'hfff;
rom[80524] = 12'hfff;
rom[80525] = 12'heee;
rom[80526] = 12'heee;
rom[80527] = 12'heee;
rom[80528] = 12'hddd;
rom[80529] = 12'hddd;
rom[80530] = 12'hccc;
rom[80531] = 12'hccc;
rom[80532] = 12'hccc;
rom[80533] = 12'hbbb;
rom[80534] = 12'hbbb;
rom[80535] = 12'hbbb;
rom[80536] = 12'hbbb;
rom[80537] = 12'haaa;
rom[80538] = 12'haaa;
rom[80539] = 12'haaa;
rom[80540] = 12'h999;
rom[80541] = 12'h999;
rom[80542] = 12'h888;
rom[80543] = 12'h888;
rom[80544] = 12'h888;
rom[80545] = 12'h777;
rom[80546] = 12'h777;
rom[80547] = 12'h777;
rom[80548] = 12'h666;
rom[80549] = 12'h666;
rom[80550] = 12'h555;
rom[80551] = 12'h555;
rom[80552] = 12'h555;
rom[80553] = 12'h555;
rom[80554] = 12'h444;
rom[80555] = 12'h444;
rom[80556] = 12'h555;
rom[80557] = 12'h555;
rom[80558] = 12'h444;
rom[80559] = 12'h444;
rom[80560] = 12'h555;
rom[80561] = 12'h444;
rom[80562] = 12'h444;
rom[80563] = 12'h444;
rom[80564] = 12'h444;
rom[80565] = 12'h444;
rom[80566] = 12'h444;
rom[80567] = 12'h444;
rom[80568] = 12'h444;
rom[80569] = 12'h444;
rom[80570] = 12'h444;
rom[80571] = 12'h444;
rom[80572] = 12'h444;
rom[80573] = 12'h444;
rom[80574] = 12'h444;
rom[80575] = 12'h444;
rom[80576] = 12'h444;
rom[80577] = 12'h444;
rom[80578] = 12'h444;
rom[80579] = 12'h444;
rom[80580] = 12'h444;
rom[80581] = 12'h444;
rom[80582] = 12'h444;
rom[80583] = 12'h444;
rom[80584] = 12'h444;
rom[80585] = 12'h444;
rom[80586] = 12'h444;
rom[80587] = 12'h444;
rom[80588] = 12'h444;
rom[80589] = 12'h444;
rom[80590] = 12'h444;
rom[80591] = 12'h444;
rom[80592] = 12'h444;
rom[80593] = 12'h444;
rom[80594] = 12'h444;
rom[80595] = 12'h444;
rom[80596] = 12'h444;
rom[80597] = 12'h555;
rom[80598] = 12'h555;
rom[80599] = 12'h555;
rom[80600] = 12'h666;
rom[80601] = 12'h777;
rom[80602] = 12'h888;
rom[80603] = 12'h999;
rom[80604] = 12'haaa;
rom[80605] = 12'haaa;
rom[80606] = 12'haaa;
rom[80607] = 12'h999;
rom[80608] = 12'h888;
rom[80609] = 12'h666;
rom[80610] = 12'h666;
rom[80611] = 12'h666;
rom[80612] = 12'h555;
rom[80613] = 12'h555;
rom[80614] = 12'h555;
rom[80615] = 12'h555;
rom[80616] = 12'h444;
rom[80617] = 12'h444;
rom[80618] = 12'h444;
rom[80619] = 12'h444;
rom[80620] = 12'h444;
rom[80621] = 12'h333;
rom[80622] = 12'h333;
rom[80623] = 12'h333;
rom[80624] = 12'h333;
rom[80625] = 12'h222;
rom[80626] = 12'h222;
rom[80627] = 12'h222;
rom[80628] = 12'h222;
rom[80629] = 12'h222;
rom[80630] = 12'h111;
rom[80631] = 12'h111;
rom[80632] = 12'h111;
rom[80633] = 12'h111;
rom[80634] = 12'h111;
rom[80635] = 12'h  0;
rom[80636] = 12'h  0;
rom[80637] = 12'h  0;
rom[80638] = 12'h  0;
rom[80639] = 12'h  0;
rom[80640] = 12'h  0;
rom[80641] = 12'h  0;
rom[80642] = 12'h  0;
rom[80643] = 12'h  0;
rom[80644] = 12'h  0;
rom[80645] = 12'h  0;
rom[80646] = 12'h  0;
rom[80647] = 12'h  0;
rom[80648] = 12'h  0;
rom[80649] = 12'h  0;
rom[80650] = 12'h  0;
rom[80651] = 12'h  0;
rom[80652] = 12'h  0;
rom[80653] = 12'h  0;
rom[80654] = 12'h  0;
rom[80655] = 12'h  0;
rom[80656] = 12'h  0;
rom[80657] = 12'h  0;
rom[80658] = 12'h  0;
rom[80659] = 12'h  0;
rom[80660] = 12'h  0;
rom[80661] = 12'h  0;
rom[80662] = 12'h  0;
rom[80663] = 12'h  0;
rom[80664] = 12'h  0;
rom[80665] = 12'h  0;
rom[80666] = 12'h  0;
rom[80667] = 12'h  0;
rom[80668] = 12'h  0;
rom[80669] = 12'h111;
rom[80670] = 12'h111;
rom[80671] = 12'h111;
rom[80672] = 12'h111;
rom[80673] = 12'h111;
rom[80674] = 12'h222;
rom[80675] = 12'h222;
rom[80676] = 12'h333;
rom[80677] = 12'h333;
rom[80678] = 12'h555;
rom[80679] = 12'h666;
rom[80680] = 12'h999;
rom[80681] = 12'h888;
rom[80682] = 12'h777;
rom[80683] = 12'h555;
rom[80684] = 12'h444;
rom[80685] = 12'h444;
rom[80686] = 12'h444;
rom[80687] = 12'h444;
rom[80688] = 12'h444;
rom[80689] = 12'h444;
rom[80690] = 12'h444;
rom[80691] = 12'h444;
rom[80692] = 12'h444;
rom[80693] = 12'h444;
rom[80694] = 12'h444;
rom[80695] = 12'h444;
rom[80696] = 12'h444;
rom[80697] = 12'h555;
rom[80698] = 12'h555;
rom[80699] = 12'h555;
rom[80700] = 12'h666;
rom[80701] = 12'h666;
rom[80702] = 12'h666;
rom[80703] = 12'h666;
rom[80704] = 12'h777;
rom[80705] = 12'h777;
rom[80706] = 12'h777;
rom[80707] = 12'h888;
rom[80708] = 12'h888;
rom[80709] = 12'h999;
rom[80710] = 12'haaa;
rom[80711] = 12'hbbb;
rom[80712] = 12'hddd;
rom[80713] = 12'hddd;
rom[80714] = 12'hddd;
rom[80715] = 12'hddd;
rom[80716] = 12'hccc;
rom[80717] = 12'hccc;
rom[80718] = 12'hbbb;
rom[80719] = 12'haaa;
rom[80720] = 12'h999;
rom[80721] = 12'h999;
rom[80722] = 12'h999;
rom[80723] = 12'h999;
rom[80724] = 12'h999;
rom[80725] = 12'h999;
rom[80726] = 12'h888;
rom[80727] = 12'h888;
rom[80728] = 12'h777;
rom[80729] = 12'h777;
rom[80730] = 12'h777;
rom[80731] = 12'h777;
rom[80732] = 12'h777;
rom[80733] = 12'h666;
rom[80734] = 12'h666;
rom[80735] = 12'h666;
rom[80736] = 12'h666;
rom[80737] = 12'h555;
rom[80738] = 12'h555;
rom[80739] = 12'h444;
rom[80740] = 12'h444;
rom[80741] = 12'h444;
rom[80742] = 12'h444;
rom[80743] = 12'h444;
rom[80744] = 12'h333;
rom[80745] = 12'h333;
rom[80746] = 12'h333;
rom[80747] = 12'h333;
rom[80748] = 12'h333;
rom[80749] = 12'h333;
rom[80750] = 12'h333;
rom[80751] = 12'h333;
rom[80752] = 12'h333;
rom[80753] = 12'h333;
rom[80754] = 12'h333;
rom[80755] = 12'h333;
rom[80756] = 12'h333;
rom[80757] = 12'h333;
rom[80758] = 12'h444;
rom[80759] = 12'h333;
rom[80760] = 12'h444;
rom[80761] = 12'h333;
rom[80762] = 12'h333;
rom[80763] = 12'h333;
rom[80764] = 12'h333;
rom[80765] = 12'h444;
rom[80766] = 12'h333;
rom[80767] = 12'h333;
rom[80768] = 12'h333;
rom[80769] = 12'h333;
rom[80770] = 12'h333;
rom[80771] = 12'h333;
rom[80772] = 12'h333;
rom[80773] = 12'h333;
rom[80774] = 12'h333;
rom[80775] = 12'h333;
rom[80776] = 12'h333;
rom[80777] = 12'h333;
rom[80778] = 12'h333;
rom[80779] = 12'h333;
rom[80780] = 12'h222;
rom[80781] = 12'h222;
rom[80782] = 12'h222;
rom[80783] = 12'h222;
rom[80784] = 12'h222;
rom[80785] = 12'h222;
rom[80786] = 12'h222;
rom[80787] = 12'h222;
rom[80788] = 12'h222;
rom[80789] = 12'h222;
rom[80790] = 12'h222;
rom[80791] = 12'h222;
rom[80792] = 12'h222;
rom[80793] = 12'h222;
rom[80794] = 12'h222;
rom[80795] = 12'h222;
rom[80796] = 12'h222;
rom[80797] = 12'h222;
rom[80798] = 12'h222;
rom[80799] = 12'h222;
rom[80800] = 12'hfff;
rom[80801] = 12'hfff;
rom[80802] = 12'hfff;
rom[80803] = 12'hfff;
rom[80804] = 12'hfff;
rom[80805] = 12'hfff;
rom[80806] = 12'hfff;
rom[80807] = 12'hfff;
rom[80808] = 12'hfff;
rom[80809] = 12'hfff;
rom[80810] = 12'hfff;
rom[80811] = 12'hfff;
rom[80812] = 12'hfff;
rom[80813] = 12'hfff;
rom[80814] = 12'hfff;
rom[80815] = 12'hfff;
rom[80816] = 12'hfff;
rom[80817] = 12'hfff;
rom[80818] = 12'hfff;
rom[80819] = 12'hfff;
rom[80820] = 12'hfff;
rom[80821] = 12'hfff;
rom[80822] = 12'hfff;
rom[80823] = 12'hfff;
rom[80824] = 12'hfff;
rom[80825] = 12'hfff;
rom[80826] = 12'hfff;
rom[80827] = 12'hfff;
rom[80828] = 12'hfff;
rom[80829] = 12'hfff;
rom[80830] = 12'hfff;
rom[80831] = 12'hfff;
rom[80832] = 12'hfff;
rom[80833] = 12'hfff;
rom[80834] = 12'hfff;
rom[80835] = 12'hfff;
rom[80836] = 12'hfff;
rom[80837] = 12'hfff;
rom[80838] = 12'hfff;
rom[80839] = 12'hfff;
rom[80840] = 12'hfff;
rom[80841] = 12'hfff;
rom[80842] = 12'hfff;
rom[80843] = 12'hfff;
rom[80844] = 12'hfff;
rom[80845] = 12'hfff;
rom[80846] = 12'hfff;
rom[80847] = 12'hfff;
rom[80848] = 12'hfff;
rom[80849] = 12'hfff;
rom[80850] = 12'hfff;
rom[80851] = 12'hfff;
rom[80852] = 12'hfff;
rom[80853] = 12'hfff;
rom[80854] = 12'hfff;
rom[80855] = 12'hfff;
rom[80856] = 12'hfff;
rom[80857] = 12'hfff;
rom[80858] = 12'hfff;
rom[80859] = 12'hfff;
rom[80860] = 12'hfff;
rom[80861] = 12'hfff;
rom[80862] = 12'hfff;
rom[80863] = 12'hfff;
rom[80864] = 12'hfff;
rom[80865] = 12'hfff;
rom[80866] = 12'hfff;
rom[80867] = 12'hfff;
rom[80868] = 12'hfff;
rom[80869] = 12'hfff;
rom[80870] = 12'hfff;
rom[80871] = 12'hfff;
rom[80872] = 12'hfff;
rom[80873] = 12'hfff;
rom[80874] = 12'hfff;
rom[80875] = 12'hfff;
rom[80876] = 12'hfff;
rom[80877] = 12'hfff;
rom[80878] = 12'hfff;
rom[80879] = 12'hfff;
rom[80880] = 12'hfff;
rom[80881] = 12'hfff;
rom[80882] = 12'hfff;
rom[80883] = 12'hfff;
rom[80884] = 12'hfff;
rom[80885] = 12'hfff;
rom[80886] = 12'hfff;
rom[80887] = 12'hfff;
rom[80888] = 12'hfff;
rom[80889] = 12'hfff;
rom[80890] = 12'hfff;
rom[80891] = 12'hfff;
rom[80892] = 12'hfff;
rom[80893] = 12'hfff;
rom[80894] = 12'hfff;
rom[80895] = 12'hfff;
rom[80896] = 12'hfff;
rom[80897] = 12'hfff;
rom[80898] = 12'hfff;
rom[80899] = 12'hfff;
rom[80900] = 12'hfff;
rom[80901] = 12'hfff;
rom[80902] = 12'hfff;
rom[80903] = 12'hfff;
rom[80904] = 12'hfff;
rom[80905] = 12'hfff;
rom[80906] = 12'hfff;
rom[80907] = 12'hfff;
rom[80908] = 12'hfff;
rom[80909] = 12'hfff;
rom[80910] = 12'hfff;
rom[80911] = 12'hfff;
rom[80912] = 12'hfff;
rom[80913] = 12'hfff;
rom[80914] = 12'hfff;
rom[80915] = 12'hfff;
rom[80916] = 12'hfff;
rom[80917] = 12'hfff;
rom[80918] = 12'hfff;
rom[80919] = 12'hfff;
rom[80920] = 12'hfff;
rom[80921] = 12'hfff;
rom[80922] = 12'hfff;
rom[80923] = 12'hfff;
rom[80924] = 12'hfff;
rom[80925] = 12'hfff;
rom[80926] = 12'hfff;
rom[80927] = 12'heee;
rom[80928] = 12'heee;
rom[80929] = 12'hddd;
rom[80930] = 12'hddd;
rom[80931] = 12'hddd;
rom[80932] = 12'hccc;
rom[80933] = 12'hccc;
rom[80934] = 12'hbbb;
rom[80935] = 12'hbbb;
rom[80936] = 12'haaa;
rom[80937] = 12'haaa;
rom[80938] = 12'haaa;
rom[80939] = 12'h999;
rom[80940] = 12'h999;
rom[80941] = 12'h999;
rom[80942] = 12'h888;
rom[80943] = 12'h888;
rom[80944] = 12'h888;
rom[80945] = 12'h777;
rom[80946] = 12'h777;
rom[80947] = 12'h777;
rom[80948] = 12'h666;
rom[80949] = 12'h666;
rom[80950] = 12'h555;
rom[80951] = 12'h555;
rom[80952] = 12'h555;
rom[80953] = 12'h555;
rom[80954] = 12'h444;
rom[80955] = 12'h444;
rom[80956] = 12'h555;
rom[80957] = 12'h555;
rom[80958] = 12'h555;
rom[80959] = 12'h444;
rom[80960] = 12'h444;
rom[80961] = 12'h444;
rom[80962] = 12'h444;
rom[80963] = 12'h444;
rom[80964] = 12'h444;
rom[80965] = 12'h444;
rom[80966] = 12'h444;
rom[80967] = 12'h444;
rom[80968] = 12'h333;
rom[80969] = 12'h333;
rom[80970] = 12'h444;
rom[80971] = 12'h444;
rom[80972] = 12'h444;
rom[80973] = 12'h444;
rom[80974] = 12'h444;
rom[80975] = 12'h444;
rom[80976] = 12'h444;
rom[80977] = 12'h444;
rom[80978] = 12'h444;
rom[80979] = 12'h444;
rom[80980] = 12'h444;
rom[80981] = 12'h444;
rom[80982] = 12'h444;
rom[80983] = 12'h444;
rom[80984] = 12'h444;
rom[80985] = 12'h444;
rom[80986] = 12'h444;
rom[80987] = 12'h444;
rom[80988] = 12'h444;
rom[80989] = 12'h444;
rom[80990] = 12'h444;
rom[80991] = 12'h444;
rom[80992] = 12'h444;
rom[80993] = 12'h444;
rom[80994] = 12'h444;
rom[80995] = 12'h444;
rom[80996] = 12'h444;
rom[80997] = 12'h444;
rom[80998] = 12'h444;
rom[80999] = 12'h444;
rom[81000] = 12'h555;
rom[81001] = 12'h555;
rom[81002] = 12'h666;
rom[81003] = 12'h888;
rom[81004] = 12'h999;
rom[81005] = 12'haaa;
rom[81006] = 12'haaa;
rom[81007] = 12'haaa;
rom[81008] = 12'h888;
rom[81009] = 12'h777;
rom[81010] = 12'h666;
rom[81011] = 12'h666;
rom[81012] = 12'h666;
rom[81013] = 12'h555;
rom[81014] = 12'h555;
rom[81015] = 12'h555;
rom[81016] = 12'h555;
rom[81017] = 12'h444;
rom[81018] = 12'h444;
rom[81019] = 12'h444;
rom[81020] = 12'h444;
rom[81021] = 12'h444;
rom[81022] = 12'h333;
rom[81023] = 12'h333;
rom[81024] = 12'h333;
rom[81025] = 12'h333;
rom[81026] = 12'h222;
rom[81027] = 12'h222;
rom[81028] = 12'h222;
rom[81029] = 12'h222;
rom[81030] = 12'h111;
rom[81031] = 12'h111;
rom[81032] = 12'h111;
rom[81033] = 12'h111;
rom[81034] = 12'h111;
rom[81035] = 12'h  0;
rom[81036] = 12'h  0;
rom[81037] = 12'h  0;
rom[81038] = 12'h  0;
rom[81039] = 12'h  0;
rom[81040] = 12'h  0;
rom[81041] = 12'h  0;
rom[81042] = 12'h  0;
rom[81043] = 12'h  0;
rom[81044] = 12'h  0;
rom[81045] = 12'h  0;
rom[81046] = 12'h  0;
rom[81047] = 12'h  0;
rom[81048] = 12'h  0;
rom[81049] = 12'h  0;
rom[81050] = 12'h  0;
rom[81051] = 12'h  0;
rom[81052] = 12'h  0;
rom[81053] = 12'h  0;
rom[81054] = 12'h  0;
rom[81055] = 12'h  0;
rom[81056] = 12'h  0;
rom[81057] = 12'h  0;
rom[81058] = 12'h  0;
rom[81059] = 12'h  0;
rom[81060] = 12'h  0;
rom[81061] = 12'h  0;
rom[81062] = 12'h  0;
rom[81063] = 12'h  0;
rom[81064] = 12'h  0;
rom[81065] = 12'h  0;
rom[81066] = 12'h  0;
rom[81067] = 12'h  0;
rom[81068] = 12'h111;
rom[81069] = 12'h111;
rom[81070] = 12'h111;
rom[81071] = 12'h111;
rom[81072] = 12'h111;
rom[81073] = 12'h111;
rom[81074] = 12'h222;
rom[81075] = 12'h222;
rom[81076] = 12'h333;
rom[81077] = 12'h333;
rom[81078] = 12'h555;
rom[81079] = 12'h666;
rom[81080] = 12'h888;
rom[81081] = 12'h999;
rom[81082] = 12'h777;
rom[81083] = 12'h555;
rom[81084] = 12'h555;
rom[81085] = 12'h555;
rom[81086] = 12'h444;
rom[81087] = 12'h555;
rom[81088] = 12'h444;
rom[81089] = 12'h444;
rom[81090] = 12'h444;
rom[81091] = 12'h444;
rom[81092] = 12'h444;
rom[81093] = 12'h444;
rom[81094] = 12'h555;
rom[81095] = 12'h555;
rom[81096] = 12'h444;
rom[81097] = 12'h555;
rom[81098] = 12'h555;
rom[81099] = 12'h555;
rom[81100] = 12'h666;
rom[81101] = 12'h666;
rom[81102] = 12'h666;
rom[81103] = 12'h666;
rom[81104] = 12'h777;
rom[81105] = 12'h777;
rom[81106] = 12'h888;
rom[81107] = 12'h888;
rom[81108] = 12'h999;
rom[81109] = 12'h999;
rom[81110] = 12'hbbb;
rom[81111] = 12'hccc;
rom[81112] = 12'hddd;
rom[81113] = 12'hddd;
rom[81114] = 12'hddd;
rom[81115] = 12'hccc;
rom[81116] = 12'hbbb;
rom[81117] = 12'haaa;
rom[81118] = 12'h999;
rom[81119] = 12'h999;
rom[81120] = 12'h999;
rom[81121] = 12'h999;
rom[81122] = 12'h999;
rom[81123] = 12'h999;
rom[81124] = 12'h999;
rom[81125] = 12'h999;
rom[81126] = 12'h888;
rom[81127] = 12'h888;
rom[81128] = 12'h777;
rom[81129] = 12'h777;
rom[81130] = 12'h777;
rom[81131] = 12'h777;
rom[81132] = 12'h666;
rom[81133] = 12'h666;
rom[81134] = 12'h666;
rom[81135] = 12'h666;
rom[81136] = 12'h555;
rom[81137] = 12'h555;
rom[81138] = 12'h555;
rom[81139] = 12'h444;
rom[81140] = 12'h444;
rom[81141] = 12'h444;
rom[81142] = 12'h444;
rom[81143] = 12'h333;
rom[81144] = 12'h333;
rom[81145] = 12'h333;
rom[81146] = 12'h333;
rom[81147] = 12'h333;
rom[81148] = 12'h333;
rom[81149] = 12'h333;
rom[81150] = 12'h333;
rom[81151] = 12'h333;
rom[81152] = 12'h333;
rom[81153] = 12'h333;
rom[81154] = 12'h333;
rom[81155] = 12'h333;
rom[81156] = 12'h333;
rom[81157] = 12'h333;
rom[81158] = 12'h444;
rom[81159] = 12'h444;
rom[81160] = 12'h444;
rom[81161] = 12'h333;
rom[81162] = 12'h333;
rom[81163] = 12'h333;
rom[81164] = 12'h333;
rom[81165] = 12'h333;
rom[81166] = 12'h333;
rom[81167] = 12'h333;
rom[81168] = 12'h333;
rom[81169] = 12'h333;
rom[81170] = 12'h333;
rom[81171] = 12'h333;
rom[81172] = 12'h333;
rom[81173] = 12'h333;
rom[81174] = 12'h333;
rom[81175] = 12'h333;
rom[81176] = 12'h333;
rom[81177] = 12'h333;
rom[81178] = 12'h333;
rom[81179] = 12'h333;
rom[81180] = 12'h222;
rom[81181] = 12'h222;
rom[81182] = 12'h222;
rom[81183] = 12'h222;
rom[81184] = 12'h222;
rom[81185] = 12'h222;
rom[81186] = 12'h222;
rom[81187] = 12'h222;
rom[81188] = 12'h222;
rom[81189] = 12'h222;
rom[81190] = 12'h222;
rom[81191] = 12'h222;
rom[81192] = 12'h222;
rom[81193] = 12'h222;
rom[81194] = 12'h222;
rom[81195] = 12'h222;
rom[81196] = 12'h222;
rom[81197] = 12'h222;
rom[81198] = 12'h222;
rom[81199] = 12'h222;
rom[81200] = 12'hfff;
rom[81201] = 12'hfff;
rom[81202] = 12'hfff;
rom[81203] = 12'hfff;
rom[81204] = 12'hfff;
rom[81205] = 12'hfff;
rom[81206] = 12'hfff;
rom[81207] = 12'hfff;
rom[81208] = 12'hfff;
rom[81209] = 12'hfff;
rom[81210] = 12'hfff;
rom[81211] = 12'hfff;
rom[81212] = 12'hfff;
rom[81213] = 12'hfff;
rom[81214] = 12'hfff;
rom[81215] = 12'hfff;
rom[81216] = 12'hfff;
rom[81217] = 12'hfff;
rom[81218] = 12'hfff;
rom[81219] = 12'hfff;
rom[81220] = 12'hfff;
rom[81221] = 12'hfff;
rom[81222] = 12'hfff;
rom[81223] = 12'hfff;
rom[81224] = 12'hfff;
rom[81225] = 12'hfff;
rom[81226] = 12'hfff;
rom[81227] = 12'hfff;
rom[81228] = 12'hfff;
rom[81229] = 12'hfff;
rom[81230] = 12'hfff;
rom[81231] = 12'hfff;
rom[81232] = 12'hfff;
rom[81233] = 12'hfff;
rom[81234] = 12'hfff;
rom[81235] = 12'hfff;
rom[81236] = 12'hfff;
rom[81237] = 12'hfff;
rom[81238] = 12'hfff;
rom[81239] = 12'hfff;
rom[81240] = 12'hfff;
rom[81241] = 12'hfff;
rom[81242] = 12'hfff;
rom[81243] = 12'hfff;
rom[81244] = 12'hfff;
rom[81245] = 12'hfff;
rom[81246] = 12'hfff;
rom[81247] = 12'hfff;
rom[81248] = 12'hfff;
rom[81249] = 12'hfff;
rom[81250] = 12'hfff;
rom[81251] = 12'hfff;
rom[81252] = 12'hfff;
rom[81253] = 12'hfff;
rom[81254] = 12'hfff;
rom[81255] = 12'hfff;
rom[81256] = 12'hfff;
rom[81257] = 12'hfff;
rom[81258] = 12'hfff;
rom[81259] = 12'hfff;
rom[81260] = 12'hfff;
rom[81261] = 12'hfff;
rom[81262] = 12'hfff;
rom[81263] = 12'hfff;
rom[81264] = 12'hfff;
rom[81265] = 12'hfff;
rom[81266] = 12'hfff;
rom[81267] = 12'hfff;
rom[81268] = 12'hfff;
rom[81269] = 12'hfff;
rom[81270] = 12'hfff;
rom[81271] = 12'hfff;
rom[81272] = 12'hfff;
rom[81273] = 12'hfff;
rom[81274] = 12'hfff;
rom[81275] = 12'hfff;
rom[81276] = 12'hfff;
rom[81277] = 12'hfff;
rom[81278] = 12'hfff;
rom[81279] = 12'hfff;
rom[81280] = 12'hfff;
rom[81281] = 12'hfff;
rom[81282] = 12'hfff;
rom[81283] = 12'hfff;
rom[81284] = 12'hfff;
rom[81285] = 12'hfff;
rom[81286] = 12'hfff;
rom[81287] = 12'hfff;
rom[81288] = 12'hfff;
rom[81289] = 12'hfff;
rom[81290] = 12'hfff;
rom[81291] = 12'hfff;
rom[81292] = 12'hfff;
rom[81293] = 12'hfff;
rom[81294] = 12'hfff;
rom[81295] = 12'hfff;
rom[81296] = 12'hfff;
rom[81297] = 12'hfff;
rom[81298] = 12'hfff;
rom[81299] = 12'hfff;
rom[81300] = 12'hfff;
rom[81301] = 12'hfff;
rom[81302] = 12'hfff;
rom[81303] = 12'hfff;
rom[81304] = 12'hfff;
rom[81305] = 12'hfff;
rom[81306] = 12'hfff;
rom[81307] = 12'hfff;
rom[81308] = 12'hfff;
rom[81309] = 12'hfff;
rom[81310] = 12'hfff;
rom[81311] = 12'hfff;
rom[81312] = 12'hfff;
rom[81313] = 12'hfff;
rom[81314] = 12'hfff;
rom[81315] = 12'hfff;
rom[81316] = 12'hfff;
rom[81317] = 12'hfff;
rom[81318] = 12'hfff;
rom[81319] = 12'hfff;
rom[81320] = 12'hfff;
rom[81321] = 12'hfff;
rom[81322] = 12'hfff;
rom[81323] = 12'hfff;
rom[81324] = 12'hfff;
rom[81325] = 12'hfff;
rom[81326] = 12'hfff;
rom[81327] = 12'hfff;
rom[81328] = 12'heee;
rom[81329] = 12'heee;
rom[81330] = 12'heee;
rom[81331] = 12'hddd;
rom[81332] = 12'hddd;
rom[81333] = 12'hccc;
rom[81334] = 12'hccc;
rom[81335] = 12'hbbb;
rom[81336] = 12'hbbb;
rom[81337] = 12'hbbb;
rom[81338] = 12'haaa;
rom[81339] = 12'haaa;
rom[81340] = 12'h999;
rom[81341] = 12'h999;
rom[81342] = 12'h999;
rom[81343] = 12'h888;
rom[81344] = 12'h888;
rom[81345] = 12'h888;
rom[81346] = 12'h777;
rom[81347] = 12'h777;
rom[81348] = 12'h666;
rom[81349] = 12'h666;
rom[81350] = 12'h555;
rom[81351] = 12'h555;
rom[81352] = 12'h555;
rom[81353] = 12'h555;
rom[81354] = 12'h555;
rom[81355] = 12'h555;
rom[81356] = 12'h555;
rom[81357] = 12'h555;
rom[81358] = 12'h555;
rom[81359] = 12'h555;
rom[81360] = 12'h444;
rom[81361] = 12'h444;
rom[81362] = 12'h444;
rom[81363] = 12'h444;
rom[81364] = 12'h444;
rom[81365] = 12'h444;
rom[81366] = 12'h444;
rom[81367] = 12'h444;
rom[81368] = 12'h333;
rom[81369] = 12'h333;
rom[81370] = 12'h333;
rom[81371] = 12'h444;
rom[81372] = 12'h444;
rom[81373] = 12'h444;
rom[81374] = 12'h444;
rom[81375] = 12'h444;
rom[81376] = 12'h444;
rom[81377] = 12'h444;
rom[81378] = 12'h444;
rom[81379] = 12'h444;
rom[81380] = 12'h444;
rom[81381] = 12'h444;
rom[81382] = 12'h444;
rom[81383] = 12'h444;
rom[81384] = 12'h444;
rom[81385] = 12'h444;
rom[81386] = 12'h444;
rom[81387] = 12'h444;
rom[81388] = 12'h444;
rom[81389] = 12'h444;
rom[81390] = 12'h444;
rom[81391] = 12'h444;
rom[81392] = 12'h444;
rom[81393] = 12'h444;
rom[81394] = 12'h444;
rom[81395] = 12'h444;
rom[81396] = 12'h444;
rom[81397] = 12'h444;
rom[81398] = 12'h444;
rom[81399] = 12'h444;
rom[81400] = 12'h444;
rom[81401] = 12'h444;
rom[81402] = 12'h555;
rom[81403] = 12'h666;
rom[81404] = 12'h888;
rom[81405] = 12'h999;
rom[81406] = 12'haaa;
rom[81407] = 12'haaa;
rom[81408] = 12'h999;
rom[81409] = 12'h888;
rom[81410] = 12'h777;
rom[81411] = 12'h666;
rom[81412] = 12'h666;
rom[81413] = 12'h555;
rom[81414] = 12'h555;
rom[81415] = 12'h555;
rom[81416] = 12'h555;
rom[81417] = 12'h444;
rom[81418] = 12'h444;
rom[81419] = 12'h444;
rom[81420] = 12'h444;
rom[81421] = 12'h444;
rom[81422] = 12'h333;
rom[81423] = 12'h333;
rom[81424] = 12'h333;
rom[81425] = 12'h333;
rom[81426] = 12'h222;
rom[81427] = 12'h222;
rom[81428] = 12'h222;
rom[81429] = 12'h222;
rom[81430] = 12'h222;
rom[81431] = 12'h111;
rom[81432] = 12'h111;
rom[81433] = 12'h111;
rom[81434] = 12'h111;
rom[81435] = 12'h111;
rom[81436] = 12'h111;
rom[81437] = 12'h  0;
rom[81438] = 12'h  0;
rom[81439] = 12'h  0;
rom[81440] = 12'h  0;
rom[81441] = 12'h  0;
rom[81442] = 12'h  0;
rom[81443] = 12'h  0;
rom[81444] = 12'h  0;
rom[81445] = 12'h  0;
rom[81446] = 12'h  0;
rom[81447] = 12'h  0;
rom[81448] = 12'h  0;
rom[81449] = 12'h  0;
rom[81450] = 12'h  0;
rom[81451] = 12'h  0;
rom[81452] = 12'h  0;
rom[81453] = 12'h  0;
rom[81454] = 12'h  0;
rom[81455] = 12'h  0;
rom[81456] = 12'h  0;
rom[81457] = 12'h  0;
rom[81458] = 12'h  0;
rom[81459] = 12'h  0;
rom[81460] = 12'h  0;
rom[81461] = 12'h  0;
rom[81462] = 12'h  0;
rom[81463] = 12'h  0;
rom[81464] = 12'h  0;
rom[81465] = 12'h  0;
rom[81466] = 12'h  0;
rom[81467] = 12'h  0;
rom[81468] = 12'h111;
rom[81469] = 12'h111;
rom[81470] = 12'h111;
rom[81471] = 12'h111;
rom[81472] = 12'h111;
rom[81473] = 12'h111;
rom[81474] = 12'h222;
rom[81475] = 12'h222;
rom[81476] = 12'h333;
rom[81477] = 12'h333;
rom[81478] = 12'h555;
rom[81479] = 12'h666;
rom[81480] = 12'h888;
rom[81481] = 12'h999;
rom[81482] = 12'h888;
rom[81483] = 12'h666;
rom[81484] = 12'h555;
rom[81485] = 12'h555;
rom[81486] = 12'h555;
rom[81487] = 12'h555;
rom[81488] = 12'h444;
rom[81489] = 12'h444;
rom[81490] = 12'h444;
rom[81491] = 12'h444;
rom[81492] = 12'h444;
rom[81493] = 12'h555;
rom[81494] = 12'h555;
rom[81495] = 12'h555;
rom[81496] = 12'h555;
rom[81497] = 12'h555;
rom[81498] = 12'h555;
rom[81499] = 12'h666;
rom[81500] = 12'h666;
rom[81501] = 12'h666;
rom[81502] = 12'h666;
rom[81503] = 12'h777;
rom[81504] = 12'h777;
rom[81505] = 12'h777;
rom[81506] = 12'h888;
rom[81507] = 12'h999;
rom[81508] = 12'h999;
rom[81509] = 12'haaa;
rom[81510] = 12'hbbb;
rom[81511] = 12'hccc;
rom[81512] = 12'hddd;
rom[81513] = 12'hddd;
rom[81514] = 12'hccc;
rom[81515] = 12'hbbb;
rom[81516] = 12'haaa;
rom[81517] = 12'h999;
rom[81518] = 12'h999;
rom[81519] = 12'h888;
rom[81520] = 12'h888;
rom[81521] = 12'h999;
rom[81522] = 12'h999;
rom[81523] = 12'h999;
rom[81524] = 12'h999;
rom[81525] = 12'h999;
rom[81526] = 12'h888;
rom[81527] = 12'h888;
rom[81528] = 12'h777;
rom[81529] = 12'h777;
rom[81530] = 12'h777;
rom[81531] = 12'h666;
rom[81532] = 12'h666;
rom[81533] = 12'h666;
rom[81534] = 12'h666;
rom[81535] = 12'h666;
rom[81536] = 12'h555;
rom[81537] = 12'h555;
rom[81538] = 12'h555;
rom[81539] = 12'h444;
rom[81540] = 12'h444;
rom[81541] = 12'h444;
rom[81542] = 12'h333;
rom[81543] = 12'h333;
rom[81544] = 12'h333;
rom[81545] = 12'h333;
rom[81546] = 12'h333;
rom[81547] = 12'h333;
rom[81548] = 12'h333;
rom[81549] = 12'h333;
rom[81550] = 12'h333;
rom[81551] = 12'h333;
rom[81552] = 12'h333;
rom[81553] = 12'h333;
rom[81554] = 12'h333;
rom[81555] = 12'h333;
rom[81556] = 12'h333;
rom[81557] = 12'h444;
rom[81558] = 12'h444;
rom[81559] = 12'h444;
rom[81560] = 12'h333;
rom[81561] = 12'h333;
rom[81562] = 12'h333;
rom[81563] = 12'h333;
rom[81564] = 12'h333;
rom[81565] = 12'h333;
rom[81566] = 12'h333;
rom[81567] = 12'h333;
rom[81568] = 12'h333;
rom[81569] = 12'h333;
rom[81570] = 12'h333;
rom[81571] = 12'h333;
rom[81572] = 12'h333;
rom[81573] = 12'h333;
rom[81574] = 12'h333;
rom[81575] = 12'h333;
rom[81576] = 12'h333;
rom[81577] = 12'h333;
rom[81578] = 12'h333;
rom[81579] = 12'h333;
rom[81580] = 12'h222;
rom[81581] = 12'h222;
rom[81582] = 12'h222;
rom[81583] = 12'h222;
rom[81584] = 12'h222;
rom[81585] = 12'h222;
rom[81586] = 12'h222;
rom[81587] = 12'h222;
rom[81588] = 12'h222;
rom[81589] = 12'h222;
rom[81590] = 12'h222;
rom[81591] = 12'h222;
rom[81592] = 12'h222;
rom[81593] = 12'h222;
rom[81594] = 12'h222;
rom[81595] = 12'h222;
rom[81596] = 12'h222;
rom[81597] = 12'h222;
rom[81598] = 12'h222;
rom[81599] = 12'h222;
rom[81600] = 12'hfff;
rom[81601] = 12'hfff;
rom[81602] = 12'hfff;
rom[81603] = 12'hfff;
rom[81604] = 12'hfff;
rom[81605] = 12'hfff;
rom[81606] = 12'hfff;
rom[81607] = 12'hfff;
rom[81608] = 12'hfff;
rom[81609] = 12'hfff;
rom[81610] = 12'hfff;
rom[81611] = 12'hfff;
rom[81612] = 12'hfff;
rom[81613] = 12'hfff;
rom[81614] = 12'hfff;
rom[81615] = 12'hfff;
rom[81616] = 12'hfff;
rom[81617] = 12'hfff;
rom[81618] = 12'hfff;
rom[81619] = 12'hfff;
rom[81620] = 12'hfff;
rom[81621] = 12'hfff;
rom[81622] = 12'hfff;
rom[81623] = 12'hfff;
rom[81624] = 12'hfff;
rom[81625] = 12'hfff;
rom[81626] = 12'hfff;
rom[81627] = 12'hfff;
rom[81628] = 12'hfff;
rom[81629] = 12'hfff;
rom[81630] = 12'hfff;
rom[81631] = 12'hfff;
rom[81632] = 12'hfff;
rom[81633] = 12'hfff;
rom[81634] = 12'hfff;
rom[81635] = 12'hfff;
rom[81636] = 12'hfff;
rom[81637] = 12'hfff;
rom[81638] = 12'hfff;
rom[81639] = 12'hfff;
rom[81640] = 12'hfff;
rom[81641] = 12'hfff;
rom[81642] = 12'hfff;
rom[81643] = 12'hfff;
rom[81644] = 12'hfff;
rom[81645] = 12'hfff;
rom[81646] = 12'hfff;
rom[81647] = 12'hfff;
rom[81648] = 12'hfff;
rom[81649] = 12'hfff;
rom[81650] = 12'hfff;
rom[81651] = 12'hfff;
rom[81652] = 12'hfff;
rom[81653] = 12'hfff;
rom[81654] = 12'hfff;
rom[81655] = 12'hfff;
rom[81656] = 12'hfff;
rom[81657] = 12'hfff;
rom[81658] = 12'hfff;
rom[81659] = 12'hfff;
rom[81660] = 12'hfff;
rom[81661] = 12'hfff;
rom[81662] = 12'hfff;
rom[81663] = 12'hfff;
rom[81664] = 12'hfff;
rom[81665] = 12'hfff;
rom[81666] = 12'hfff;
rom[81667] = 12'hfff;
rom[81668] = 12'hfff;
rom[81669] = 12'hfff;
rom[81670] = 12'hfff;
rom[81671] = 12'hfff;
rom[81672] = 12'hfff;
rom[81673] = 12'hfff;
rom[81674] = 12'hfff;
rom[81675] = 12'hfff;
rom[81676] = 12'hfff;
rom[81677] = 12'hfff;
rom[81678] = 12'hfff;
rom[81679] = 12'hfff;
rom[81680] = 12'hfff;
rom[81681] = 12'hfff;
rom[81682] = 12'hfff;
rom[81683] = 12'hfff;
rom[81684] = 12'hfff;
rom[81685] = 12'hfff;
rom[81686] = 12'hfff;
rom[81687] = 12'hfff;
rom[81688] = 12'hfff;
rom[81689] = 12'hfff;
rom[81690] = 12'hfff;
rom[81691] = 12'hfff;
rom[81692] = 12'hfff;
rom[81693] = 12'hfff;
rom[81694] = 12'hfff;
rom[81695] = 12'hfff;
rom[81696] = 12'hfff;
rom[81697] = 12'hfff;
rom[81698] = 12'hfff;
rom[81699] = 12'hfff;
rom[81700] = 12'hfff;
rom[81701] = 12'hfff;
rom[81702] = 12'hfff;
rom[81703] = 12'hfff;
rom[81704] = 12'hfff;
rom[81705] = 12'hfff;
rom[81706] = 12'hfff;
rom[81707] = 12'hfff;
rom[81708] = 12'hfff;
rom[81709] = 12'hfff;
rom[81710] = 12'hfff;
rom[81711] = 12'hfff;
rom[81712] = 12'hfff;
rom[81713] = 12'hfff;
rom[81714] = 12'hfff;
rom[81715] = 12'hfff;
rom[81716] = 12'hfff;
rom[81717] = 12'hfff;
rom[81718] = 12'hfff;
rom[81719] = 12'hfff;
rom[81720] = 12'hfff;
rom[81721] = 12'hfff;
rom[81722] = 12'hfff;
rom[81723] = 12'hfff;
rom[81724] = 12'hfff;
rom[81725] = 12'hfff;
rom[81726] = 12'hfff;
rom[81727] = 12'hfff;
rom[81728] = 12'hfff;
rom[81729] = 12'hfff;
rom[81730] = 12'heee;
rom[81731] = 12'heee;
rom[81732] = 12'hddd;
rom[81733] = 12'hddd;
rom[81734] = 12'hccc;
rom[81735] = 12'hccc;
rom[81736] = 12'hbbb;
rom[81737] = 12'hbbb;
rom[81738] = 12'hbbb;
rom[81739] = 12'haaa;
rom[81740] = 12'haaa;
rom[81741] = 12'h999;
rom[81742] = 12'h999;
rom[81743] = 12'h888;
rom[81744] = 12'h888;
rom[81745] = 12'h888;
rom[81746] = 12'h777;
rom[81747] = 12'h777;
rom[81748] = 12'h777;
rom[81749] = 12'h666;
rom[81750] = 12'h666;
rom[81751] = 12'h555;
rom[81752] = 12'h555;
rom[81753] = 12'h555;
rom[81754] = 12'h555;
rom[81755] = 12'h555;
rom[81756] = 12'h555;
rom[81757] = 12'h555;
rom[81758] = 12'h555;
rom[81759] = 12'h555;
rom[81760] = 12'h444;
rom[81761] = 12'h444;
rom[81762] = 12'h444;
rom[81763] = 12'h444;
rom[81764] = 12'h444;
rom[81765] = 12'h444;
rom[81766] = 12'h444;
rom[81767] = 12'h444;
rom[81768] = 12'h333;
rom[81769] = 12'h333;
rom[81770] = 12'h333;
rom[81771] = 12'h333;
rom[81772] = 12'h444;
rom[81773] = 12'h444;
rom[81774] = 12'h444;
rom[81775] = 12'h444;
rom[81776] = 12'h444;
rom[81777] = 12'h444;
rom[81778] = 12'h444;
rom[81779] = 12'h444;
rom[81780] = 12'h444;
rom[81781] = 12'h444;
rom[81782] = 12'h444;
rom[81783] = 12'h444;
rom[81784] = 12'h444;
rom[81785] = 12'h444;
rom[81786] = 12'h444;
rom[81787] = 12'h444;
rom[81788] = 12'h444;
rom[81789] = 12'h444;
rom[81790] = 12'h444;
rom[81791] = 12'h444;
rom[81792] = 12'h444;
rom[81793] = 12'h444;
rom[81794] = 12'h444;
rom[81795] = 12'h444;
rom[81796] = 12'h444;
rom[81797] = 12'h444;
rom[81798] = 12'h444;
rom[81799] = 12'h444;
rom[81800] = 12'h444;
rom[81801] = 12'h444;
rom[81802] = 12'h444;
rom[81803] = 12'h555;
rom[81804] = 12'h777;
rom[81805] = 12'h888;
rom[81806] = 12'haaa;
rom[81807] = 12'haaa;
rom[81808] = 12'haaa;
rom[81809] = 12'h999;
rom[81810] = 12'h888;
rom[81811] = 12'h777;
rom[81812] = 12'h666;
rom[81813] = 12'h555;
rom[81814] = 12'h555;
rom[81815] = 12'h555;
rom[81816] = 12'h555;
rom[81817] = 12'h444;
rom[81818] = 12'h444;
rom[81819] = 12'h444;
rom[81820] = 12'h444;
rom[81821] = 12'h444;
rom[81822] = 12'h333;
rom[81823] = 12'h333;
rom[81824] = 12'h333;
rom[81825] = 12'h222;
rom[81826] = 12'h222;
rom[81827] = 12'h222;
rom[81828] = 12'h222;
rom[81829] = 12'h222;
rom[81830] = 12'h222;
rom[81831] = 12'h111;
rom[81832] = 12'h111;
rom[81833] = 12'h111;
rom[81834] = 12'h111;
rom[81835] = 12'h111;
rom[81836] = 12'h111;
rom[81837] = 12'h111;
rom[81838] = 12'h111;
rom[81839] = 12'h  0;
rom[81840] = 12'h  0;
rom[81841] = 12'h  0;
rom[81842] = 12'h  0;
rom[81843] = 12'h  0;
rom[81844] = 12'h  0;
rom[81845] = 12'h  0;
rom[81846] = 12'h  0;
rom[81847] = 12'h  0;
rom[81848] = 12'h  0;
rom[81849] = 12'h  0;
rom[81850] = 12'h  0;
rom[81851] = 12'h  0;
rom[81852] = 12'h  0;
rom[81853] = 12'h  0;
rom[81854] = 12'h  0;
rom[81855] = 12'h  0;
rom[81856] = 12'h  0;
rom[81857] = 12'h  0;
rom[81858] = 12'h  0;
rom[81859] = 12'h  0;
rom[81860] = 12'h  0;
rom[81861] = 12'h  0;
rom[81862] = 12'h  0;
rom[81863] = 12'h  0;
rom[81864] = 12'h  0;
rom[81865] = 12'h  0;
rom[81866] = 12'h  0;
rom[81867] = 12'h111;
rom[81868] = 12'h111;
rom[81869] = 12'h111;
rom[81870] = 12'h111;
rom[81871] = 12'h111;
rom[81872] = 12'h111;
rom[81873] = 12'h222;
rom[81874] = 12'h222;
rom[81875] = 12'h222;
rom[81876] = 12'h333;
rom[81877] = 12'h333;
rom[81878] = 12'h444;
rom[81879] = 12'h666;
rom[81880] = 12'h888;
rom[81881] = 12'h999;
rom[81882] = 12'h888;
rom[81883] = 12'h666;
rom[81884] = 12'h555;
rom[81885] = 12'h555;
rom[81886] = 12'h555;
rom[81887] = 12'h555;
rom[81888] = 12'h555;
rom[81889] = 12'h555;
rom[81890] = 12'h555;
rom[81891] = 12'h555;
rom[81892] = 12'h555;
rom[81893] = 12'h555;
rom[81894] = 12'h555;
rom[81895] = 12'h555;
rom[81896] = 12'h555;
rom[81897] = 12'h666;
rom[81898] = 12'h666;
rom[81899] = 12'h666;
rom[81900] = 12'h666;
rom[81901] = 12'h666;
rom[81902] = 12'h666;
rom[81903] = 12'h777;
rom[81904] = 12'h777;
rom[81905] = 12'h888;
rom[81906] = 12'h888;
rom[81907] = 12'h999;
rom[81908] = 12'haaa;
rom[81909] = 12'hbbb;
rom[81910] = 12'hccc;
rom[81911] = 12'hddd;
rom[81912] = 12'hccc;
rom[81913] = 12'hccc;
rom[81914] = 12'hbbb;
rom[81915] = 12'haaa;
rom[81916] = 12'h999;
rom[81917] = 12'h999;
rom[81918] = 12'h888;
rom[81919] = 12'h888;
rom[81920] = 12'h888;
rom[81921] = 12'h888;
rom[81922] = 12'h999;
rom[81923] = 12'h999;
rom[81924] = 12'h999;
rom[81925] = 12'h999;
rom[81926] = 12'h888;
rom[81927] = 12'h888;
rom[81928] = 12'h777;
rom[81929] = 12'h777;
rom[81930] = 12'h666;
rom[81931] = 12'h666;
rom[81932] = 12'h666;
rom[81933] = 12'h666;
rom[81934] = 12'h666;
rom[81935] = 12'h555;
rom[81936] = 12'h555;
rom[81937] = 12'h555;
rom[81938] = 12'h555;
rom[81939] = 12'h444;
rom[81940] = 12'h444;
rom[81941] = 12'h444;
rom[81942] = 12'h333;
rom[81943] = 12'h333;
rom[81944] = 12'h333;
rom[81945] = 12'h333;
rom[81946] = 12'h333;
rom[81947] = 12'h333;
rom[81948] = 12'h333;
rom[81949] = 12'h333;
rom[81950] = 12'h333;
rom[81951] = 12'h333;
rom[81952] = 12'h333;
rom[81953] = 12'h333;
rom[81954] = 12'h333;
rom[81955] = 12'h333;
rom[81956] = 12'h333;
rom[81957] = 12'h444;
rom[81958] = 12'h444;
rom[81959] = 12'h444;
rom[81960] = 12'h333;
rom[81961] = 12'h333;
rom[81962] = 12'h333;
rom[81963] = 12'h333;
rom[81964] = 12'h333;
rom[81965] = 12'h333;
rom[81966] = 12'h333;
rom[81967] = 12'h333;
rom[81968] = 12'h333;
rom[81969] = 12'h333;
rom[81970] = 12'h333;
rom[81971] = 12'h333;
rom[81972] = 12'h333;
rom[81973] = 12'h333;
rom[81974] = 12'h333;
rom[81975] = 12'h333;
rom[81976] = 12'h333;
rom[81977] = 12'h333;
rom[81978] = 12'h333;
rom[81979] = 12'h333;
rom[81980] = 12'h222;
rom[81981] = 12'h222;
rom[81982] = 12'h222;
rom[81983] = 12'h222;
rom[81984] = 12'h222;
rom[81985] = 12'h222;
rom[81986] = 12'h222;
rom[81987] = 12'h222;
rom[81988] = 12'h222;
rom[81989] = 12'h222;
rom[81990] = 12'h222;
rom[81991] = 12'h222;
rom[81992] = 12'h222;
rom[81993] = 12'h222;
rom[81994] = 12'h222;
rom[81995] = 12'h222;
rom[81996] = 12'h222;
rom[81997] = 12'h222;
rom[81998] = 12'h222;
rom[81999] = 12'h222;
rom[82000] = 12'hfff;
rom[82001] = 12'hfff;
rom[82002] = 12'hfff;
rom[82003] = 12'hfff;
rom[82004] = 12'hfff;
rom[82005] = 12'hfff;
rom[82006] = 12'hfff;
rom[82007] = 12'hfff;
rom[82008] = 12'hfff;
rom[82009] = 12'hfff;
rom[82010] = 12'hfff;
rom[82011] = 12'hfff;
rom[82012] = 12'hfff;
rom[82013] = 12'hfff;
rom[82014] = 12'hfff;
rom[82015] = 12'hfff;
rom[82016] = 12'hfff;
rom[82017] = 12'hfff;
rom[82018] = 12'hfff;
rom[82019] = 12'hfff;
rom[82020] = 12'hfff;
rom[82021] = 12'hfff;
rom[82022] = 12'hfff;
rom[82023] = 12'hfff;
rom[82024] = 12'hfff;
rom[82025] = 12'hfff;
rom[82026] = 12'hfff;
rom[82027] = 12'hfff;
rom[82028] = 12'hfff;
rom[82029] = 12'hfff;
rom[82030] = 12'hfff;
rom[82031] = 12'hfff;
rom[82032] = 12'hfff;
rom[82033] = 12'hfff;
rom[82034] = 12'hfff;
rom[82035] = 12'hfff;
rom[82036] = 12'hfff;
rom[82037] = 12'hfff;
rom[82038] = 12'hfff;
rom[82039] = 12'hfff;
rom[82040] = 12'hfff;
rom[82041] = 12'hfff;
rom[82042] = 12'hfff;
rom[82043] = 12'hfff;
rom[82044] = 12'hfff;
rom[82045] = 12'hfff;
rom[82046] = 12'hfff;
rom[82047] = 12'hfff;
rom[82048] = 12'hfff;
rom[82049] = 12'hfff;
rom[82050] = 12'hfff;
rom[82051] = 12'hfff;
rom[82052] = 12'hfff;
rom[82053] = 12'hfff;
rom[82054] = 12'hfff;
rom[82055] = 12'hfff;
rom[82056] = 12'hfff;
rom[82057] = 12'hfff;
rom[82058] = 12'hfff;
rom[82059] = 12'hfff;
rom[82060] = 12'hfff;
rom[82061] = 12'hfff;
rom[82062] = 12'hfff;
rom[82063] = 12'hfff;
rom[82064] = 12'hfff;
rom[82065] = 12'hfff;
rom[82066] = 12'hfff;
rom[82067] = 12'hfff;
rom[82068] = 12'hfff;
rom[82069] = 12'hfff;
rom[82070] = 12'hfff;
rom[82071] = 12'hfff;
rom[82072] = 12'hfff;
rom[82073] = 12'hfff;
rom[82074] = 12'hfff;
rom[82075] = 12'hfff;
rom[82076] = 12'hfff;
rom[82077] = 12'hfff;
rom[82078] = 12'hfff;
rom[82079] = 12'hfff;
rom[82080] = 12'hfff;
rom[82081] = 12'hfff;
rom[82082] = 12'hfff;
rom[82083] = 12'hfff;
rom[82084] = 12'hfff;
rom[82085] = 12'hfff;
rom[82086] = 12'hfff;
rom[82087] = 12'hfff;
rom[82088] = 12'hfff;
rom[82089] = 12'hfff;
rom[82090] = 12'hfff;
rom[82091] = 12'hfff;
rom[82092] = 12'hfff;
rom[82093] = 12'hfff;
rom[82094] = 12'hfff;
rom[82095] = 12'hfff;
rom[82096] = 12'hfff;
rom[82097] = 12'hfff;
rom[82098] = 12'hfff;
rom[82099] = 12'hfff;
rom[82100] = 12'hfff;
rom[82101] = 12'hfff;
rom[82102] = 12'hfff;
rom[82103] = 12'hfff;
rom[82104] = 12'hfff;
rom[82105] = 12'hfff;
rom[82106] = 12'hfff;
rom[82107] = 12'hfff;
rom[82108] = 12'hfff;
rom[82109] = 12'hfff;
rom[82110] = 12'hfff;
rom[82111] = 12'hfff;
rom[82112] = 12'hfff;
rom[82113] = 12'hfff;
rom[82114] = 12'hfff;
rom[82115] = 12'hfff;
rom[82116] = 12'hfff;
rom[82117] = 12'hfff;
rom[82118] = 12'hfff;
rom[82119] = 12'hfff;
rom[82120] = 12'hfff;
rom[82121] = 12'hfff;
rom[82122] = 12'hfff;
rom[82123] = 12'hfff;
rom[82124] = 12'hfff;
rom[82125] = 12'hfff;
rom[82126] = 12'hfff;
rom[82127] = 12'hfff;
rom[82128] = 12'hfff;
rom[82129] = 12'hfff;
rom[82130] = 12'hfff;
rom[82131] = 12'heee;
rom[82132] = 12'heee;
rom[82133] = 12'heee;
rom[82134] = 12'hddd;
rom[82135] = 12'hddd;
rom[82136] = 12'hccc;
rom[82137] = 12'hccc;
rom[82138] = 12'hbbb;
rom[82139] = 12'hbbb;
rom[82140] = 12'haaa;
rom[82141] = 12'haaa;
rom[82142] = 12'h999;
rom[82143] = 12'h999;
rom[82144] = 12'h999;
rom[82145] = 12'h888;
rom[82146] = 12'h888;
rom[82147] = 12'h777;
rom[82148] = 12'h777;
rom[82149] = 12'h666;
rom[82150] = 12'h666;
rom[82151] = 12'h555;
rom[82152] = 12'h666;
rom[82153] = 12'h555;
rom[82154] = 12'h555;
rom[82155] = 12'h555;
rom[82156] = 12'h555;
rom[82157] = 12'h555;
rom[82158] = 12'h555;
rom[82159] = 12'h555;
rom[82160] = 12'h444;
rom[82161] = 12'h444;
rom[82162] = 12'h444;
rom[82163] = 12'h444;
rom[82164] = 12'h444;
rom[82165] = 12'h444;
rom[82166] = 12'h444;
rom[82167] = 12'h444;
rom[82168] = 12'h333;
rom[82169] = 12'h333;
rom[82170] = 12'h333;
rom[82171] = 12'h333;
rom[82172] = 12'h444;
rom[82173] = 12'h444;
rom[82174] = 12'h444;
rom[82175] = 12'h444;
rom[82176] = 12'h444;
rom[82177] = 12'h444;
rom[82178] = 12'h444;
rom[82179] = 12'h444;
rom[82180] = 12'h444;
rom[82181] = 12'h444;
rom[82182] = 12'h444;
rom[82183] = 12'h444;
rom[82184] = 12'h444;
rom[82185] = 12'h444;
rom[82186] = 12'h444;
rom[82187] = 12'h444;
rom[82188] = 12'h444;
rom[82189] = 12'h444;
rom[82190] = 12'h444;
rom[82191] = 12'h444;
rom[82192] = 12'h444;
rom[82193] = 12'h444;
rom[82194] = 12'h444;
rom[82195] = 12'h444;
rom[82196] = 12'h444;
rom[82197] = 12'h444;
rom[82198] = 12'h333;
rom[82199] = 12'h333;
rom[82200] = 12'h444;
rom[82201] = 12'h444;
rom[82202] = 12'h444;
rom[82203] = 12'h444;
rom[82204] = 12'h555;
rom[82205] = 12'h777;
rom[82206] = 12'h888;
rom[82207] = 12'haaa;
rom[82208] = 12'haaa;
rom[82209] = 12'haaa;
rom[82210] = 12'h888;
rom[82211] = 12'h777;
rom[82212] = 12'h666;
rom[82213] = 12'h555;
rom[82214] = 12'h555;
rom[82215] = 12'h555;
rom[82216] = 12'h555;
rom[82217] = 12'h555;
rom[82218] = 12'h444;
rom[82219] = 12'h444;
rom[82220] = 12'h444;
rom[82221] = 12'h444;
rom[82222] = 12'h333;
rom[82223] = 12'h333;
rom[82224] = 12'h333;
rom[82225] = 12'h222;
rom[82226] = 12'h222;
rom[82227] = 12'h222;
rom[82228] = 12'h222;
rom[82229] = 12'h222;
rom[82230] = 12'h111;
rom[82231] = 12'h111;
rom[82232] = 12'h111;
rom[82233] = 12'h111;
rom[82234] = 12'h111;
rom[82235] = 12'h111;
rom[82236] = 12'h111;
rom[82237] = 12'h111;
rom[82238] = 12'h111;
rom[82239] = 12'h111;
rom[82240] = 12'h  0;
rom[82241] = 12'h  0;
rom[82242] = 12'h  0;
rom[82243] = 12'h  0;
rom[82244] = 12'h  0;
rom[82245] = 12'h  0;
rom[82246] = 12'h  0;
rom[82247] = 12'h  0;
rom[82248] = 12'h  0;
rom[82249] = 12'h  0;
rom[82250] = 12'h  0;
rom[82251] = 12'h  0;
rom[82252] = 12'h  0;
rom[82253] = 12'h  0;
rom[82254] = 12'h  0;
rom[82255] = 12'h  0;
rom[82256] = 12'h  0;
rom[82257] = 12'h  0;
rom[82258] = 12'h  0;
rom[82259] = 12'h  0;
rom[82260] = 12'h  0;
rom[82261] = 12'h  0;
rom[82262] = 12'h  0;
rom[82263] = 12'h  0;
rom[82264] = 12'h  0;
rom[82265] = 12'h  0;
rom[82266] = 12'h  0;
rom[82267] = 12'h111;
rom[82268] = 12'h111;
rom[82269] = 12'h111;
rom[82270] = 12'h111;
rom[82271] = 12'h111;
rom[82272] = 12'h222;
rom[82273] = 12'h222;
rom[82274] = 12'h222;
rom[82275] = 12'h222;
rom[82276] = 12'h333;
rom[82277] = 12'h333;
rom[82278] = 12'h444;
rom[82279] = 12'h555;
rom[82280] = 12'h888;
rom[82281] = 12'haaa;
rom[82282] = 12'h999;
rom[82283] = 12'h777;
rom[82284] = 12'h666;
rom[82285] = 12'h555;
rom[82286] = 12'h555;
rom[82287] = 12'h555;
rom[82288] = 12'h555;
rom[82289] = 12'h555;
rom[82290] = 12'h555;
rom[82291] = 12'h555;
rom[82292] = 12'h555;
rom[82293] = 12'h555;
rom[82294] = 12'h555;
rom[82295] = 12'h555;
rom[82296] = 12'h555;
rom[82297] = 12'h666;
rom[82298] = 12'h666;
rom[82299] = 12'h666;
rom[82300] = 12'h666;
rom[82301] = 12'h666;
rom[82302] = 12'h666;
rom[82303] = 12'h777;
rom[82304] = 12'h777;
rom[82305] = 12'h888;
rom[82306] = 12'h999;
rom[82307] = 12'h999;
rom[82308] = 12'haaa;
rom[82309] = 12'hbbb;
rom[82310] = 12'hccc;
rom[82311] = 12'hccc;
rom[82312] = 12'hccc;
rom[82313] = 12'hbbb;
rom[82314] = 12'haaa;
rom[82315] = 12'h999;
rom[82316] = 12'h999;
rom[82317] = 12'h999;
rom[82318] = 12'h888;
rom[82319] = 12'h888;
rom[82320] = 12'h888;
rom[82321] = 12'h888;
rom[82322] = 12'h888;
rom[82323] = 12'h888;
rom[82324] = 12'h888;
rom[82325] = 12'h888;
rom[82326] = 12'h888;
rom[82327] = 12'h777;
rom[82328] = 12'h777;
rom[82329] = 12'h777;
rom[82330] = 12'h666;
rom[82331] = 12'h666;
rom[82332] = 12'h666;
rom[82333] = 12'h666;
rom[82334] = 12'h666;
rom[82335] = 12'h555;
rom[82336] = 12'h555;
rom[82337] = 12'h555;
rom[82338] = 12'h555;
rom[82339] = 12'h444;
rom[82340] = 12'h444;
rom[82341] = 12'h444;
rom[82342] = 12'h333;
rom[82343] = 12'h333;
rom[82344] = 12'h333;
rom[82345] = 12'h333;
rom[82346] = 12'h333;
rom[82347] = 12'h333;
rom[82348] = 12'h333;
rom[82349] = 12'h333;
rom[82350] = 12'h333;
rom[82351] = 12'h333;
rom[82352] = 12'h333;
rom[82353] = 12'h333;
rom[82354] = 12'h333;
rom[82355] = 12'h333;
rom[82356] = 12'h333;
rom[82357] = 12'h444;
rom[82358] = 12'h444;
rom[82359] = 12'h444;
rom[82360] = 12'h444;
rom[82361] = 12'h333;
rom[82362] = 12'h333;
rom[82363] = 12'h333;
rom[82364] = 12'h333;
rom[82365] = 12'h333;
rom[82366] = 12'h333;
rom[82367] = 12'h333;
rom[82368] = 12'h333;
rom[82369] = 12'h333;
rom[82370] = 12'h333;
rom[82371] = 12'h333;
rom[82372] = 12'h333;
rom[82373] = 12'h333;
rom[82374] = 12'h333;
rom[82375] = 12'h333;
rom[82376] = 12'h333;
rom[82377] = 12'h333;
rom[82378] = 12'h333;
rom[82379] = 12'h333;
rom[82380] = 12'h222;
rom[82381] = 12'h222;
rom[82382] = 12'h222;
rom[82383] = 12'h222;
rom[82384] = 12'h222;
rom[82385] = 12'h222;
rom[82386] = 12'h222;
rom[82387] = 12'h222;
rom[82388] = 12'h222;
rom[82389] = 12'h222;
rom[82390] = 12'h222;
rom[82391] = 12'h222;
rom[82392] = 12'h222;
rom[82393] = 12'h222;
rom[82394] = 12'h222;
rom[82395] = 12'h222;
rom[82396] = 12'h222;
rom[82397] = 12'h222;
rom[82398] = 12'h222;
rom[82399] = 12'h222;
rom[82400] = 12'hfff;
rom[82401] = 12'hfff;
rom[82402] = 12'hfff;
rom[82403] = 12'hfff;
rom[82404] = 12'hfff;
rom[82405] = 12'hfff;
rom[82406] = 12'hfff;
rom[82407] = 12'hfff;
rom[82408] = 12'hfff;
rom[82409] = 12'hfff;
rom[82410] = 12'hfff;
rom[82411] = 12'hfff;
rom[82412] = 12'hfff;
rom[82413] = 12'hfff;
rom[82414] = 12'hfff;
rom[82415] = 12'hfff;
rom[82416] = 12'hfff;
rom[82417] = 12'hfff;
rom[82418] = 12'hfff;
rom[82419] = 12'hfff;
rom[82420] = 12'hfff;
rom[82421] = 12'hfff;
rom[82422] = 12'hfff;
rom[82423] = 12'hfff;
rom[82424] = 12'hfff;
rom[82425] = 12'hfff;
rom[82426] = 12'hfff;
rom[82427] = 12'hfff;
rom[82428] = 12'hfff;
rom[82429] = 12'hfff;
rom[82430] = 12'hfff;
rom[82431] = 12'hfff;
rom[82432] = 12'hfff;
rom[82433] = 12'hfff;
rom[82434] = 12'hfff;
rom[82435] = 12'hfff;
rom[82436] = 12'hfff;
rom[82437] = 12'hfff;
rom[82438] = 12'hfff;
rom[82439] = 12'hfff;
rom[82440] = 12'hfff;
rom[82441] = 12'hfff;
rom[82442] = 12'hfff;
rom[82443] = 12'hfff;
rom[82444] = 12'hfff;
rom[82445] = 12'hfff;
rom[82446] = 12'hfff;
rom[82447] = 12'hfff;
rom[82448] = 12'hfff;
rom[82449] = 12'hfff;
rom[82450] = 12'hfff;
rom[82451] = 12'hfff;
rom[82452] = 12'hfff;
rom[82453] = 12'hfff;
rom[82454] = 12'hfff;
rom[82455] = 12'hfff;
rom[82456] = 12'hfff;
rom[82457] = 12'hfff;
rom[82458] = 12'hfff;
rom[82459] = 12'hfff;
rom[82460] = 12'hfff;
rom[82461] = 12'hfff;
rom[82462] = 12'hfff;
rom[82463] = 12'hfff;
rom[82464] = 12'hfff;
rom[82465] = 12'hfff;
rom[82466] = 12'hfff;
rom[82467] = 12'hfff;
rom[82468] = 12'hfff;
rom[82469] = 12'hfff;
rom[82470] = 12'hfff;
rom[82471] = 12'hfff;
rom[82472] = 12'hfff;
rom[82473] = 12'hfff;
rom[82474] = 12'hfff;
rom[82475] = 12'hfff;
rom[82476] = 12'hfff;
rom[82477] = 12'hfff;
rom[82478] = 12'hfff;
rom[82479] = 12'hfff;
rom[82480] = 12'hfff;
rom[82481] = 12'hfff;
rom[82482] = 12'hfff;
rom[82483] = 12'hfff;
rom[82484] = 12'hfff;
rom[82485] = 12'hfff;
rom[82486] = 12'hfff;
rom[82487] = 12'hfff;
rom[82488] = 12'hfff;
rom[82489] = 12'hfff;
rom[82490] = 12'hfff;
rom[82491] = 12'hfff;
rom[82492] = 12'hfff;
rom[82493] = 12'hfff;
rom[82494] = 12'hfff;
rom[82495] = 12'hfff;
rom[82496] = 12'hfff;
rom[82497] = 12'hfff;
rom[82498] = 12'hfff;
rom[82499] = 12'hfff;
rom[82500] = 12'hfff;
rom[82501] = 12'hfff;
rom[82502] = 12'hfff;
rom[82503] = 12'hfff;
rom[82504] = 12'hfff;
rom[82505] = 12'hfff;
rom[82506] = 12'hfff;
rom[82507] = 12'hfff;
rom[82508] = 12'hfff;
rom[82509] = 12'hfff;
rom[82510] = 12'hfff;
rom[82511] = 12'hfff;
rom[82512] = 12'hfff;
rom[82513] = 12'hfff;
rom[82514] = 12'hfff;
rom[82515] = 12'hfff;
rom[82516] = 12'hfff;
rom[82517] = 12'hfff;
rom[82518] = 12'hfff;
rom[82519] = 12'hfff;
rom[82520] = 12'hfff;
rom[82521] = 12'hfff;
rom[82522] = 12'hfff;
rom[82523] = 12'hfff;
rom[82524] = 12'hfff;
rom[82525] = 12'hfff;
rom[82526] = 12'hfff;
rom[82527] = 12'hfff;
rom[82528] = 12'hfff;
rom[82529] = 12'hfff;
rom[82530] = 12'hfff;
rom[82531] = 12'hfff;
rom[82532] = 12'hfff;
rom[82533] = 12'heee;
rom[82534] = 12'heee;
rom[82535] = 12'heee;
rom[82536] = 12'hddd;
rom[82537] = 12'hddd;
rom[82538] = 12'hccc;
rom[82539] = 12'hccc;
rom[82540] = 12'hbbb;
rom[82541] = 12'haaa;
rom[82542] = 12'haaa;
rom[82543] = 12'haaa;
rom[82544] = 12'h999;
rom[82545] = 12'h999;
rom[82546] = 12'h888;
rom[82547] = 12'h888;
rom[82548] = 12'h777;
rom[82549] = 12'h777;
rom[82550] = 12'h666;
rom[82551] = 12'h666;
rom[82552] = 12'h666;
rom[82553] = 12'h666;
rom[82554] = 12'h555;
rom[82555] = 12'h555;
rom[82556] = 12'h555;
rom[82557] = 12'h555;
rom[82558] = 12'h555;
rom[82559] = 12'h555;
rom[82560] = 12'h555;
rom[82561] = 12'h444;
rom[82562] = 12'h444;
rom[82563] = 12'h444;
rom[82564] = 12'h444;
rom[82565] = 12'h444;
rom[82566] = 12'h444;
rom[82567] = 12'h444;
rom[82568] = 12'h333;
rom[82569] = 12'h333;
rom[82570] = 12'h333;
rom[82571] = 12'h333;
rom[82572] = 12'h333;
rom[82573] = 12'h333;
rom[82574] = 12'h444;
rom[82575] = 12'h444;
rom[82576] = 12'h444;
rom[82577] = 12'h444;
rom[82578] = 12'h444;
rom[82579] = 12'h444;
rom[82580] = 12'h444;
rom[82581] = 12'h444;
rom[82582] = 12'h444;
rom[82583] = 12'h444;
rom[82584] = 12'h444;
rom[82585] = 12'h444;
rom[82586] = 12'h444;
rom[82587] = 12'h444;
rom[82588] = 12'h444;
rom[82589] = 12'h444;
rom[82590] = 12'h555;
rom[82591] = 12'h444;
rom[82592] = 12'h444;
rom[82593] = 12'h444;
rom[82594] = 12'h444;
rom[82595] = 12'h444;
rom[82596] = 12'h444;
rom[82597] = 12'h333;
rom[82598] = 12'h333;
rom[82599] = 12'h333;
rom[82600] = 12'h444;
rom[82601] = 12'h333;
rom[82602] = 12'h333;
rom[82603] = 12'h444;
rom[82604] = 12'h444;
rom[82605] = 12'h555;
rom[82606] = 12'h777;
rom[82607] = 12'h999;
rom[82608] = 12'haaa;
rom[82609] = 12'haaa;
rom[82610] = 12'h999;
rom[82611] = 12'h888;
rom[82612] = 12'h777;
rom[82613] = 12'h666;
rom[82614] = 12'h555;
rom[82615] = 12'h555;
rom[82616] = 12'h444;
rom[82617] = 12'h444;
rom[82618] = 12'h444;
rom[82619] = 12'h444;
rom[82620] = 12'h333;
rom[82621] = 12'h333;
rom[82622] = 12'h333;
rom[82623] = 12'h333;
rom[82624] = 12'h222;
rom[82625] = 12'h222;
rom[82626] = 12'h222;
rom[82627] = 12'h222;
rom[82628] = 12'h222;
rom[82629] = 12'h222;
rom[82630] = 12'h111;
rom[82631] = 12'h111;
rom[82632] = 12'h111;
rom[82633] = 12'h111;
rom[82634] = 12'h111;
rom[82635] = 12'h111;
rom[82636] = 12'h111;
rom[82637] = 12'h111;
rom[82638] = 12'h111;
rom[82639] = 12'h111;
rom[82640] = 12'h111;
rom[82641] = 12'h111;
rom[82642] = 12'h  0;
rom[82643] = 12'h  0;
rom[82644] = 12'h  0;
rom[82645] = 12'h  0;
rom[82646] = 12'h  0;
rom[82647] = 12'h  0;
rom[82648] = 12'h  0;
rom[82649] = 12'h  0;
rom[82650] = 12'h  0;
rom[82651] = 12'h  0;
rom[82652] = 12'h  0;
rom[82653] = 12'h  0;
rom[82654] = 12'h  0;
rom[82655] = 12'h  0;
rom[82656] = 12'h  0;
rom[82657] = 12'h  0;
rom[82658] = 12'h  0;
rom[82659] = 12'h  0;
rom[82660] = 12'h  0;
rom[82661] = 12'h  0;
rom[82662] = 12'h  0;
rom[82663] = 12'h  0;
rom[82664] = 12'h  0;
rom[82665] = 12'h  0;
rom[82666] = 12'h111;
rom[82667] = 12'h111;
rom[82668] = 12'h111;
rom[82669] = 12'h111;
rom[82670] = 12'h111;
rom[82671] = 12'h111;
rom[82672] = 12'h222;
rom[82673] = 12'h222;
rom[82674] = 12'h222;
rom[82675] = 12'h333;
rom[82676] = 12'h333;
rom[82677] = 12'h333;
rom[82678] = 12'h444;
rom[82679] = 12'h555;
rom[82680] = 12'h888;
rom[82681] = 12'haaa;
rom[82682] = 12'h999;
rom[82683] = 12'h777;
rom[82684] = 12'h666;
rom[82685] = 12'h666;
rom[82686] = 12'h555;
rom[82687] = 12'h555;
rom[82688] = 12'h555;
rom[82689] = 12'h555;
rom[82690] = 12'h555;
rom[82691] = 12'h555;
rom[82692] = 12'h555;
rom[82693] = 12'h555;
rom[82694] = 12'h555;
rom[82695] = 12'h555;
rom[82696] = 12'h555;
rom[82697] = 12'h666;
rom[82698] = 12'h666;
rom[82699] = 12'h666;
rom[82700] = 12'h666;
rom[82701] = 12'h666;
rom[82702] = 12'h777;
rom[82703] = 12'h777;
rom[82704] = 12'h888;
rom[82705] = 12'h888;
rom[82706] = 12'h999;
rom[82707] = 12'h999;
rom[82708] = 12'hbbb;
rom[82709] = 12'hccc;
rom[82710] = 12'hccc;
rom[82711] = 12'hbbb;
rom[82712] = 12'hbbb;
rom[82713] = 12'haaa;
rom[82714] = 12'h999;
rom[82715] = 12'h999;
rom[82716] = 12'h888;
rom[82717] = 12'h888;
rom[82718] = 12'h888;
rom[82719] = 12'h888;
rom[82720] = 12'h888;
rom[82721] = 12'h888;
rom[82722] = 12'h888;
rom[82723] = 12'h888;
rom[82724] = 12'h888;
rom[82725] = 12'h888;
rom[82726] = 12'h888;
rom[82727] = 12'h777;
rom[82728] = 12'h777;
rom[82729] = 12'h777;
rom[82730] = 12'h666;
rom[82731] = 12'h666;
rom[82732] = 12'h666;
rom[82733] = 12'h666;
rom[82734] = 12'h666;
rom[82735] = 12'h555;
rom[82736] = 12'h666;
rom[82737] = 12'h555;
rom[82738] = 12'h555;
rom[82739] = 12'h444;
rom[82740] = 12'h444;
rom[82741] = 12'h444;
rom[82742] = 12'h444;
rom[82743] = 12'h333;
rom[82744] = 12'h333;
rom[82745] = 12'h333;
rom[82746] = 12'h333;
rom[82747] = 12'h333;
rom[82748] = 12'h333;
rom[82749] = 12'h333;
rom[82750] = 12'h333;
rom[82751] = 12'h333;
rom[82752] = 12'h333;
rom[82753] = 12'h333;
rom[82754] = 12'h333;
rom[82755] = 12'h333;
rom[82756] = 12'h444;
rom[82757] = 12'h444;
rom[82758] = 12'h444;
rom[82759] = 12'h444;
rom[82760] = 12'h444;
rom[82761] = 12'h333;
rom[82762] = 12'h333;
rom[82763] = 12'h333;
rom[82764] = 12'h333;
rom[82765] = 12'h444;
rom[82766] = 12'h333;
rom[82767] = 12'h333;
rom[82768] = 12'h333;
rom[82769] = 12'h333;
rom[82770] = 12'h333;
rom[82771] = 12'h333;
rom[82772] = 12'h333;
rom[82773] = 12'h333;
rom[82774] = 12'h333;
rom[82775] = 12'h333;
rom[82776] = 12'h333;
rom[82777] = 12'h333;
rom[82778] = 12'h333;
rom[82779] = 12'h333;
rom[82780] = 12'h222;
rom[82781] = 12'h222;
rom[82782] = 12'h222;
rom[82783] = 12'h222;
rom[82784] = 12'h222;
rom[82785] = 12'h222;
rom[82786] = 12'h222;
rom[82787] = 12'h222;
rom[82788] = 12'h222;
rom[82789] = 12'h222;
rom[82790] = 12'h222;
rom[82791] = 12'h222;
rom[82792] = 12'h222;
rom[82793] = 12'h222;
rom[82794] = 12'h222;
rom[82795] = 12'h222;
rom[82796] = 12'h222;
rom[82797] = 12'h222;
rom[82798] = 12'h222;
rom[82799] = 12'h222;
rom[82800] = 12'hfff;
rom[82801] = 12'hfff;
rom[82802] = 12'hfff;
rom[82803] = 12'hfff;
rom[82804] = 12'hfff;
rom[82805] = 12'hfff;
rom[82806] = 12'hfff;
rom[82807] = 12'hfff;
rom[82808] = 12'hfff;
rom[82809] = 12'hfff;
rom[82810] = 12'hfff;
rom[82811] = 12'hfff;
rom[82812] = 12'hfff;
rom[82813] = 12'hfff;
rom[82814] = 12'hfff;
rom[82815] = 12'hfff;
rom[82816] = 12'hfff;
rom[82817] = 12'hfff;
rom[82818] = 12'hfff;
rom[82819] = 12'hfff;
rom[82820] = 12'hfff;
rom[82821] = 12'hfff;
rom[82822] = 12'hfff;
rom[82823] = 12'hfff;
rom[82824] = 12'hfff;
rom[82825] = 12'hfff;
rom[82826] = 12'hfff;
rom[82827] = 12'hfff;
rom[82828] = 12'hfff;
rom[82829] = 12'hfff;
rom[82830] = 12'hfff;
rom[82831] = 12'hfff;
rom[82832] = 12'hfff;
rom[82833] = 12'hfff;
rom[82834] = 12'hfff;
rom[82835] = 12'hfff;
rom[82836] = 12'hfff;
rom[82837] = 12'hfff;
rom[82838] = 12'hfff;
rom[82839] = 12'hfff;
rom[82840] = 12'hfff;
rom[82841] = 12'hfff;
rom[82842] = 12'hfff;
rom[82843] = 12'hfff;
rom[82844] = 12'hfff;
rom[82845] = 12'hfff;
rom[82846] = 12'hfff;
rom[82847] = 12'hfff;
rom[82848] = 12'hfff;
rom[82849] = 12'hfff;
rom[82850] = 12'hfff;
rom[82851] = 12'hfff;
rom[82852] = 12'hfff;
rom[82853] = 12'hfff;
rom[82854] = 12'hfff;
rom[82855] = 12'hfff;
rom[82856] = 12'hfff;
rom[82857] = 12'hfff;
rom[82858] = 12'hfff;
rom[82859] = 12'hfff;
rom[82860] = 12'hfff;
rom[82861] = 12'hfff;
rom[82862] = 12'hfff;
rom[82863] = 12'hfff;
rom[82864] = 12'hfff;
rom[82865] = 12'hfff;
rom[82866] = 12'hfff;
rom[82867] = 12'hfff;
rom[82868] = 12'hfff;
rom[82869] = 12'hfff;
rom[82870] = 12'hfff;
rom[82871] = 12'hfff;
rom[82872] = 12'hfff;
rom[82873] = 12'hfff;
rom[82874] = 12'hfff;
rom[82875] = 12'hfff;
rom[82876] = 12'hfff;
rom[82877] = 12'hfff;
rom[82878] = 12'hfff;
rom[82879] = 12'hfff;
rom[82880] = 12'hfff;
rom[82881] = 12'hfff;
rom[82882] = 12'hfff;
rom[82883] = 12'hfff;
rom[82884] = 12'hfff;
rom[82885] = 12'hfff;
rom[82886] = 12'hfff;
rom[82887] = 12'hfff;
rom[82888] = 12'hfff;
rom[82889] = 12'hfff;
rom[82890] = 12'hfff;
rom[82891] = 12'hfff;
rom[82892] = 12'hfff;
rom[82893] = 12'hfff;
rom[82894] = 12'hfff;
rom[82895] = 12'hfff;
rom[82896] = 12'hfff;
rom[82897] = 12'hfff;
rom[82898] = 12'hfff;
rom[82899] = 12'hfff;
rom[82900] = 12'hfff;
rom[82901] = 12'hfff;
rom[82902] = 12'hfff;
rom[82903] = 12'hfff;
rom[82904] = 12'hfff;
rom[82905] = 12'hfff;
rom[82906] = 12'hfff;
rom[82907] = 12'hfff;
rom[82908] = 12'hfff;
rom[82909] = 12'hfff;
rom[82910] = 12'hfff;
rom[82911] = 12'hfff;
rom[82912] = 12'hfff;
rom[82913] = 12'hfff;
rom[82914] = 12'hfff;
rom[82915] = 12'hfff;
rom[82916] = 12'hfff;
rom[82917] = 12'hfff;
rom[82918] = 12'hfff;
rom[82919] = 12'hfff;
rom[82920] = 12'hfff;
rom[82921] = 12'hfff;
rom[82922] = 12'hfff;
rom[82923] = 12'hfff;
rom[82924] = 12'hfff;
rom[82925] = 12'hfff;
rom[82926] = 12'hfff;
rom[82927] = 12'hfff;
rom[82928] = 12'hfff;
rom[82929] = 12'hfff;
rom[82930] = 12'hfff;
rom[82931] = 12'hfff;
rom[82932] = 12'hfff;
rom[82933] = 12'heee;
rom[82934] = 12'heee;
rom[82935] = 12'heee;
rom[82936] = 12'heee;
rom[82937] = 12'hddd;
rom[82938] = 12'hddd;
rom[82939] = 12'hccc;
rom[82940] = 12'hccc;
rom[82941] = 12'hbbb;
rom[82942] = 12'hbbb;
rom[82943] = 12'hbbb;
rom[82944] = 12'haaa;
rom[82945] = 12'h999;
rom[82946] = 12'h999;
rom[82947] = 12'h888;
rom[82948] = 12'h888;
rom[82949] = 12'h777;
rom[82950] = 12'h777;
rom[82951] = 12'h777;
rom[82952] = 12'h666;
rom[82953] = 12'h666;
rom[82954] = 12'h666;
rom[82955] = 12'h555;
rom[82956] = 12'h555;
rom[82957] = 12'h555;
rom[82958] = 12'h555;
rom[82959] = 12'h555;
rom[82960] = 12'h555;
rom[82961] = 12'h555;
rom[82962] = 12'h444;
rom[82963] = 12'h444;
rom[82964] = 12'h444;
rom[82965] = 12'h444;
rom[82966] = 12'h444;
rom[82967] = 12'h444;
rom[82968] = 12'h333;
rom[82969] = 12'h333;
rom[82970] = 12'h333;
rom[82971] = 12'h333;
rom[82972] = 12'h333;
rom[82973] = 12'h333;
rom[82974] = 12'h333;
rom[82975] = 12'h444;
rom[82976] = 12'h444;
rom[82977] = 12'h444;
rom[82978] = 12'h444;
rom[82979] = 12'h444;
rom[82980] = 12'h444;
rom[82981] = 12'h444;
rom[82982] = 12'h444;
rom[82983] = 12'h444;
rom[82984] = 12'h444;
rom[82985] = 12'h444;
rom[82986] = 12'h444;
rom[82987] = 12'h444;
rom[82988] = 12'h444;
rom[82989] = 12'h555;
rom[82990] = 12'h555;
rom[82991] = 12'h555;
rom[82992] = 12'h444;
rom[82993] = 12'h444;
rom[82994] = 12'h444;
rom[82995] = 12'h444;
rom[82996] = 12'h333;
rom[82997] = 12'h333;
rom[82998] = 12'h333;
rom[82999] = 12'h333;
rom[83000] = 12'h333;
rom[83001] = 12'h333;
rom[83002] = 12'h333;
rom[83003] = 12'h444;
rom[83004] = 12'h444;
rom[83005] = 12'h555;
rom[83006] = 12'h777;
rom[83007] = 12'h888;
rom[83008] = 12'haaa;
rom[83009] = 12'haaa;
rom[83010] = 12'h999;
rom[83011] = 12'h999;
rom[83012] = 12'h777;
rom[83013] = 12'h666;
rom[83014] = 12'h555;
rom[83015] = 12'h444;
rom[83016] = 12'h444;
rom[83017] = 12'h444;
rom[83018] = 12'h444;
rom[83019] = 12'h444;
rom[83020] = 12'h333;
rom[83021] = 12'h333;
rom[83022] = 12'h333;
rom[83023] = 12'h333;
rom[83024] = 12'h222;
rom[83025] = 12'h222;
rom[83026] = 12'h222;
rom[83027] = 12'h222;
rom[83028] = 12'h222;
rom[83029] = 12'h222;
rom[83030] = 12'h111;
rom[83031] = 12'h111;
rom[83032] = 12'h111;
rom[83033] = 12'h111;
rom[83034] = 12'h111;
rom[83035] = 12'h111;
rom[83036] = 12'h111;
rom[83037] = 12'h111;
rom[83038] = 12'h111;
rom[83039] = 12'h111;
rom[83040] = 12'h111;
rom[83041] = 12'h111;
rom[83042] = 12'h111;
rom[83043] = 12'h  0;
rom[83044] = 12'h  0;
rom[83045] = 12'h  0;
rom[83046] = 12'h  0;
rom[83047] = 12'h  0;
rom[83048] = 12'h  0;
rom[83049] = 12'h  0;
rom[83050] = 12'h  0;
rom[83051] = 12'h  0;
rom[83052] = 12'h  0;
rom[83053] = 12'h  0;
rom[83054] = 12'h  0;
rom[83055] = 12'h  0;
rom[83056] = 12'h  0;
rom[83057] = 12'h  0;
rom[83058] = 12'h  0;
rom[83059] = 12'h  0;
rom[83060] = 12'h  0;
rom[83061] = 12'h  0;
rom[83062] = 12'h  0;
rom[83063] = 12'h  0;
rom[83064] = 12'h  0;
rom[83065] = 12'h  0;
rom[83066] = 12'h111;
rom[83067] = 12'h111;
rom[83068] = 12'h111;
rom[83069] = 12'h111;
rom[83070] = 12'h111;
rom[83071] = 12'h111;
rom[83072] = 12'h222;
rom[83073] = 12'h222;
rom[83074] = 12'h222;
rom[83075] = 12'h333;
rom[83076] = 12'h333;
rom[83077] = 12'h333;
rom[83078] = 12'h444;
rom[83079] = 12'h555;
rom[83080] = 12'h888;
rom[83081] = 12'haaa;
rom[83082] = 12'h999;
rom[83083] = 12'h777;
rom[83084] = 12'h666;
rom[83085] = 12'h666;
rom[83086] = 12'h666;
rom[83087] = 12'h555;
rom[83088] = 12'h555;
rom[83089] = 12'h555;
rom[83090] = 12'h555;
rom[83091] = 12'h555;
rom[83092] = 12'h555;
rom[83093] = 12'h555;
rom[83094] = 12'h555;
rom[83095] = 12'h555;
rom[83096] = 12'h666;
rom[83097] = 12'h666;
rom[83098] = 12'h666;
rom[83099] = 12'h666;
rom[83100] = 12'h666;
rom[83101] = 12'h666;
rom[83102] = 12'h777;
rom[83103] = 12'h888;
rom[83104] = 12'h888;
rom[83105] = 12'h999;
rom[83106] = 12'h999;
rom[83107] = 12'haaa;
rom[83108] = 12'hbbb;
rom[83109] = 12'hccc;
rom[83110] = 12'hccc;
rom[83111] = 12'hbbb;
rom[83112] = 12'haaa;
rom[83113] = 12'h999;
rom[83114] = 12'h888;
rom[83115] = 12'h888;
rom[83116] = 12'h888;
rom[83117] = 12'h777;
rom[83118] = 12'h777;
rom[83119] = 12'h777;
rom[83120] = 12'h888;
rom[83121] = 12'h888;
rom[83122] = 12'h888;
rom[83123] = 12'h888;
rom[83124] = 12'h888;
rom[83125] = 12'h888;
rom[83126] = 12'h888;
rom[83127] = 12'h777;
rom[83128] = 12'h777;
rom[83129] = 12'h777;
rom[83130] = 12'h666;
rom[83131] = 12'h666;
rom[83132] = 12'h666;
rom[83133] = 12'h666;
rom[83134] = 12'h666;
rom[83135] = 12'h555;
rom[83136] = 12'h666;
rom[83137] = 12'h555;
rom[83138] = 12'h555;
rom[83139] = 12'h444;
rom[83140] = 12'h444;
rom[83141] = 12'h444;
rom[83142] = 12'h444;
rom[83143] = 12'h333;
rom[83144] = 12'h333;
rom[83145] = 12'h333;
rom[83146] = 12'h333;
rom[83147] = 12'h333;
rom[83148] = 12'h333;
rom[83149] = 12'h333;
rom[83150] = 12'h333;
rom[83151] = 12'h333;
rom[83152] = 12'h333;
rom[83153] = 12'h333;
rom[83154] = 12'h333;
rom[83155] = 12'h333;
rom[83156] = 12'h444;
rom[83157] = 12'h444;
rom[83158] = 12'h444;
rom[83159] = 12'h444;
rom[83160] = 12'h444;
rom[83161] = 12'h333;
rom[83162] = 12'h333;
rom[83163] = 12'h333;
rom[83164] = 12'h333;
rom[83165] = 12'h444;
rom[83166] = 12'h444;
rom[83167] = 12'h333;
rom[83168] = 12'h333;
rom[83169] = 12'h333;
rom[83170] = 12'h333;
rom[83171] = 12'h333;
rom[83172] = 12'h333;
rom[83173] = 12'h333;
rom[83174] = 12'h333;
rom[83175] = 12'h333;
rom[83176] = 12'h333;
rom[83177] = 12'h333;
rom[83178] = 12'h333;
rom[83179] = 12'h333;
rom[83180] = 12'h222;
rom[83181] = 12'h222;
rom[83182] = 12'h222;
rom[83183] = 12'h222;
rom[83184] = 12'h222;
rom[83185] = 12'h222;
rom[83186] = 12'h222;
rom[83187] = 12'h222;
rom[83188] = 12'h222;
rom[83189] = 12'h222;
rom[83190] = 12'h222;
rom[83191] = 12'h222;
rom[83192] = 12'h222;
rom[83193] = 12'h222;
rom[83194] = 12'h222;
rom[83195] = 12'h222;
rom[83196] = 12'h222;
rom[83197] = 12'h222;
rom[83198] = 12'h222;
rom[83199] = 12'h222;
rom[83200] = 12'hfff;
rom[83201] = 12'hfff;
rom[83202] = 12'hfff;
rom[83203] = 12'hfff;
rom[83204] = 12'hfff;
rom[83205] = 12'hfff;
rom[83206] = 12'hfff;
rom[83207] = 12'hfff;
rom[83208] = 12'hfff;
rom[83209] = 12'hfff;
rom[83210] = 12'hfff;
rom[83211] = 12'hfff;
rom[83212] = 12'hfff;
rom[83213] = 12'hfff;
rom[83214] = 12'hfff;
rom[83215] = 12'hfff;
rom[83216] = 12'hfff;
rom[83217] = 12'hfff;
rom[83218] = 12'hfff;
rom[83219] = 12'hfff;
rom[83220] = 12'hfff;
rom[83221] = 12'hfff;
rom[83222] = 12'hfff;
rom[83223] = 12'hfff;
rom[83224] = 12'hfff;
rom[83225] = 12'hfff;
rom[83226] = 12'hfff;
rom[83227] = 12'hfff;
rom[83228] = 12'hfff;
rom[83229] = 12'hfff;
rom[83230] = 12'hfff;
rom[83231] = 12'hfff;
rom[83232] = 12'hfff;
rom[83233] = 12'hfff;
rom[83234] = 12'hfff;
rom[83235] = 12'hfff;
rom[83236] = 12'hfff;
rom[83237] = 12'hfff;
rom[83238] = 12'hfff;
rom[83239] = 12'hfff;
rom[83240] = 12'hfff;
rom[83241] = 12'hfff;
rom[83242] = 12'hfff;
rom[83243] = 12'hfff;
rom[83244] = 12'hfff;
rom[83245] = 12'hfff;
rom[83246] = 12'hfff;
rom[83247] = 12'hfff;
rom[83248] = 12'hfff;
rom[83249] = 12'hfff;
rom[83250] = 12'hfff;
rom[83251] = 12'hfff;
rom[83252] = 12'hfff;
rom[83253] = 12'hfff;
rom[83254] = 12'hfff;
rom[83255] = 12'hfff;
rom[83256] = 12'hfff;
rom[83257] = 12'hfff;
rom[83258] = 12'hfff;
rom[83259] = 12'hfff;
rom[83260] = 12'hfff;
rom[83261] = 12'hfff;
rom[83262] = 12'hfff;
rom[83263] = 12'hfff;
rom[83264] = 12'hfff;
rom[83265] = 12'hfff;
rom[83266] = 12'hfff;
rom[83267] = 12'hfff;
rom[83268] = 12'hfff;
rom[83269] = 12'hfff;
rom[83270] = 12'hfff;
rom[83271] = 12'hfff;
rom[83272] = 12'hfff;
rom[83273] = 12'hfff;
rom[83274] = 12'hfff;
rom[83275] = 12'hfff;
rom[83276] = 12'hfff;
rom[83277] = 12'hfff;
rom[83278] = 12'hfff;
rom[83279] = 12'hfff;
rom[83280] = 12'hfff;
rom[83281] = 12'hfff;
rom[83282] = 12'hfff;
rom[83283] = 12'hfff;
rom[83284] = 12'hfff;
rom[83285] = 12'hfff;
rom[83286] = 12'hfff;
rom[83287] = 12'hfff;
rom[83288] = 12'hfff;
rom[83289] = 12'hfff;
rom[83290] = 12'hfff;
rom[83291] = 12'hfff;
rom[83292] = 12'hfff;
rom[83293] = 12'hfff;
rom[83294] = 12'hfff;
rom[83295] = 12'hfff;
rom[83296] = 12'hfff;
rom[83297] = 12'hfff;
rom[83298] = 12'hfff;
rom[83299] = 12'hfff;
rom[83300] = 12'hfff;
rom[83301] = 12'hfff;
rom[83302] = 12'hfff;
rom[83303] = 12'hfff;
rom[83304] = 12'hfff;
rom[83305] = 12'hfff;
rom[83306] = 12'hfff;
rom[83307] = 12'hfff;
rom[83308] = 12'hfff;
rom[83309] = 12'hfff;
rom[83310] = 12'hfff;
rom[83311] = 12'hfff;
rom[83312] = 12'hfff;
rom[83313] = 12'hfff;
rom[83314] = 12'hfff;
rom[83315] = 12'hfff;
rom[83316] = 12'hfff;
rom[83317] = 12'hfff;
rom[83318] = 12'hfff;
rom[83319] = 12'hfff;
rom[83320] = 12'hfff;
rom[83321] = 12'hfff;
rom[83322] = 12'heee;
rom[83323] = 12'heee;
rom[83324] = 12'heee;
rom[83325] = 12'heee;
rom[83326] = 12'heee;
rom[83327] = 12'heee;
rom[83328] = 12'heee;
rom[83329] = 12'heee;
rom[83330] = 12'heee;
rom[83331] = 12'heee;
rom[83332] = 12'heee;
rom[83333] = 12'heee;
rom[83334] = 12'heee;
rom[83335] = 12'heee;
rom[83336] = 12'heee;
rom[83337] = 12'heee;
rom[83338] = 12'heee;
rom[83339] = 12'hddd;
rom[83340] = 12'hddd;
rom[83341] = 12'hccc;
rom[83342] = 12'hccc;
rom[83343] = 12'hbbb;
rom[83344] = 12'hbbb;
rom[83345] = 12'hbbb;
rom[83346] = 12'haaa;
rom[83347] = 12'h999;
rom[83348] = 12'h999;
rom[83349] = 12'h888;
rom[83350] = 12'h888;
rom[83351] = 12'h777;
rom[83352] = 12'h777;
rom[83353] = 12'h666;
rom[83354] = 12'h666;
rom[83355] = 12'h555;
rom[83356] = 12'h555;
rom[83357] = 12'h555;
rom[83358] = 12'h555;
rom[83359] = 12'h555;
rom[83360] = 12'h555;
rom[83361] = 12'h444;
rom[83362] = 12'h444;
rom[83363] = 12'h444;
rom[83364] = 12'h444;
rom[83365] = 12'h444;
rom[83366] = 12'h444;
rom[83367] = 12'h444;
rom[83368] = 12'h333;
rom[83369] = 12'h333;
rom[83370] = 12'h333;
rom[83371] = 12'h333;
rom[83372] = 12'h333;
rom[83373] = 12'h444;
rom[83374] = 12'h444;
rom[83375] = 12'h444;
rom[83376] = 12'h444;
rom[83377] = 12'h444;
rom[83378] = 12'h444;
rom[83379] = 12'h444;
rom[83380] = 12'h444;
rom[83381] = 12'h444;
rom[83382] = 12'h444;
rom[83383] = 12'h444;
rom[83384] = 12'h444;
rom[83385] = 12'h444;
rom[83386] = 12'h444;
rom[83387] = 12'h555;
rom[83388] = 12'h555;
rom[83389] = 12'h555;
rom[83390] = 12'h555;
rom[83391] = 12'h444;
rom[83392] = 12'h444;
rom[83393] = 12'h444;
rom[83394] = 12'h444;
rom[83395] = 12'h444;
rom[83396] = 12'h333;
rom[83397] = 12'h333;
rom[83398] = 12'h333;
rom[83399] = 12'h333;
rom[83400] = 12'h333;
rom[83401] = 12'h333;
rom[83402] = 12'h333;
rom[83403] = 12'h444;
rom[83404] = 12'h444;
rom[83405] = 12'h555;
rom[83406] = 12'h666;
rom[83407] = 12'h777;
rom[83408] = 12'h888;
rom[83409] = 12'haaa;
rom[83410] = 12'haaa;
rom[83411] = 12'h999;
rom[83412] = 12'h888;
rom[83413] = 12'h777;
rom[83414] = 12'h666;
rom[83415] = 12'h444;
rom[83416] = 12'h444;
rom[83417] = 12'h444;
rom[83418] = 12'h444;
rom[83419] = 12'h333;
rom[83420] = 12'h333;
rom[83421] = 12'h333;
rom[83422] = 12'h333;
rom[83423] = 12'h222;
rom[83424] = 12'h222;
rom[83425] = 12'h222;
rom[83426] = 12'h222;
rom[83427] = 12'h222;
rom[83428] = 12'h111;
rom[83429] = 12'h111;
rom[83430] = 12'h111;
rom[83431] = 12'h111;
rom[83432] = 12'h111;
rom[83433] = 12'h111;
rom[83434] = 12'h111;
rom[83435] = 12'h  0;
rom[83436] = 12'h  0;
rom[83437] = 12'h111;
rom[83438] = 12'h111;
rom[83439] = 12'h111;
rom[83440] = 12'h111;
rom[83441] = 12'h111;
rom[83442] = 12'h111;
rom[83443] = 12'h  0;
rom[83444] = 12'h  0;
rom[83445] = 12'h  0;
rom[83446] = 12'h  0;
rom[83447] = 12'h  0;
rom[83448] = 12'h  0;
rom[83449] = 12'h  0;
rom[83450] = 12'h  0;
rom[83451] = 12'h  0;
rom[83452] = 12'h  0;
rom[83453] = 12'h  0;
rom[83454] = 12'h  0;
rom[83455] = 12'h  0;
rom[83456] = 12'h  0;
rom[83457] = 12'h  0;
rom[83458] = 12'h  0;
rom[83459] = 12'h  0;
rom[83460] = 12'h  0;
rom[83461] = 12'h  0;
rom[83462] = 12'h  0;
rom[83463] = 12'h111;
rom[83464] = 12'h111;
rom[83465] = 12'h111;
rom[83466] = 12'h111;
rom[83467] = 12'h111;
rom[83468] = 12'h111;
rom[83469] = 12'h111;
rom[83470] = 12'h111;
rom[83471] = 12'h111;
rom[83472] = 12'h222;
rom[83473] = 12'h222;
rom[83474] = 12'h222;
rom[83475] = 12'h222;
rom[83476] = 12'h333;
rom[83477] = 12'h333;
rom[83478] = 12'h444;
rom[83479] = 12'h555;
rom[83480] = 12'h777;
rom[83481] = 12'h999;
rom[83482] = 12'haaa;
rom[83483] = 12'h888;
rom[83484] = 12'h666;
rom[83485] = 12'h666;
rom[83486] = 12'h666;
rom[83487] = 12'h666;
rom[83488] = 12'h555;
rom[83489] = 12'h555;
rom[83490] = 12'h555;
rom[83491] = 12'h555;
rom[83492] = 12'h555;
rom[83493] = 12'h555;
rom[83494] = 12'h555;
rom[83495] = 12'h555;
rom[83496] = 12'h666;
rom[83497] = 12'h666;
rom[83498] = 12'h666;
rom[83499] = 12'h666;
rom[83500] = 12'h666;
rom[83501] = 12'h777;
rom[83502] = 12'h777;
rom[83503] = 12'h888;
rom[83504] = 12'h888;
rom[83505] = 12'h888;
rom[83506] = 12'h999;
rom[83507] = 12'haaa;
rom[83508] = 12'hbbb;
rom[83509] = 12'hccc;
rom[83510] = 12'hbbb;
rom[83511] = 12'haaa;
rom[83512] = 12'h999;
rom[83513] = 12'h888;
rom[83514] = 12'h888;
rom[83515] = 12'h777;
rom[83516] = 12'h888;
rom[83517] = 12'h888;
rom[83518] = 12'h777;
rom[83519] = 12'h777;
rom[83520] = 12'h777;
rom[83521] = 12'h777;
rom[83522] = 12'h888;
rom[83523] = 12'h888;
rom[83524] = 12'h888;
rom[83525] = 12'h888;
rom[83526] = 12'h888;
rom[83527] = 12'h777;
rom[83528] = 12'h777;
rom[83529] = 12'h777;
rom[83530] = 12'h777;
rom[83531] = 12'h666;
rom[83532] = 12'h666;
rom[83533] = 12'h666;
rom[83534] = 12'h666;
rom[83535] = 12'h666;
rom[83536] = 12'h555;
rom[83537] = 12'h555;
rom[83538] = 12'h555;
rom[83539] = 12'h555;
rom[83540] = 12'h444;
rom[83541] = 12'h444;
rom[83542] = 12'h444;
rom[83543] = 12'h444;
rom[83544] = 12'h333;
rom[83545] = 12'h333;
rom[83546] = 12'h333;
rom[83547] = 12'h333;
rom[83548] = 12'h333;
rom[83549] = 12'h333;
rom[83550] = 12'h333;
rom[83551] = 12'h333;
rom[83552] = 12'h333;
rom[83553] = 12'h333;
rom[83554] = 12'h333;
rom[83555] = 12'h444;
rom[83556] = 12'h444;
rom[83557] = 12'h444;
rom[83558] = 12'h444;
rom[83559] = 12'h444;
rom[83560] = 12'h444;
rom[83561] = 12'h444;
rom[83562] = 12'h444;
rom[83563] = 12'h333;
rom[83564] = 12'h333;
rom[83565] = 12'h333;
rom[83566] = 12'h333;
rom[83567] = 12'h333;
rom[83568] = 12'h333;
rom[83569] = 12'h333;
rom[83570] = 12'h333;
rom[83571] = 12'h333;
rom[83572] = 12'h333;
rom[83573] = 12'h333;
rom[83574] = 12'h333;
rom[83575] = 12'h333;
rom[83576] = 12'h333;
rom[83577] = 12'h333;
rom[83578] = 12'h333;
rom[83579] = 12'h333;
rom[83580] = 12'h222;
rom[83581] = 12'h222;
rom[83582] = 12'h222;
rom[83583] = 12'h222;
rom[83584] = 12'h222;
rom[83585] = 12'h222;
rom[83586] = 12'h222;
rom[83587] = 12'h222;
rom[83588] = 12'h222;
rom[83589] = 12'h222;
rom[83590] = 12'h222;
rom[83591] = 12'h222;
rom[83592] = 12'h222;
rom[83593] = 12'h222;
rom[83594] = 12'h222;
rom[83595] = 12'h222;
rom[83596] = 12'h222;
rom[83597] = 12'h222;
rom[83598] = 12'h222;
rom[83599] = 12'h222;
rom[83600] = 12'hfff;
rom[83601] = 12'hfff;
rom[83602] = 12'hfff;
rom[83603] = 12'hfff;
rom[83604] = 12'hfff;
rom[83605] = 12'hfff;
rom[83606] = 12'hfff;
rom[83607] = 12'hfff;
rom[83608] = 12'hfff;
rom[83609] = 12'hfff;
rom[83610] = 12'hfff;
rom[83611] = 12'hfff;
rom[83612] = 12'hfff;
rom[83613] = 12'hfff;
rom[83614] = 12'hfff;
rom[83615] = 12'hfff;
rom[83616] = 12'hfff;
rom[83617] = 12'hfff;
rom[83618] = 12'hfff;
rom[83619] = 12'hfff;
rom[83620] = 12'hfff;
rom[83621] = 12'hfff;
rom[83622] = 12'hfff;
rom[83623] = 12'hfff;
rom[83624] = 12'hfff;
rom[83625] = 12'hfff;
rom[83626] = 12'hfff;
rom[83627] = 12'hfff;
rom[83628] = 12'hfff;
rom[83629] = 12'hfff;
rom[83630] = 12'hfff;
rom[83631] = 12'hfff;
rom[83632] = 12'hfff;
rom[83633] = 12'hfff;
rom[83634] = 12'hfff;
rom[83635] = 12'hfff;
rom[83636] = 12'hfff;
rom[83637] = 12'hfff;
rom[83638] = 12'hfff;
rom[83639] = 12'hfff;
rom[83640] = 12'hfff;
rom[83641] = 12'hfff;
rom[83642] = 12'hfff;
rom[83643] = 12'hfff;
rom[83644] = 12'hfff;
rom[83645] = 12'hfff;
rom[83646] = 12'hfff;
rom[83647] = 12'hfff;
rom[83648] = 12'hfff;
rom[83649] = 12'hfff;
rom[83650] = 12'hfff;
rom[83651] = 12'hfff;
rom[83652] = 12'hfff;
rom[83653] = 12'hfff;
rom[83654] = 12'hfff;
rom[83655] = 12'hfff;
rom[83656] = 12'hfff;
rom[83657] = 12'hfff;
rom[83658] = 12'hfff;
rom[83659] = 12'hfff;
rom[83660] = 12'hfff;
rom[83661] = 12'hfff;
rom[83662] = 12'hfff;
rom[83663] = 12'hfff;
rom[83664] = 12'hfff;
rom[83665] = 12'hfff;
rom[83666] = 12'hfff;
rom[83667] = 12'hfff;
rom[83668] = 12'hfff;
rom[83669] = 12'hfff;
rom[83670] = 12'hfff;
rom[83671] = 12'hfff;
rom[83672] = 12'hfff;
rom[83673] = 12'hfff;
rom[83674] = 12'hfff;
rom[83675] = 12'hfff;
rom[83676] = 12'hfff;
rom[83677] = 12'hfff;
rom[83678] = 12'hfff;
rom[83679] = 12'hfff;
rom[83680] = 12'hfff;
rom[83681] = 12'hfff;
rom[83682] = 12'hfff;
rom[83683] = 12'hfff;
rom[83684] = 12'hfff;
rom[83685] = 12'hfff;
rom[83686] = 12'hfff;
rom[83687] = 12'hfff;
rom[83688] = 12'hfff;
rom[83689] = 12'hfff;
rom[83690] = 12'hfff;
rom[83691] = 12'hfff;
rom[83692] = 12'hfff;
rom[83693] = 12'hfff;
rom[83694] = 12'hfff;
rom[83695] = 12'hfff;
rom[83696] = 12'hfff;
rom[83697] = 12'hfff;
rom[83698] = 12'hfff;
rom[83699] = 12'hfff;
rom[83700] = 12'hfff;
rom[83701] = 12'hfff;
rom[83702] = 12'hfff;
rom[83703] = 12'hfff;
rom[83704] = 12'hfff;
rom[83705] = 12'hfff;
rom[83706] = 12'hfff;
rom[83707] = 12'hfff;
rom[83708] = 12'hfff;
rom[83709] = 12'hfff;
rom[83710] = 12'hfff;
rom[83711] = 12'hfff;
rom[83712] = 12'hfff;
rom[83713] = 12'hfff;
rom[83714] = 12'hfff;
rom[83715] = 12'hfff;
rom[83716] = 12'hfff;
rom[83717] = 12'hfff;
rom[83718] = 12'hfff;
rom[83719] = 12'hfff;
rom[83720] = 12'hfff;
rom[83721] = 12'hfff;
rom[83722] = 12'heee;
rom[83723] = 12'heee;
rom[83724] = 12'heee;
rom[83725] = 12'heee;
rom[83726] = 12'heee;
rom[83727] = 12'heee;
rom[83728] = 12'heee;
rom[83729] = 12'heee;
rom[83730] = 12'heee;
rom[83731] = 12'heee;
rom[83732] = 12'heee;
rom[83733] = 12'heee;
rom[83734] = 12'heee;
rom[83735] = 12'heee;
rom[83736] = 12'heee;
rom[83737] = 12'heee;
rom[83738] = 12'heee;
rom[83739] = 12'heee;
rom[83740] = 12'hddd;
rom[83741] = 12'hddd;
rom[83742] = 12'hddd;
rom[83743] = 12'hccc;
rom[83744] = 12'hccc;
rom[83745] = 12'hbbb;
rom[83746] = 12'hbbb;
rom[83747] = 12'haaa;
rom[83748] = 12'haaa;
rom[83749] = 12'h999;
rom[83750] = 12'h888;
rom[83751] = 12'h888;
rom[83752] = 12'h777;
rom[83753] = 12'h777;
rom[83754] = 12'h666;
rom[83755] = 12'h666;
rom[83756] = 12'h555;
rom[83757] = 12'h555;
rom[83758] = 12'h555;
rom[83759] = 12'h555;
rom[83760] = 12'h555;
rom[83761] = 12'h444;
rom[83762] = 12'h444;
rom[83763] = 12'h444;
rom[83764] = 12'h444;
rom[83765] = 12'h444;
rom[83766] = 12'h444;
rom[83767] = 12'h333;
rom[83768] = 12'h333;
rom[83769] = 12'h333;
rom[83770] = 12'h333;
rom[83771] = 12'h333;
rom[83772] = 12'h333;
rom[83773] = 12'h333;
rom[83774] = 12'h444;
rom[83775] = 12'h444;
rom[83776] = 12'h444;
rom[83777] = 12'h444;
rom[83778] = 12'h444;
rom[83779] = 12'h444;
rom[83780] = 12'h444;
rom[83781] = 12'h444;
rom[83782] = 12'h555;
rom[83783] = 12'h555;
rom[83784] = 12'h444;
rom[83785] = 12'h444;
rom[83786] = 12'h444;
rom[83787] = 12'h555;
rom[83788] = 12'h555;
rom[83789] = 12'h555;
rom[83790] = 12'h555;
rom[83791] = 12'h555;
rom[83792] = 12'h444;
rom[83793] = 12'h444;
rom[83794] = 12'h444;
rom[83795] = 12'h333;
rom[83796] = 12'h333;
rom[83797] = 12'h333;
rom[83798] = 12'h333;
rom[83799] = 12'h333;
rom[83800] = 12'h333;
rom[83801] = 12'h333;
rom[83802] = 12'h333;
rom[83803] = 12'h444;
rom[83804] = 12'h444;
rom[83805] = 12'h555;
rom[83806] = 12'h666;
rom[83807] = 12'h666;
rom[83808] = 12'h777;
rom[83809] = 12'h888;
rom[83810] = 12'h999;
rom[83811] = 12'h999;
rom[83812] = 12'h999;
rom[83813] = 12'h888;
rom[83814] = 12'h666;
rom[83815] = 12'h555;
rom[83816] = 12'h444;
rom[83817] = 12'h444;
rom[83818] = 12'h333;
rom[83819] = 12'h333;
rom[83820] = 12'h333;
rom[83821] = 12'h333;
rom[83822] = 12'h222;
rom[83823] = 12'h222;
rom[83824] = 12'h222;
rom[83825] = 12'h222;
rom[83826] = 12'h222;
rom[83827] = 12'h222;
rom[83828] = 12'h111;
rom[83829] = 12'h111;
rom[83830] = 12'h111;
rom[83831] = 12'h111;
rom[83832] = 12'h111;
rom[83833] = 12'h  0;
rom[83834] = 12'h  0;
rom[83835] = 12'h  0;
rom[83836] = 12'h  0;
rom[83837] = 12'h  0;
rom[83838] = 12'h  0;
rom[83839] = 12'h  0;
rom[83840] = 12'h  0;
rom[83841] = 12'h  0;
rom[83842] = 12'h  0;
rom[83843] = 12'h  0;
rom[83844] = 12'h  0;
rom[83845] = 12'h  0;
rom[83846] = 12'h  0;
rom[83847] = 12'h  0;
rom[83848] = 12'h  0;
rom[83849] = 12'h  0;
rom[83850] = 12'h  0;
rom[83851] = 12'h  0;
rom[83852] = 12'h  0;
rom[83853] = 12'h  0;
rom[83854] = 12'h  0;
rom[83855] = 12'h  0;
rom[83856] = 12'h  0;
rom[83857] = 12'h  0;
rom[83858] = 12'h  0;
rom[83859] = 12'h  0;
rom[83860] = 12'h  0;
rom[83861] = 12'h111;
rom[83862] = 12'h111;
rom[83863] = 12'h111;
rom[83864] = 12'h111;
rom[83865] = 12'h111;
rom[83866] = 12'h111;
rom[83867] = 12'h111;
rom[83868] = 12'h111;
rom[83869] = 12'h111;
rom[83870] = 12'h222;
rom[83871] = 12'h222;
rom[83872] = 12'h222;
rom[83873] = 12'h222;
rom[83874] = 12'h222;
rom[83875] = 12'h222;
rom[83876] = 12'h333;
rom[83877] = 12'h333;
rom[83878] = 12'h444;
rom[83879] = 12'h555;
rom[83880] = 12'h777;
rom[83881] = 12'h999;
rom[83882] = 12'haaa;
rom[83883] = 12'h888;
rom[83884] = 12'h666;
rom[83885] = 12'h666;
rom[83886] = 12'h666;
rom[83887] = 12'h666;
rom[83888] = 12'h666;
rom[83889] = 12'h666;
rom[83890] = 12'h555;
rom[83891] = 12'h555;
rom[83892] = 12'h555;
rom[83893] = 12'h666;
rom[83894] = 12'h666;
rom[83895] = 12'h666;
rom[83896] = 12'h666;
rom[83897] = 12'h666;
rom[83898] = 12'h777;
rom[83899] = 12'h777;
rom[83900] = 12'h777;
rom[83901] = 12'h777;
rom[83902] = 12'h777;
rom[83903] = 12'h888;
rom[83904] = 12'h888;
rom[83905] = 12'h888;
rom[83906] = 12'h999;
rom[83907] = 12'hbbb;
rom[83908] = 12'hccc;
rom[83909] = 12'hccc;
rom[83910] = 12'hbbb;
rom[83911] = 12'haaa;
rom[83912] = 12'h999;
rom[83913] = 12'h888;
rom[83914] = 12'h888;
rom[83915] = 12'h777;
rom[83916] = 12'h777;
rom[83917] = 12'h777;
rom[83918] = 12'h777;
rom[83919] = 12'h777;
rom[83920] = 12'h777;
rom[83921] = 12'h777;
rom[83922] = 12'h777;
rom[83923] = 12'h777;
rom[83924] = 12'h888;
rom[83925] = 12'h888;
rom[83926] = 12'h888;
rom[83927] = 12'h888;
rom[83928] = 12'h777;
rom[83929] = 12'h777;
rom[83930] = 12'h777;
rom[83931] = 12'h777;
rom[83932] = 12'h666;
rom[83933] = 12'h666;
rom[83934] = 12'h666;
rom[83935] = 12'h666;
rom[83936] = 12'h555;
rom[83937] = 12'h555;
rom[83938] = 12'h555;
rom[83939] = 12'h555;
rom[83940] = 12'h444;
rom[83941] = 12'h444;
rom[83942] = 12'h444;
rom[83943] = 12'h444;
rom[83944] = 12'h444;
rom[83945] = 12'h444;
rom[83946] = 12'h333;
rom[83947] = 12'h333;
rom[83948] = 12'h333;
rom[83949] = 12'h333;
rom[83950] = 12'h333;
rom[83951] = 12'h333;
rom[83952] = 12'h333;
rom[83953] = 12'h333;
rom[83954] = 12'h333;
rom[83955] = 12'h444;
rom[83956] = 12'h444;
rom[83957] = 12'h444;
rom[83958] = 12'h444;
rom[83959] = 12'h444;
rom[83960] = 12'h444;
rom[83961] = 12'h444;
rom[83962] = 12'h444;
rom[83963] = 12'h333;
rom[83964] = 12'h333;
rom[83965] = 12'h333;
rom[83966] = 12'h333;
rom[83967] = 12'h333;
rom[83968] = 12'h333;
rom[83969] = 12'h333;
rom[83970] = 12'h333;
rom[83971] = 12'h333;
rom[83972] = 12'h333;
rom[83973] = 12'h333;
rom[83974] = 12'h333;
rom[83975] = 12'h333;
rom[83976] = 12'h333;
rom[83977] = 12'h333;
rom[83978] = 12'h333;
rom[83979] = 12'h333;
rom[83980] = 12'h222;
rom[83981] = 12'h222;
rom[83982] = 12'h222;
rom[83983] = 12'h222;
rom[83984] = 12'h222;
rom[83985] = 12'h222;
rom[83986] = 12'h222;
rom[83987] = 12'h222;
rom[83988] = 12'h222;
rom[83989] = 12'h222;
rom[83990] = 12'h222;
rom[83991] = 12'h222;
rom[83992] = 12'h222;
rom[83993] = 12'h222;
rom[83994] = 12'h222;
rom[83995] = 12'h222;
rom[83996] = 12'h111;
rom[83997] = 12'h222;
rom[83998] = 12'h222;
rom[83999] = 12'h222;
rom[84000] = 12'hfff;
rom[84001] = 12'hfff;
rom[84002] = 12'hfff;
rom[84003] = 12'hfff;
rom[84004] = 12'hfff;
rom[84005] = 12'hfff;
rom[84006] = 12'hfff;
rom[84007] = 12'hfff;
rom[84008] = 12'hfff;
rom[84009] = 12'hfff;
rom[84010] = 12'hfff;
rom[84011] = 12'hfff;
rom[84012] = 12'hfff;
rom[84013] = 12'hfff;
rom[84014] = 12'hfff;
rom[84015] = 12'hfff;
rom[84016] = 12'hfff;
rom[84017] = 12'hfff;
rom[84018] = 12'hfff;
rom[84019] = 12'hfff;
rom[84020] = 12'hfff;
rom[84021] = 12'hfff;
rom[84022] = 12'hfff;
rom[84023] = 12'hfff;
rom[84024] = 12'hfff;
rom[84025] = 12'hfff;
rom[84026] = 12'hfff;
rom[84027] = 12'hfff;
rom[84028] = 12'hfff;
rom[84029] = 12'hfff;
rom[84030] = 12'hfff;
rom[84031] = 12'hfff;
rom[84032] = 12'hfff;
rom[84033] = 12'hfff;
rom[84034] = 12'hfff;
rom[84035] = 12'hfff;
rom[84036] = 12'hfff;
rom[84037] = 12'hfff;
rom[84038] = 12'hfff;
rom[84039] = 12'hfff;
rom[84040] = 12'hfff;
rom[84041] = 12'hfff;
rom[84042] = 12'hfff;
rom[84043] = 12'hfff;
rom[84044] = 12'hfff;
rom[84045] = 12'hfff;
rom[84046] = 12'hfff;
rom[84047] = 12'hfff;
rom[84048] = 12'hfff;
rom[84049] = 12'hfff;
rom[84050] = 12'hfff;
rom[84051] = 12'hfff;
rom[84052] = 12'hfff;
rom[84053] = 12'hfff;
rom[84054] = 12'hfff;
rom[84055] = 12'hfff;
rom[84056] = 12'hfff;
rom[84057] = 12'hfff;
rom[84058] = 12'hfff;
rom[84059] = 12'hfff;
rom[84060] = 12'hfff;
rom[84061] = 12'hfff;
rom[84062] = 12'hfff;
rom[84063] = 12'hfff;
rom[84064] = 12'hfff;
rom[84065] = 12'hfff;
rom[84066] = 12'hfff;
rom[84067] = 12'hfff;
rom[84068] = 12'hfff;
rom[84069] = 12'hfff;
rom[84070] = 12'hfff;
rom[84071] = 12'hfff;
rom[84072] = 12'hfff;
rom[84073] = 12'hfff;
rom[84074] = 12'hfff;
rom[84075] = 12'hfff;
rom[84076] = 12'hfff;
rom[84077] = 12'hfff;
rom[84078] = 12'hfff;
rom[84079] = 12'hfff;
rom[84080] = 12'hfff;
rom[84081] = 12'hfff;
rom[84082] = 12'hfff;
rom[84083] = 12'hfff;
rom[84084] = 12'hfff;
rom[84085] = 12'hfff;
rom[84086] = 12'hfff;
rom[84087] = 12'hfff;
rom[84088] = 12'hfff;
rom[84089] = 12'hfff;
rom[84090] = 12'hfff;
rom[84091] = 12'hfff;
rom[84092] = 12'hfff;
rom[84093] = 12'hfff;
rom[84094] = 12'hfff;
rom[84095] = 12'hfff;
rom[84096] = 12'hfff;
rom[84097] = 12'hfff;
rom[84098] = 12'hfff;
rom[84099] = 12'hfff;
rom[84100] = 12'hfff;
rom[84101] = 12'hfff;
rom[84102] = 12'hfff;
rom[84103] = 12'hfff;
rom[84104] = 12'hfff;
rom[84105] = 12'hfff;
rom[84106] = 12'hfff;
rom[84107] = 12'hfff;
rom[84108] = 12'hfff;
rom[84109] = 12'hfff;
rom[84110] = 12'hfff;
rom[84111] = 12'hfff;
rom[84112] = 12'hfff;
rom[84113] = 12'hfff;
rom[84114] = 12'hfff;
rom[84115] = 12'hfff;
rom[84116] = 12'hfff;
rom[84117] = 12'hfff;
rom[84118] = 12'hfff;
rom[84119] = 12'hfff;
rom[84120] = 12'hfff;
rom[84121] = 12'hfff;
rom[84122] = 12'hfff;
rom[84123] = 12'heee;
rom[84124] = 12'heee;
rom[84125] = 12'heee;
rom[84126] = 12'heee;
rom[84127] = 12'heee;
rom[84128] = 12'heee;
rom[84129] = 12'heee;
rom[84130] = 12'heee;
rom[84131] = 12'heee;
rom[84132] = 12'heee;
rom[84133] = 12'heee;
rom[84134] = 12'heee;
rom[84135] = 12'heee;
rom[84136] = 12'heee;
rom[84137] = 12'heee;
rom[84138] = 12'heee;
rom[84139] = 12'hddd;
rom[84140] = 12'hddd;
rom[84141] = 12'hddd;
rom[84142] = 12'hddd;
rom[84143] = 12'hddd;
rom[84144] = 12'hddd;
rom[84145] = 12'hccc;
rom[84146] = 12'hccc;
rom[84147] = 12'hbbb;
rom[84148] = 12'hbbb;
rom[84149] = 12'haaa;
rom[84150] = 12'h999;
rom[84151] = 12'h999;
rom[84152] = 12'h888;
rom[84153] = 12'h777;
rom[84154] = 12'h777;
rom[84155] = 12'h666;
rom[84156] = 12'h666;
rom[84157] = 12'h666;
rom[84158] = 12'h555;
rom[84159] = 12'h555;
rom[84160] = 12'h555;
rom[84161] = 12'h555;
rom[84162] = 12'h444;
rom[84163] = 12'h444;
rom[84164] = 12'h444;
rom[84165] = 12'h444;
rom[84166] = 12'h444;
rom[84167] = 12'h333;
rom[84168] = 12'h333;
rom[84169] = 12'h333;
rom[84170] = 12'h333;
rom[84171] = 12'h333;
rom[84172] = 12'h444;
rom[84173] = 12'h444;
rom[84174] = 12'h444;
rom[84175] = 12'h444;
rom[84176] = 12'h444;
rom[84177] = 12'h444;
rom[84178] = 12'h444;
rom[84179] = 12'h444;
rom[84180] = 12'h444;
rom[84181] = 12'h555;
rom[84182] = 12'h555;
rom[84183] = 12'h555;
rom[84184] = 12'h555;
rom[84185] = 12'h444;
rom[84186] = 12'h555;
rom[84187] = 12'h555;
rom[84188] = 12'h555;
rom[84189] = 12'h555;
rom[84190] = 12'h555;
rom[84191] = 12'h555;
rom[84192] = 12'h444;
rom[84193] = 12'h444;
rom[84194] = 12'h444;
rom[84195] = 12'h333;
rom[84196] = 12'h333;
rom[84197] = 12'h333;
rom[84198] = 12'h333;
rom[84199] = 12'h444;
rom[84200] = 12'h444;
rom[84201] = 12'h444;
rom[84202] = 12'h444;
rom[84203] = 12'h444;
rom[84204] = 12'h555;
rom[84205] = 12'h555;
rom[84206] = 12'h555;
rom[84207] = 12'h555;
rom[84208] = 12'h666;
rom[84209] = 12'h777;
rom[84210] = 12'h888;
rom[84211] = 12'h999;
rom[84212] = 12'h999;
rom[84213] = 12'h888;
rom[84214] = 12'h777;
rom[84215] = 12'h666;
rom[84216] = 12'h555;
rom[84217] = 12'h444;
rom[84218] = 12'h333;
rom[84219] = 12'h333;
rom[84220] = 12'h333;
rom[84221] = 12'h333;
rom[84222] = 12'h222;
rom[84223] = 12'h222;
rom[84224] = 12'h222;
rom[84225] = 12'h222;
rom[84226] = 12'h222;
rom[84227] = 12'h222;
rom[84228] = 12'h111;
rom[84229] = 12'h111;
rom[84230] = 12'h111;
rom[84231] = 12'h111;
rom[84232] = 12'h  0;
rom[84233] = 12'h  0;
rom[84234] = 12'h  0;
rom[84235] = 12'h  0;
rom[84236] = 12'h  0;
rom[84237] = 12'h  0;
rom[84238] = 12'h  0;
rom[84239] = 12'h  0;
rom[84240] = 12'h  0;
rom[84241] = 12'h  0;
rom[84242] = 12'h  0;
rom[84243] = 12'h  0;
rom[84244] = 12'h  0;
rom[84245] = 12'h  0;
rom[84246] = 12'h111;
rom[84247] = 12'h111;
rom[84248] = 12'h  0;
rom[84249] = 12'h  0;
rom[84250] = 12'h  0;
rom[84251] = 12'h  0;
rom[84252] = 12'h111;
rom[84253] = 12'h111;
rom[84254] = 12'h111;
rom[84255] = 12'h111;
rom[84256] = 12'h111;
rom[84257] = 12'h111;
rom[84258] = 12'h111;
rom[84259] = 12'h111;
rom[84260] = 12'h111;
rom[84261] = 12'h111;
rom[84262] = 12'h111;
rom[84263] = 12'h111;
rom[84264] = 12'h111;
rom[84265] = 12'h111;
rom[84266] = 12'h111;
rom[84267] = 12'h111;
rom[84268] = 12'h222;
rom[84269] = 12'h222;
rom[84270] = 12'h222;
rom[84271] = 12'h222;
rom[84272] = 12'h222;
rom[84273] = 12'h222;
rom[84274] = 12'h333;
rom[84275] = 12'h333;
rom[84276] = 12'h333;
rom[84277] = 12'h333;
rom[84278] = 12'h444;
rom[84279] = 12'h444;
rom[84280] = 12'h777;
rom[84281] = 12'h999;
rom[84282] = 12'haaa;
rom[84283] = 12'h888;
rom[84284] = 12'h777;
rom[84285] = 12'h777;
rom[84286] = 12'h777;
rom[84287] = 12'h666;
rom[84288] = 12'h666;
rom[84289] = 12'h666;
rom[84290] = 12'h666;
rom[84291] = 12'h666;
rom[84292] = 12'h666;
rom[84293] = 12'h666;
rom[84294] = 12'h666;
rom[84295] = 12'h666;
rom[84296] = 12'h666;
rom[84297] = 12'h666;
rom[84298] = 12'h777;
rom[84299] = 12'h777;
rom[84300] = 12'h888;
rom[84301] = 12'h888;
rom[84302] = 12'h888;
rom[84303] = 12'h777;
rom[84304] = 12'h777;
rom[84305] = 12'h999;
rom[84306] = 12'haaa;
rom[84307] = 12'hbbb;
rom[84308] = 12'hbbb;
rom[84309] = 12'hbbb;
rom[84310] = 12'haaa;
rom[84311] = 12'h999;
rom[84312] = 12'h888;
rom[84313] = 12'h888;
rom[84314] = 12'h888;
rom[84315] = 12'h777;
rom[84316] = 12'h777;
rom[84317] = 12'h777;
rom[84318] = 12'h777;
rom[84319] = 12'h777;
rom[84320] = 12'h777;
rom[84321] = 12'h777;
rom[84322] = 12'h777;
rom[84323] = 12'h777;
rom[84324] = 12'h888;
rom[84325] = 12'h888;
rom[84326] = 12'h888;
rom[84327] = 12'h888;
rom[84328] = 12'h888;
rom[84329] = 12'h888;
rom[84330] = 12'h777;
rom[84331] = 12'h777;
rom[84332] = 12'h777;
rom[84333] = 12'h666;
rom[84334] = 12'h666;
rom[84335] = 12'h666;
rom[84336] = 12'h555;
rom[84337] = 12'h555;
rom[84338] = 12'h555;
rom[84339] = 12'h555;
rom[84340] = 12'h555;
rom[84341] = 12'h555;
rom[84342] = 12'h555;
rom[84343] = 12'h555;
rom[84344] = 12'h444;
rom[84345] = 12'h444;
rom[84346] = 12'h444;
rom[84347] = 12'h333;
rom[84348] = 12'h333;
rom[84349] = 12'h333;
rom[84350] = 12'h333;
rom[84351] = 12'h333;
rom[84352] = 12'h333;
rom[84353] = 12'h333;
rom[84354] = 12'h444;
rom[84355] = 12'h444;
rom[84356] = 12'h444;
rom[84357] = 12'h444;
rom[84358] = 12'h444;
rom[84359] = 12'h444;
rom[84360] = 12'h444;
rom[84361] = 12'h444;
rom[84362] = 12'h444;
rom[84363] = 12'h444;
rom[84364] = 12'h444;
rom[84365] = 12'h333;
rom[84366] = 12'h333;
rom[84367] = 12'h444;
rom[84368] = 12'h333;
rom[84369] = 12'h333;
rom[84370] = 12'h333;
rom[84371] = 12'h333;
rom[84372] = 12'h333;
rom[84373] = 12'h333;
rom[84374] = 12'h333;
rom[84375] = 12'h333;
rom[84376] = 12'h333;
rom[84377] = 12'h333;
rom[84378] = 12'h333;
rom[84379] = 12'h333;
rom[84380] = 12'h222;
rom[84381] = 12'h222;
rom[84382] = 12'h222;
rom[84383] = 12'h222;
rom[84384] = 12'h222;
rom[84385] = 12'h222;
rom[84386] = 12'h222;
rom[84387] = 12'h222;
rom[84388] = 12'h222;
rom[84389] = 12'h222;
rom[84390] = 12'h222;
rom[84391] = 12'h222;
rom[84392] = 12'h222;
rom[84393] = 12'h222;
rom[84394] = 12'h222;
rom[84395] = 12'h111;
rom[84396] = 12'h111;
rom[84397] = 12'h111;
rom[84398] = 12'h111;
rom[84399] = 12'h111;
rom[84400] = 12'hfff;
rom[84401] = 12'hfff;
rom[84402] = 12'hfff;
rom[84403] = 12'hfff;
rom[84404] = 12'hfff;
rom[84405] = 12'hfff;
rom[84406] = 12'hfff;
rom[84407] = 12'hfff;
rom[84408] = 12'hfff;
rom[84409] = 12'hfff;
rom[84410] = 12'hfff;
rom[84411] = 12'hfff;
rom[84412] = 12'hfff;
rom[84413] = 12'hfff;
rom[84414] = 12'hfff;
rom[84415] = 12'hfff;
rom[84416] = 12'hfff;
rom[84417] = 12'hfff;
rom[84418] = 12'hfff;
rom[84419] = 12'hfff;
rom[84420] = 12'hfff;
rom[84421] = 12'hfff;
rom[84422] = 12'hfff;
rom[84423] = 12'hfff;
rom[84424] = 12'hfff;
rom[84425] = 12'hfff;
rom[84426] = 12'hfff;
rom[84427] = 12'hfff;
rom[84428] = 12'hfff;
rom[84429] = 12'hfff;
rom[84430] = 12'hfff;
rom[84431] = 12'hfff;
rom[84432] = 12'hfff;
rom[84433] = 12'hfff;
rom[84434] = 12'hfff;
rom[84435] = 12'hfff;
rom[84436] = 12'hfff;
rom[84437] = 12'hfff;
rom[84438] = 12'hfff;
rom[84439] = 12'hfff;
rom[84440] = 12'hfff;
rom[84441] = 12'hfff;
rom[84442] = 12'hfff;
rom[84443] = 12'hfff;
rom[84444] = 12'hfff;
rom[84445] = 12'hfff;
rom[84446] = 12'hfff;
rom[84447] = 12'hfff;
rom[84448] = 12'hfff;
rom[84449] = 12'hfff;
rom[84450] = 12'hfff;
rom[84451] = 12'hfff;
rom[84452] = 12'hfff;
rom[84453] = 12'hfff;
rom[84454] = 12'hfff;
rom[84455] = 12'hfff;
rom[84456] = 12'hfff;
rom[84457] = 12'hfff;
rom[84458] = 12'hfff;
rom[84459] = 12'hfff;
rom[84460] = 12'hfff;
rom[84461] = 12'hfff;
rom[84462] = 12'hfff;
rom[84463] = 12'hfff;
rom[84464] = 12'hfff;
rom[84465] = 12'hfff;
rom[84466] = 12'hfff;
rom[84467] = 12'hfff;
rom[84468] = 12'hfff;
rom[84469] = 12'hfff;
rom[84470] = 12'hfff;
rom[84471] = 12'hfff;
rom[84472] = 12'hfff;
rom[84473] = 12'hfff;
rom[84474] = 12'hfff;
rom[84475] = 12'hfff;
rom[84476] = 12'hfff;
rom[84477] = 12'hfff;
rom[84478] = 12'hfff;
rom[84479] = 12'hfff;
rom[84480] = 12'hfff;
rom[84481] = 12'hfff;
rom[84482] = 12'hfff;
rom[84483] = 12'hfff;
rom[84484] = 12'hfff;
rom[84485] = 12'hfff;
rom[84486] = 12'hfff;
rom[84487] = 12'hfff;
rom[84488] = 12'hfff;
rom[84489] = 12'hfff;
rom[84490] = 12'hfff;
rom[84491] = 12'hfff;
rom[84492] = 12'hfff;
rom[84493] = 12'hfff;
rom[84494] = 12'hfff;
rom[84495] = 12'hfff;
rom[84496] = 12'hfff;
rom[84497] = 12'hfff;
rom[84498] = 12'hfff;
rom[84499] = 12'hfff;
rom[84500] = 12'hfff;
rom[84501] = 12'hfff;
rom[84502] = 12'hfff;
rom[84503] = 12'hfff;
rom[84504] = 12'hfff;
rom[84505] = 12'hfff;
rom[84506] = 12'hfff;
rom[84507] = 12'hfff;
rom[84508] = 12'hfff;
rom[84509] = 12'hfff;
rom[84510] = 12'hfff;
rom[84511] = 12'hfff;
rom[84512] = 12'hfff;
rom[84513] = 12'hfff;
rom[84514] = 12'hfff;
rom[84515] = 12'hfff;
rom[84516] = 12'hfff;
rom[84517] = 12'hfff;
rom[84518] = 12'hfff;
rom[84519] = 12'hfff;
rom[84520] = 12'hfff;
rom[84521] = 12'hfff;
rom[84522] = 12'hfff;
rom[84523] = 12'hfff;
rom[84524] = 12'heee;
rom[84525] = 12'heee;
rom[84526] = 12'heee;
rom[84527] = 12'heee;
rom[84528] = 12'heee;
rom[84529] = 12'heee;
rom[84530] = 12'heee;
rom[84531] = 12'heee;
rom[84532] = 12'hddd;
rom[84533] = 12'hddd;
rom[84534] = 12'hddd;
rom[84535] = 12'hddd;
rom[84536] = 12'hddd;
rom[84537] = 12'hddd;
rom[84538] = 12'hddd;
rom[84539] = 12'hddd;
rom[84540] = 12'hddd;
rom[84541] = 12'hddd;
rom[84542] = 12'hddd;
rom[84543] = 12'hddd;
rom[84544] = 12'hddd;
rom[84545] = 12'hddd;
rom[84546] = 12'hccc;
rom[84547] = 12'hccc;
rom[84548] = 12'hbbb;
rom[84549] = 12'hbbb;
rom[84550] = 12'haaa;
rom[84551] = 12'haaa;
rom[84552] = 12'h999;
rom[84553] = 12'h888;
rom[84554] = 12'h888;
rom[84555] = 12'h777;
rom[84556] = 12'h777;
rom[84557] = 12'h666;
rom[84558] = 12'h666;
rom[84559] = 12'h555;
rom[84560] = 12'h555;
rom[84561] = 12'h555;
rom[84562] = 12'h555;
rom[84563] = 12'h444;
rom[84564] = 12'h444;
rom[84565] = 12'h444;
rom[84566] = 12'h444;
rom[84567] = 12'h444;
rom[84568] = 12'h444;
rom[84569] = 12'h444;
rom[84570] = 12'h444;
rom[84571] = 12'h444;
rom[84572] = 12'h444;
rom[84573] = 12'h444;
rom[84574] = 12'h444;
rom[84575] = 12'h444;
rom[84576] = 12'h444;
rom[84577] = 12'h444;
rom[84578] = 12'h444;
rom[84579] = 12'h444;
rom[84580] = 12'h555;
rom[84581] = 12'h555;
rom[84582] = 12'h555;
rom[84583] = 12'h555;
rom[84584] = 12'h555;
rom[84585] = 12'h555;
rom[84586] = 12'h555;
rom[84587] = 12'h555;
rom[84588] = 12'h555;
rom[84589] = 12'h555;
rom[84590] = 12'h555;
rom[84591] = 12'h555;
rom[84592] = 12'h444;
rom[84593] = 12'h444;
rom[84594] = 12'h444;
rom[84595] = 12'h333;
rom[84596] = 12'h333;
rom[84597] = 12'h444;
rom[84598] = 12'h444;
rom[84599] = 12'h444;
rom[84600] = 12'h444;
rom[84601] = 12'h444;
rom[84602] = 12'h444;
rom[84603] = 12'h444;
rom[84604] = 12'h555;
rom[84605] = 12'h666;
rom[84606] = 12'h666;
rom[84607] = 12'h666;
rom[84608] = 12'h555;
rom[84609] = 12'h666;
rom[84610] = 12'h777;
rom[84611] = 12'h888;
rom[84612] = 12'h999;
rom[84613] = 12'h999;
rom[84614] = 12'h777;
rom[84615] = 12'h777;
rom[84616] = 12'h666;
rom[84617] = 12'h555;
rom[84618] = 12'h444;
rom[84619] = 12'h333;
rom[84620] = 12'h333;
rom[84621] = 12'h333;
rom[84622] = 12'h222;
rom[84623] = 12'h222;
rom[84624] = 12'h222;
rom[84625] = 12'h222;
rom[84626] = 12'h111;
rom[84627] = 12'h111;
rom[84628] = 12'h111;
rom[84629] = 12'h111;
rom[84630] = 12'h111;
rom[84631] = 12'h111;
rom[84632] = 12'h  0;
rom[84633] = 12'h  0;
rom[84634] = 12'h  0;
rom[84635] = 12'h  0;
rom[84636] = 12'h  0;
rom[84637] = 12'h  0;
rom[84638] = 12'h  0;
rom[84639] = 12'h  0;
rom[84640] = 12'h  0;
rom[84641] = 12'h  0;
rom[84642] = 12'h  0;
rom[84643] = 12'h  0;
rom[84644] = 12'h  0;
rom[84645] = 12'h  0;
rom[84646] = 12'h  0;
rom[84647] = 12'h  0;
rom[84648] = 12'h  0;
rom[84649] = 12'h  0;
rom[84650] = 12'h  0;
rom[84651] = 12'h  0;
rom[84652] = 12'h  0;
rom[84653] = 12'h111;
rom[84654] = 12'h111;
rom[84655] = 12'h111;
rom[84656] = 12'h111;
rom[84657] = 12'h111;
rom[84658] = 12'h111;
rom[84659] = 12'h111;
rom[84660] = 12'h111;
rom[84661] = 12'h111;
rom[84662] = 12'h111;
rom[84663] = 12'h111;
rom[84664] = 12'h111;
rom[84665] = 12'h111;
rom[84666] = 12'h222;
rom[84667] = 12'h222;
rom[84668] = 12'h222;
rom[84669] = 12'h222;
rom[84670] = 12'h222;
rom[84671] = 12'h333;
rom[84672] = 12'h222;
rom[84673] = 12'h333;
rom[84674] = 12'h333;
rom[84675] = 12'h333;
rom[84676] = 12'h333;
rom[84677] = 12'h333;
rom[84678] = 12'h444;
rom[84679] = 12'h444;
rom[84680] = 12'h777;
rom[84681] = 12'h999;
rom[84682] = 12'haaa;
rom[84683] = 12'h999;
rom[84684] = 12'h777;
rom[84685] = 12'h777;
rom[84686] = 12'h777;
rom[84687] = 12'h777;
rom[84688] = 12'h666;
rom[84689] = 12'h666;
rom[84690] = 12'h666;
rom[84691] = 12'h666;
rom[84692] = 12'h666;
rom[84693] = 12'h666;
rom[84694] = 12'h666;
rom[84695] = 12'h666;
rom[84696] = 12'h666;
rom[84697] = 12'h666;
rom[84698] = 12'h777;
rom[84699] = 12'h777;
rom[84700] = 12'h888;
rom[84701] = 12'h888;
rom[84702] = 12'h888;
rom[84703] = 12'h888;
rom[84704] = 12'h888;
rom[84705] = 12'h999;
rom[84706] = 12'hbbb;
rom[84707] = 12'hbbb;
rom[84708] = 12'hbbb;
rom[84709] = 12'hbbb;
rom[84710] = 12'haaa;
rom[84711] = 12'h999;
rom[84712] = 12'h999;
rom[84713] = 12'h999;
rom[84714] = 12'h999;
rom[84715] = 12'h999;
rom[84716] = 12'h888;
rom[84717] = 12'h888;
rom[84718] = 12'h888;
rom[84719] = 12'h888;
rom[84720] = 12'h888;
rom[84721] = 12'h777;
rom[84722] = 12'h777;
rom[84723] = 12'h777;
rom[84724] = 12'h777;
rom[84725] = 12'h888;
rom[84726] = 12'h888;
rom[84727] = 12'h888;
rom[84728] = 12'h888;
rom[84729] = 12'h888;
rom[84730] = 12'h888;
rom[84731] = 12'h888;
rom[84732] = 12'h777;
rom[84733] = 12'h777;
rom[84734] = 12'h777;
rom[84735] = 12'h666;
rom[84736] = 12'h666;
rom[84737] = 12'h666;
rom[84738] = 12'h666;
rom[84739] = 12'h555;
rom[84740] = 12'h555;
rom[84741] = 12'h555;
rom[84742] = 12'h555;
rom[84743] = 12'h555;
rom[84744] = 12'h444;
rom[84745] = 12'h444;
rom[84746] = 12'h444;
rom[84747] = 12'h333;
rom[84748] = 12'h333;
rom[84749] = 12'h333;
rom[84750] = 12'h333;
rom[84751] = 12'h333;
rom[84752] = 12'h333;
rom[84753] = 12'h444;
rom[84754] = 12'h444;
rom[84755] = 12'h444;
rom[84756] = 12'h444;
rom[84757] = 12'h444;
rom[84758] = 12'h444;
rom[84759] = 12'h444;
rom[84760] = 12'h444;
rom[84761] = 12'h444;
rom[84762] = 12'h444;
rom[84763] = 12'h444;
rom[84764] = 12'h444;
rom[84765] = 12'h444;
rom[84766] = 12'h444;
rom[84767] = 12'h444;
rom[84768] = 12'h333;
rom[84769] = 12'h333;
rom[84770] = 12'h333;
rom[84771] = 12'h333;
rom[84772] = 12'h333;
rom[84773] = 12'h333;
rom[84774] = 12'h333;
rom[84775] = 12'h333;
rom[84776] = 12'h333;
rom[84777] = 12'h333;
rom[84778] = 12'h333;
rom[84779] = 12'h333;
rom[84780] = 12'h222;
rom[84781] = 12'h222;
rom[84782] = 12'h222;
rom[84783] = 12'h222;
rom[84784] = 12'h222;
rom[84785] = 12'h222;
rom[84786] = 12'h222;
rom[84787] = 12'h222;
rom[84788] = 12'h222;
rom[84789] = 12'h222;
rom[84790] = 12'h222;
rom[84791] = 12'h222;
rom[84792] = 12'h222;
rom[84793] = 12'h222;
rom[84794] = 12'h222;
rom[84795] = 12'h111;
rom[84796] = 12'h111;
rom[84797] = 12'h111;
rom[84798] = 12'h111;
rom[84799] = 12'h111;
rom[84800] = 12'hfff;
rom[84801] = 12'hfff;
rom[84802] = 12'hfff;
rom[84803] = 12'hfff;
rom[84804] = 12'hfff;
rom[84805] = 12'hfff;
rom[84806] = 12'hfff;
rom[84807] = 12'hfff;
rom[84808] = 12'hfff;
rom[84809] = 12'hfff;
rom[84810] = 12'hfff;
rom[84811] = 12'hfff;
rom[84812] = 12'hfff;
rom[84813] = 12'hfff;
rom[84814] = 12'hfff;
rom[84815] = 12'hfff;
rom[84816] = 12'hfff;
rom[84817] = 12'hfff;
rom[84818] = 12'hfff;
rom[84819] = 12'hfff;
rom[84820] = 12'hfff;
rom[84821] = 12'hfff;
rom[84822] = 12'hfff;
rom[84823] = 12'hfff;
rom[84824] = 12'hfff;
rom[84825] = 12'hfff;
rom[84826] = 12'hfff;
rom[84827] = 12'hfff;
rom[84828] = 12'hfff;
rom[84829] = 12'hfff;
rom[84830] = 12'hfff;
rom[84831] = 12'hfff;
rom[84832] = 12'hfff;
rom[84833] = 12'hfff;
rom[84834] = 12'hfff;
rom[84835] = 12'hfff;
rom[84836] = 12'hfff;
rom[84837] = 12'hfff;
rom[84838] = 12'hfff;
rom[84839] = 12'hfff;
rom[84840] = 12'hfff;
rom[84841] = 12'hfff;
rom[84842] = 12'hfff;
rom[84843] = 12'hfff;
rom[84844] = 12'hfff;
rom[84845] = 12'hfff;
rom[84846] = 12'hfff;
rom[84847] = 12'hfff;
rom[84848] = 12'hfff;
rom[84849] = 12'hfff;
rom[84850] = 12'hfff;
rom[84851] = 12'hfff;
rom[84852] = 12'hfff;
rom[84853] = 12'hfff;
rom[84854] = 12'hfff;
rom[84855] = 12'hfff;
rom[84856] = 12'hfff;
rom[84857] = 12'hfff;
rom[84858] = 12'hfff;
rom[84859] = 12'hfff;
rom[84860] = 12'hfff;
rom[84861] = 12'hfff;
rom[84862] = 12'hfff;
rom[84863] = 12'hfff;
rom[84864] = 12'hfff;
rom[84865] = 12'hfff;
rom[84866] = 12'hfff;
rom[84867] = 12'hfff;
rom[84868] = 12'hfff;
rom[84869] = 12'hfff;
rom[84870] = 12'hfff;
rom[84871] = 12'hfff;
rom[84872] = 12'hfff;
rom[84873] = 12'hfff;
rom[84874] = 12'hfff;
rom[84875] = 12'hfff;
rom[84876] = 12'hfff;
rom[84877] = 12'hfff;
rom[84878] = 12'hfff;
rom[84879] = 12'hfff;
rom[84880] = 12'hfff;
rom[84881] = 12'hfff;
rom[84882] = 12'hfff;
rom[84883] = 12'hfff;
rom[84884] = 12'hfff;
rom[84885] = 12'hfff;
rom[84886] = 12'hfff;
rom[84887] = 12'hfff;
rom[84888] = 12'hfff;
rom[84889] = 12'hfff;
rom[84890] = 12'hfff;
rom[84891] = 12'hfff;
rom[84892] = 12'hfff;
rom[84893] = 12'hfff;
rom[84894] = 12'hfff;
rom[84895] = 12'hfff;
rom[84896] = 12'hfff;
rom[84897] = 12'hfff;
rom[84898] = 12'hfff;
rom[84899] = 12'hfff;
rom[84900] = 12'hfff;
rom[84901] = 12'hfff;
rom[84902] = 12'hfff;
rom[84903] = 12'hfff;
rom[84904] = 12'hfff;
rom[84905] = 12'hfff;
rom[84906] = 12'hfff;
rom[84907] = 12'hfff;
rom[84908] = 12'hfff;
rom[84909] = 12'hfff;
rom[84910] = 12'hfff;
rom[84911] = 12'hfff;
rom[84912] = 12'hfff;
rom[84913] = 12'hfff;
rom[84914] = 12'hfff;
rom[84915] = 12'hfff;
rom[84916] = 12'hfff;
rom[84917] = 12'hfff;
rom[84918] = 12'hfff;
rom[84919] = 12'hfff;
rom[84920] = 12'hfff;
rom[84921] = 12'hfff;
rom[84922] = 12'hfff;
rom[84923] = 12'hfff;
rom[84924] = 12'hfff;
rom[84925] = 12'heee;
rom[84926] = 12'heee;
rom[84927] = 12'heee;
rom[84928] = 12'heee;
rom[84929] = 12'heee;
rom[84930] = 12'hddd;
rom[84931] = 12'hddd;
rom[84932] = 12'hddd;
rom[84933] = 12'hddd;
rom[84934] = 12'hccc;
rom[84935] = 12'hccc;
rom[84936] = 12'hccc;
rom[84937] = 12'hccc;
rom[84938] = 12'hccc;
rom[84939] = 12'hddd;
rom[84940] = 12'hddd;
rom[84941] = 12'hddd;
rom[84942] = 12'hddd;
rom[84943] = 12'hddd;
rom[84944] = 12'hddd;
rom[84945] = 12'hddd;
rom[84946] = 12'hddd;
rom[84947] = 12'hccc;
rom[84948] = 12'hccc;
rom[84949] = 12'hbbb;
rom[84950] = 12'hbbb;
rom[84951] = 12'hbbb;
rom[84952] = 12'haaa;
rom[84953] = 12'haaa;
rom[84954] = 12'h999;
rom[84955] = 12'h888;
rom[84956] = 12'h888;
rom[84957] = 12'h777;
rom[84958] = 12'h666;
rom[84959] = 12'h666;
rom[84960] = 12'h666;
rom[84961] = 12'h555;
rom[84962] = 12'h555;
rom[84963] = 12'h555;
rom[84964] = 12'h555;
rom[84965] = 12'h555;
rom[84966] = 12'h555;
rom[84967] = 12'h444;
rom[84968] = 12'h444;
rom[84969] = 12'h444;
rom[84970] = 12'h444;
rom[84971] = 12'h444;
rom[84972] = 12'h444;
rom[84973] = 12'h444;
rom[84974] = 12'h444;
rom[84975] = 12'h444;
rom[84976] = 12'h444;
rom[84977] = 12'h444;
rom[84978] = 12'h444;
rom[84979] = 12'h555;
rom[84980] = 12'h555;
rom[84981] = 12'h555;
rom[84982] = 12'h555;
rom[84983] = 12'h555;
rom[84984] = 12'h555;
rom[84985] = 12'h555;
rom[84986] = 12'h555;
rom[84987] = 12'h555;
rom[84988] = 12'h555;
rom[84989] = 12'h555;
rom[84990] = 12'h555;
rom[84991] = 12'h555;
rom[84992] = 12'h444;
rom[84993] = 12'h444;
rom[84994] = 12'h444;
rom[84995] = 12'h444;
rom[84996] = 12'h444;
rom[84997] = 12'h444;
rom[84998] = 12'h444;
rom[84999] = 12'h444;
rom[85000] = 12'h444;
rom[85001] = 12'h444;
rom[85002] = 12'h444;
rom[85003] = 12'h444;
rom[85004] = 12'h555;
rom[85005] = 12'h666;
rom[85006] = 12'h666;
rom[85007] = 12'h666;
rom[85008] = 12'h555;
rom[85009] = 12'h555;
rom[85010] = 12'h666;
rom[85011] = 12'h777;
rom[85012] = 12'h888;
rom[85013] = 12'h888;
rom[85014] = 12'h888;
rom[85015] = 12'h888;
rom[85016] = 12'h777;
rom[85017] = 12'h555;
rom[85018] = 12'h444;
rom[85019] = 12'h333;
rom[85020] = 12'h333;
rom[85021] = 12'h333;
rom[85022] = 12'h222;
rom[85023] = 12'h222;
rom[85024] = 12'h222;
rom[85025] = 12'h222;
rom[85026] = 12'h111;
rom[85027] = 12'h111;
rom[85028] = 12'h111;
rom[85029] = 12'h111;
rom[85030] = 12'h111;
rom[85031] = 12'h111;
rom[85032] = 12'h  0;
rom[85033] = 12'h  0;
rom[85034] = 12'h  0;
rom[85035] = 12'h  0;
rom[85036] = 12'h  0;
rom[85037] = 12'h  0;
rom[85038] = 12'h  0;
rom[85039] = 12'h  0;
rom[85040] = 12'h  0;
rom[85041] = 12'h  0;
rom[85042] = 12'h  0;
rom[85043] = 12'h  0;
rom[85044] = 12'h  0;
rom[85045] = 12'h  0;
rom[85046] = 12'h  0;
rom[85047] = 12'h  0;
rom[85048] = 12'h  0;
rom[85049] = 12'h  0;
rom[85050] = 12'h  0;
rom[85051] = 12'h  0;
rom[85052] = 12'h  0;
rom[85053] = 12'h  0;
rom[85054] = 12'h  0;
rom[85055] = 12'h  0;
rom[85056] = 12'h111;
rom[85057] = 12'h111;
rom[85058] = 12'h111;
rom[85059] = 12'h111;
rom[85060] = 12'h111;
rom[85061] = 12'h111;
rom[85062] = 12'h111;
rom[85063] = 12'h222;
rom[85064] = 12'h111;
rom[85065] = 12'h111;
rom[85066] = 12'h222;
rom[85067] = 12'h222;
rom[85068] = 12'h222;
rom[85069] = 12'h222;
rom[85070] = 12'h333;
rom[85071] = 12'h333;
rom[85072] = 12'h333;
rom[85073] = 12'h333;
rom[85074] = 12'h333;
rom[85075] = 12'h333;
rom[85076] = 12'h333;
rom[85077] = 12'h444;
rom[85078] = 12'h444;
rom[85079] = 12'h444;
rom[85080] = 12'h777;
rom[85081] = 12'h999;
rom[85082] = 12'haaa;
rom[85083] = 12'h999;
rom[85084] = 12'h888;
rom[85085] = 12'h777;
rom[85086] = 12'h777;
rom[85087] = 12'h777;
rom[85088] = 12'h666;
rom[85089] = 12'h666;
rom[85090] = 12'h666;
rom[85091] = 12'h666;
rom[85092] = 12'h666;
rom[85093] = 12'h666;
rom[85094] = 12'h666;
rom[85095] = 12'h666;
rom[85096] = 12'h777;
rom[85097] = 12'h777;
rom[85098] = 12'h777;
rom[85099] = 12'h777;
rom[85100] = 12'h888;
rom[85101] = 12'h888;
rom[85102] = 12'h888;
rom[85103] = 12'h888;
rom[85104] = 12'h999;
rom[85105] = 12'haaa;
rom[85106] = 12'hbbb;
rom[85107] = 12'hbbb;
rom[85108] = 12'hbbb;
rom[85109] = 12'hbbb;
rom[85110] = 12'hbbb;
rom[85111] = 12'hbbb;
rom[85112] = 12'hbbb;
rom[85113] = 12'hbbb;
rom[85114] = 12'hbbb;
rom[85115] = 12'hbbb;
rom[85116] = 12'haaa;
rom[85117] = 12'haaa;
rom[85118] = 12'h999;
rom[85119] = 12'h999;
rom[85120] = 12'h888;
rom[85121] = 12'h888;
rom[85122] = 12'h888;
rom[85123] = 12'h888;
rom[85124] = 12'h888;
rom[85125] = 12'h888;
rom[85126] = 12'h888;
rom[85127] = 12'h888;
rom[85128] = 12'h888;
rom[85129] = 12'h888;
rom[85130] = 12'h888;
rom[85131] = 12'h888;
rom[85132] = 12'h888;
rom[85133] = 12'h777;
rom[85134] = 12'h777;
rom[85135] = 12'h777;
rom[85136] = 12'h777;
rom[85137] = 12'h777;
rom[85138] = 12'h666;
rom[85139] = 12'h666;
rom[85140] = 12'h666;
rom[85141] = 12'h555;
rom[85142] = 12'h555;
rom[85143] = 12'h555;
rom[85144] = 12'h444;
rom[85145] = 12'h444;
rom[85146] = 12'h444;
rom[85147] = 12'h444;
rom[85148] = 12'h444;
rom[85149] = 12'h444;
rom[85150] = 12'h444;
rom[85151] = 12'h444;
rom[85152] = 12'h444;
rom[85153] = 12'h444;
rom[85154] = 12'h444;
rom[85155] = 12'h444;
rom[85156] = 12'h444;
rom[85157] = 12'h444;
rom[85158] = 12'h444;
rom[85159] = 12'h444;
rom[85160] = 12'h444;
rom[85161] = 12'h444;
rom[85162] = 12'h444;
rom[85163] = 12'h444;
rom[85164] = 12'h444;
rom[85165] = 12'h444;
rom[85166] = 12'h444;
rom[85167] = 12'h444;
rom[85168] = 12'h333;
rom[85169] = 12'h333;
rom[85170] = 12'h444;
rom[85171] = 12'h444;
rom[85172] = 12'h444;
rom[85173] = 12'h333;
rom[85174] = 12'h333;
rom[85175] = 12'h333;
rom[85176] = 12'h333;
rom[85177] = 12'h333;
rom[85178] = 12'h333;
rom[85179] = 12'h333;
rom[85180] = 12'h333;
rom[85181] = 12'h222;
rom[85182] = 12'h222;
rom[85183] = 12'h222;
rom[85184] = 12'h222;
rom[85185] = 12'h222;
rom[85186] = 12'h222;
rom[85187] = 12'h222;
rom[85188] = 12'h222;
rom[85189] = 12'h222;
rom[85190] = 12'h222;
rom[85191] = 12'h222;
rom[85192] = 12'h222;
rom[85193] = 12'h222;
rom[85194] = 12'h222;
rom[85195] = 12'h111;
rom[85196] = 12'h111;
rom[85197] = 12'h111;
rom[85198] = 12'h111;
rom[85199] = 12'h222;
rom[85200] = 12'hfff;
rom[85201] = 12'hfff;
rom[85202] = 12'hfff;
rom[85203] = 12'hfff;
rom[85204] = 12'hfff;
rom[85205] = 12'hfff;
rom[85206] = 12'hfff;
rom[85207] = 12'hfff;
rom[85208] = 12'hfff;
rom[85209] = 12'hfff;
rom[85210] = 12'hfff;
rom[85211] = 12'hfff;
rom[85212] = 12'hfff;
rom[85213] = 12'hfff;
rom[85214] = 12'hfff;
rom[85215] = 12'hfff;
rom[85216] = 12'hfff;
rom[85217] = 12'hfff;
rom[85218] = 12'hfff;
rom[85219] = 12'hfff;
rom[85220] = 12'hfff;
rom[85221] = 12'hfff;
rom[85222] = 12'hfff;
rom[85223] = 12'hfff;
rom[85224] = 12'hfff;
rom[85225] = 12'hfff;
rom[85226] = 12'hfff;
rom[85227] = 12'hfff;
rom[85228] = 12'hfff;
rom[85229] = 12'hfff;
rom[85230] = 12'hfff;
rom[85231] = 12'hfff;
rom[85232] = 12'hfff;
rom[85233] = 12'hfff;
rom[85234] = 12'hfff;
rom[85235] = 12'hfff;
rom[85236] = 12'hfff;
rom[85237] = 12'hfff;
rom[85238] = 12'hfff;
rom[85239] = 12'hfff;
rom[85240] = 12'hfff;
rom[85241] = 12'hfff;
rom[85242] = 12'hfff;
rom[85243] = 12'hfff;
rom[85244] = 12'hfff;
rom[85245] = 12'hfff;
rom[85246] = 12'hfff;
rom[85247] = 12'hfff;
rom[85248] = 12'hfff;
rom[85249] = 12'hfff;
rom[85250] = 12'hfff;
rom[85251] = 12'hfff;
rom[85252] = 12'hfff;
rom[85253] = 12'hfff;
rom[85254] = 12'hfff;
rom[85255] = 12'hfff;
rom[85256] = 12'hfff;
rom[85257] = 12'hfff;
rom[85258] = 12'hfff;
rom[85259] = 12'hfff;
rom[85260] = 12'hfff;
rom[85261] = 12'hfff;
rom[85262] = 12'hfff;
rom[85263] = 12'hfff;
rom[85264] = 12'hfff;
rom[85265] = 12'hfff;
rom[85266] = 12'hfff;
rom[85267] = 12'hfff;
rom[85268] = 12'hfff;
rom[85269] = 12'hfff;
rom[85270] = 12'hfff;
rom[85271] = 12'hfff;
rom[85272] = 12'hfff;
rom[85273] = 12'hfff;
rom[85274] = 12'hfff;
rom[85275] = 12'hfff;
rom[85276] = 12'hfff;
rom[85277] = 12'hfff;
rom[85278] = 12'hfff;
rom[85279] = 12'hfff;
rom[85280] = 12'hfff;
rom[85281] = 12'hfff;
rom[85282] = 12'hfff;
rom[85283] = 12'hfff;
rom[85284] = 12'hfff;
rom[85285] = 12'hfff;
rom[85286] = 12'hfff;
rom[85287] = 12'hfff;
rom[85288] = 12'hfff;
rom[85289] = 12'hfff;
rom[85290] = 12'hfff;
rom[85291] = 12'hfff;
rom[85292] = 12'hfff;
rom[85293] = 12'hfff;
rom[85294] = 12'hfff;
rom[85295] = 12'hfff;
rom[85296] = 12'hfff;
rom[85297] = 12'hfff;
rom[85298] = 12'hfff;
rom[85299] = 12'hfff;
rom[85300] = 12'hfff;
rom[85301] = 12'hfff;
rom[85302] = 12'hfff;
rom[85303] = 12'hfff;
rom[85304] = 12'hfff;
rom[85305] = 12'hfff;
rom[85306] = 12'hfff;
rom[85307] = 12'hfff;
rom[85308] = 12'hfff;
rom[85309] = 12'hfff;
rom[85310] = 12'hfff;
rom[85311] = 12'hfff;
rom[85312] = 12'hfff;
rom[85313] = 12'hfff;
rom[85314] = 12'hfff;
rom[85315] = 12'hfff;
rom[85316] = 12'hfff;
rom[85317] = 12'hfff;
rom[85318] = 12'hfff;
rom[85319] = 12'hfff;
rom[85320] = 12'hfff;
rom[85321] = 12'hfff;
rom[85322] = 12'hfff;
rom[85323] = 12'hfff;
rom[85324] = 12'hfff;
rom[85325] = 12'hfff;
rom[85326] = 12'heee;
rom[85327] = 12'heee;
rom[85328] = 12'heee;
rom[85329] = 12'hddd;
rom[85330] = 12'hddd;
rom[85331] = 12'hddd;
rom[85332] = 12'hccc;
rom[85333] = 12'hccc;
rom[85334] = 12'hccc;
rom[85335] = 12'hccc;
rom[85336] = 12'hbbb;
rom[85337] = 12'hbbb;
rom[85338] = 12'hbbb;
rom[85339] = 12'hbbb;
rom[85340] = 12'hccc;
rom[85341] = 12'hccc;
rom[85342] = 12'hccc;
rom[85343] = 12'hccc;
rom[85344] = 12'hddd;
rom[85345] = 12'hddd;
rom[85346] = 12'hddd;
rom[85347] = 12'hccc;
rom[85348] = 12'hccc;
rom[85349] = 12'hccc;
rom[85350] = 12'hccc;
rom[85351] = 12'hccc;
rom[85352] = 12'hbbb;
rom[85353] = 12'hbbb;
rom[85354] = 12'haaa;
rom[85355] = 12'h999;
rom[85356] = 12'h999;
rom[85357] = 12'h888;
rom[85358] = 12'h777;
rom[85359] = 12'h777;
rom[85360] = 12'h666;
rom[85361] = 12'h666;
rom[85362] = 12'h555;
rom[85363] = 12'h555;
rom[85364] = 12'h555;
rom[85365] = 12'h555;
rom[85366] = 12'h555;
rom[85367] = 12'h555;
rom[85368] = 12'h444;
rom[85369] = 12'h444;
rom[85370] = 12'h444;
rom[85371] = 12'h444;
rom[85372] = 12'h444;
rom[85373] = 12'h444;
rom[85374] = 12'h444;
rom[85375] = 12'h444;
rom[85376] = 12'h444;
rom[85377] = 12'h555;
rom[85378] = 12'h555;
rom[85379] = 12'h555;
rom[85380] = 12'h555;
rom[85381] = 12'h555;
rom[85382] = 12'h555;
rom[85383] = 12'h555;
rom[85384] = 12'h555;
rom[85385] = 12'h555;
rom[85386] = 12'h555;
rom[85387] = 12'h555;
rom[85388] = 12'h555;
rom[85389] = 12'h555;
rom[85390] = 12'h555;
rom[85391] = 12'h555;
rom[85392] = 12'h444;
rom[85393] = 12'h444;
rom[85394] = 12'h444;
rom[85395] = 12'h444;
rom[85396] = 12'h444;
rom[85397] = 12'h444;
rom[85398] = 12'h444;
rom[85399] = 12'h444;
rom[85400] = 12'h444;
rom[85401] = 12'h444;
rom[85402] = 12'h444;
rom[85403] = 12'h555;
rom[85404] = 12'h555;
rom[85405] = 12'h666;
rom[85406] = 12'h666;
rom[85407] = 12'h666;
rom[85408] = 12'h555;
rom[85409] = 12'h555;
rom[85410] = 12'h555;
rom[85411] = 12'h666;
rom[85412] = 12'h777;
rom[85413] = 12'h888;
rom[85414] = 12'h888;
rom[85415] = 12'h888;
rom[85416] = 12'h777;
rom[85417] = 12'h666;
rom[85418] = 12'h555;
rom[85419] = 12'h333;
rom[85420] = 12'h333;
rom[85421] = 12'h333;
rom[85422] = 12'h222;
rom[85423] = 12'h222;
rom[85424] = 12'h222;
rom[85425] = 12'h222;
rom[85426] = 12'h222;
rom[85427] = 12'h222;
rom[85428] = 12'h222;
rom[85429] = 12'h222;
rom[85430] = 12'h111;
rom[85431] = 12'h111;
rom[85432] = 12'h111;
rom[85433] = 12'h111;
rom[85434] = 12'h  0;
rom[85435] = 12'h  0;
rom[85436] = 12'h  0;
rom[85437] = 12'h  0;
rom[85438] = 12'h  0;
rom[85439] = 12'h  0;
rom[85440] = 12'h  0;
rom[85441] = 12'h  0;
rom[85442] = 12'h  0;
rom[85443] = 12'h  0;
rom[85444] = 12'h  0;
rom[85445] = 12'h  0;
rom[85446] = 12'h  0;
rom[85447] = 12'h  0;
rom[85448] = 12'h  0;
rom[85449] = 12'h  0;
rom[85450] = 12'h  0;
rom[85451] = 12'h  0;
rom[85452] = 12'h  0;
rom[85453] = 12'h  0;
rom[85454] = 12'h  0;
rom[85455] = 12'h  0;
rom[85456] = 12'h  0;
rom[85457] = 12'h111;
rom[85458] = 12'h111;
rom[85459] = 12'h111;
rom[85460] = 12'h111;
rom[85461] = 12'h111;
rom[85462] = 12'h111;
rom[85463] = 12'h111;
rom[85464] = 12'h111;
rom[85465] = 12'h111;
rom[85466] = 12'h222;
rom[85467] = 12'h222;
rom[85468] = 12'h222;
rom[85469] = 12'h222;
rom[85470] = 12'h222;
rom[85471] = 12'h333;
rom[85472] = 12'h333;
rom[85473] = 12'h333;
rom[85474] = 12'h333;
rom[85475] = 12'h333;
rom[85476] = 12'h333;
rom[85477] = 12'h444;
rom[85478] = 12'h444;
rom[85479] = 12'h444;
rom[85480] = 12'h777;
rom[85481] = 12'h888;
rom[85482] = 12'haaa;
rom[85483] = 12'h999;
rom[85484] = 12'h888;
rom[85485] = 12'h777;
rom[85486] = 12'h777;
rom[85487] = 12'h666;
rom[85488] = 12'h666;
rom[85489] = 12'h666;
rom[85490] = 12'h666;
rom[85491] = 12'h666;
rom[85492] = 12'h666;
rom[85493] = 12'h666;
rom[85494] = 12'h666;
rom[85495] = 12'h666;
rom[85496] = 12'h777;
rom[85497] = 12'h777;
rom[85498] = 12'h777;
rom[85499] = 12'h777;
rom[85500] = 12'h777;
rom[85501] = 12'h777;
rom[85502] = 12'h888;
rom[85503] = 12'h888;
rom[85504] = 12'haaa;
rom[85505] = 12'haaa;
rom[85506] = 12'hbbb;
rom[85507] = 12'hbbb;
rom[85508] = 12'haaa;
rom[85509] = 12'haaa;
rom[85510] = 12'hbbb;
rom[85511] = 12'hbbb;
rom[85512] = 12'hbbb;
rom[85513] = 12'hccc;
rom[85514] = 12'hddd;
rom[85515] = 12'hddd;
rom[85516] = 12'hddd;
rom[85517] = 12'hddd;
rom[85518] = 12'hccc;
rom[85519] = 12'hccc;
rom[85520] = 12'hccc;
rom[85521] = 12'hbbb;
rom[85522] = 12'hbbb;
rom[85523] = 12'haaa;
rom[85524] = 12'haaa;
rom[85525] = 12'haaa;
rom[85526] = 12'h999;
rom[85527] = 12'h999;
rom[85528] = 12'h999;
rom[85529] = 12'h999;
rom[85530] = 12'h999;
rom[85531] = 12'h999;
rom[85532] = 12'h888;
rom[85533] = 12'h888;
rom[85534] = 12'h777;
rom[85535] = 12'h777;
rom[85536] = 12'h777;
rom[85537] = 12'h777;
rom[85538] = 12'h666;
rom[85539] = 12'h666;
rom[85540] = 12'h666;
rom[85541] = 12'h666;
rom[85542] = 12'h555;
rom[85543] = 12'h555;
rom[85544] = 12'h555;
rom[85545] = 12'h444;
rom[85546] = 12'h444;
rom[85547] = 12'h444;
rom[85548] = 12'h444;
rom[85549] = 12'h444;
rom[85550] = 12'h444;
rom[85551] = 12'h444;
rom[85552] = 12'h444;
rom[85553] = 12'h444;
rom[85554] = 12'h444;
rom[85555] = 12'h444;
rom[85556] = 12'h444;
rom[85557] = 12'h444;
rom[85558] = 12'h444;
rom[85559] = 12'h444;
rom[85560] = 12'h444;
rom[85561] = 12'h444;
rom[85562] = 12'h444;
rom[85563] = 12'h444;
rom[85564] = 12'h444;
rom[85565] = 12'h444;
rom[85566] = 12'h444;
rom[85567] = 12'h444;
rom[85568] = 12'h444;
rom[85569] = 12'h444;
rom[85570] = 12'h444;
rom[85571] = 12'h444;
rom[85572] = 12'h444;
rom[85573] = 12'h333;
rom[85574] = 12'h333;
rom[85575] = 12'h333;
rom[85576] = 12'h333;
rom[85577] = 12'h333;
rom[85578] = 12'h333;
rom[85579] = 12'h333;
rom[85580] = 12'h333;
rom[85581] = 12'h333;
rom[85582] = 12'h222;
rom[85583] = 12'h222;
rom[85584] = 12'h222;
rom[85585] = 12'h222;
rom[85586] = 12'h222;
rom[85587] = 12'h222;
rom[85588] = 12'h222;
rom[85589] = 12'h222;
rom[85590] = 12'h222;
rom[85591] = 12'h222;
rom[85592] = 12'h222;
rom[85593] = 12'h222;
rom[85594] = 12'h222;
rom[85595] = 12'h222;
rom[85596] = 12'h222;
rom[85597] = 12'h222;
rom[85598] = 12'h222;
rom[85599] = 12'h222;
rom[85600] = 12'hfff;
rom[85601] = 12'hfff;
rom[85602] = 12'hfff;
rom[85603] = 12'hfff;
rom[85604] = 12'hfff;
rom[85605] = 12'hfff;
rom[85606] = 12'hfff;
rom[85607] = 12'hfff;
rom[85608] = 12'hfff;
rom[85609] = 12'hfff;
rom[85610] = 12'hfff;
rom[85611] = 12'hfff;
rom[85612] = 12'hfff;
rom[85613] = 12'hfff;
rom[85614] = 12'hfff;
rom[85615] = 12'hfff;
rom[85616] = 12'hfff;
rom[85617] = 12'hfff;
rom[85618] = 12'hfff;
rom[85619] = 12'hfff;
rom[85620] = 12'hfff;
rom[85621] = 12'hfff;
rom[85622] = 12'hfff;
rom[85623] = 12'hfff;
rom[85624] = 12'hfff;
rom[85625] = 12'hfff;
rom[85626] = 12'hfff;
rom[85627] = 12'hfff;
rom[85628] = 12'hfff;
rom[85629] = 12'hfff;
rom[85630] = 12'hfff;
rom[85631] = 12'hfff;
rom[85632] = 12'hfff;
rom[85633] = 12'hfff;
rom[85634] = 12'hfff;
rom[85635] = 12'hfff;
rom[85636] = 12'hfff;
rom[85637] = 12'hfff;
rom[85638] = 12'hfff;
rom[85639] = 12'hfff;
rom[85640] = 12'hfff;
rom[85641] = 12'hfff;
rom[85642] = 12'hfff;
rom[85643] = 12'hfff;
rom[85644] = 12'hfff;
rom[85645] = 12'hfff;
rom[85646] = 12'hfff;
rom[85647] = 12'hfff;
rom[85648] = 12'hfff;
rom[85649] = 12'hfff;
rom[85650] = 12'hfff;
rom[85651] = 12'hfff;
rom[85652] = 12'hfff;
rom[85653] = 12'hfff;
rom[85654] = 12'hfff;
rom[85655] = 12'hfff;
rom[85656] = 12'hfff;
rom[85657] = 12'hfff;
rom[85658] = 12'hfff;
rom[85659] = 12'hfff;
rom[85660] = 12'hfff;
rom[85661] = 12'hfff;
rom[85662] = 12'hfff;
rom[85663] = 12'hfff;
rom[85664] = 12'hfff;
rom[85665] = 12'hfff;
rom[85666] = 12'hfff;
rom[85667] = 12'hfff;
rom[85668] = 12'hfff;
rom[85669] = 12'hfff;
rom[85670] = 12'hfff;
rom[85671] = 12'hfff;
rom[85672] = 12'hfff;
rom[85673] = 12'hfff;
rom[85674] = 12'hfff;
rom[85675] = 12'hfff;
rom[85676] = 12'hfff;
rom[85677] = 12'hfff;
rom[85678] = 12'hfff;
rom[85679] = 12'hfff;
rom[85680] = 12'hfff;
rom[85681] = 12'hfff;
rom[85682] = 12'hfff;
rom[85683] = 12'hfff;
rom[85684] = 12'hfff;
rom[85685] = 12'hfff;
rom[85686] = 12'hfff;
rom[85687] = 12'hfff;
rom[85688] = 12'hfff;
rom[85689] = 12'hfff;
rom[85690] = 12'hfff;
rom[85691] = 12'hfff;
rom[85692] = 12'hfff;
rom[85693] = 12'hfff;
rom[85694] = 12'hfff;
rom[85695] = 12'hfff;
rom[85696] = 12'hfff;
rom[85697] = 12'hfff;
rom[85698] = 12'hfff;
rom[85699] = 12'hfff;
rom[85700] = 12'hfff;
rom[85701] = 12'hfff;
rom[85702] = 12'hfff;
rom[85703] = 12'hfff;
rom[85704] = 12'hfff;
rom[85705] = 12'hfff;
rom[85706] = 12'hfff;
rom[85707] = 12'hfff;
rom[85708] = 12'hfff;
rom[85709] = 12'hfff;
rom[85710] = 12'hfff;
rom[85711] = 12'hfff;
rom[85712] = 12'hfff;
rom[85713] = 12'hfff;
rom[85714] = 12'hfff;
rom[85715] = 12'hfff;
rom[85716] = 12'hfff;
rom[85717] = 12'hfff;
rom[85718] = 12'hfff;
rom[85719] = 12'hfff;
rom[85720] = 12'hfff;
rom[85721] = 12'hfff;
rom[85722] = 12'hfff;
rom[85723] = 12'hfff;
rom[85724] = 12'hfff;
rom[85725] = 12'heee;
rom[85726] = 12'heee;
rom[85727] = 12'heee;
rom[85728] = 12'hddd;
rom[85729] = 12'hddd;
rom[85730] = 12'hddd;
rom[85731] = 12'hccc;
rom[85732] = 12'hccc;
rom[85733] = 12'hccc;
rom[85734] = 12'hccc;
rom[85735] = 12'hccc;
rom[85736] = 12'hbbb;
rom[85737] = 12'hbbb;
rom[85738] = 12'hbbb;
rom[85739] = 12'hbbb;
rom[85740] = 12'hbbb;
rom[85741] = 12'hbbb;
rom[85742] = 12'hbbb;
rom[85743] = 12'hbbb;
rom[85744] = 12'hbbb;
rom[85745] = 12'hbbb;
rom[85746] = 12'hbbb;
rom[85747] = 12'hccc;
rom[85748] = 12'hccc;
rom[85749] = 12'hccc;
rom[85750] = 12'hccc;
rom[85751] = 12'hccc;
rom[85752] = 12'hbbb;
rom[85753] = 12'hbbb;
rom[85754] = 12'hbbb;
rom[85755] = 12'haaa;
rom[85756] = 12'haaa;
rom[85757] = 12'h999;
rom[85758] = 12'h999;
rom[85759] = 12'h888;
rom[85760] = 12'h777;
rom[85761] = 12'h777;
rom[85762] = 12'h666;
rom[85763] = 12'h666;
rom[85764] = 12'h666;
rom[85765] = 12'h666;
rom[85766] = 12'h666;
rom[85767] = 12'h666;
rom[85768] = 12'h555;
rom[85769] = 12'h555;
rom[85770] = 12'h555;
rom[85771] = 12'h555;
rom[85772] = 12'h555;
rom[85773] = 12'h555;
rom[85774] = 12'h555;
rom[85775] = 12'h555;
rom[85776] = 12'h555;
rom[85777] = 12'h555;
rom[85778] = 12'h555;
rom[85779] = 12'h555;
rom[85780] = 12'h555;
rom[85781] = 12'h555;
rom[85782] = 12'h555;
rom[85783] = 12'h555;
rom[85784] = 12'h555;
rom[85785] = 12'h555;
rom[85786] = 12'h555;
rom[85787] = 12'h555;
rom[85788] = 12'h555;
rom[85789] = 12'h555;
rom[85790] = 12'h555;
rom[85791] = 12'h555;
rom[85792] = 12'h555;
rom[85793] = 12'h444;
rom[85794] = 12'h444;
rom[85795] = 12'h444;
rom[85796] = 12'h444;
rom[85797] = 12'h444;
rom[85798] = 12'h444;
rom[85799] = 12'h444;
rom[85800] = 12'h444;
rom[85801] = 12'h444;
rom[85802] = 12'h555;
rom[85803] = 12'h555;
rom[85804] = 12'h555;
rom[85805] = 12'h555;
rom[85806] = 12'h555;
rom[85807] = 12'h555;
rom[85808] = 12'h555;
rom[85809] = 12'h555;
rom[85810] = 12'h555;
rom[85811] = 12'h555;
rom[85812] = 12'h666;
rom[85813] = 12'h777;
rom[85814] = 12'h888;
rom[85815] = 12'h888;
rom[85816] = 12'h777;
rom[85817] = 12'h777;
rom[85818] = 12'h666;
rom[85819] = 12'h444;
rom[85820] = 12'h444;
rom[85821] = 12'h333;
rom[85822] = 12'h333;
rom[85823] = 12'h222;
rom[85824] = 12'h222;
rom[85825] = 12'h222;
rom[85826] = 12'h222;
rom[85827] = 12'h222;
rom[85828] = 12'h222;
rom[85829] = 12'h222;
rom[85830] = 12'h111;
rom[85831] = 12'h111;
rom[85832] = 12'h111;
rom[85833] = 12'h111;
rom[85834] = 12'h111;
rom[85835] = 12'h  0;
rom[85836] = 12'h  0;
rom[85837] = 12'h  0;
rom[85838] = 12'h  0;
rom[85839] = 12'h  0;
rom[85840] = 12'h  0;
rom[85841] = 12'h  0;
rom[85842] = 12'h  0;
rom[85843] = 12'h  0;
rom[85844] = 12'h  0;
rom[85845] = 12'h  0;
rom[85846] = 12'h  0;
rom[85847] = 12'h  0;
rom[85848] = 12'h  0;
rom[85849] = 12'h  0;
rom[85850] = 12'h  0;
rom[85851] = 12'h  0;
rom[85852] = 12'h  0;
rom[85853] = 12'h  0;
rom[85854] = 12'h  0;
rom[85855] = 12'h  0;
rom[85856] = 12'h  0;
rom[85857] = 12'h  0;
rom[85858] = 12'h  0;
rom[85859] = 12'h  0;
rom[85860] = 12'h111;
rom[85861] = 12'h111;
rom[85862] = 12'h111;
rom[85863] = 12'h111;
rom[85864] = 12'h111;
rom[85865] = 12'h111;
rom[85866] = 12'h111;
rom[85867] = 12'h111;
rom[85868] = 12'h222;
rom[85869] = 12'h222;
rom[85870] = 12'h222;
rom[85871] = 12'h222;
rom[85872] = 12'h222;
rom[85873] = 12'h333;
rom[85874] = 12'h333;
rom[85875] = 12'h333;
rom[85876] = 12'h333;
rom[85877] = 12'h333;
rom[85878] = 12'h444;
rom[85879] = 12'h444;
rom[85880] = 12'h666;
rom[85881] = 12'h888;
rom[85882] = 12'h999;
rom[85883] = 12'h999;
rom[85884] = 12'h888;
rom[85885] = 12'h777;
rom[85886] = 12'h777;
rom[85887] = 12'h666;
rom[85888] = 12'h666;
rom[85889] = 12'h666;
rom[85890] = 12'h666;
rom[85891] = 12'h666;
rom[85892] = 12'h666;
rom[85893] = 12'h666;
rom[85894] = 12'h666;
rom[85895] = 12'h666;
rom[85896] = 12'h666;
rom[85897] = 12'h777;
rom[85898] = 12'h777;
rom[85899] = 12'h777;
rom[85900] = 12'h777;
rom[85901] = 12'h777;
rom[85902] = 12'h777;
rom[85903] = 12'h888;
rom[85904] = 12'haaa;
rom[85905] = 12'haaa;
rom[85906] = 12'hbbb;
rom[85907] = 12'haaa;
rom[85908] = 12'h999;
rom[85909] = 12'h999;
rom[85910] = 12'h999;
rom[85911] = 12'h999;
rom[85912] = 12'h999;
rom[85913] = 12'haaa;
rom[85914] = 12'hbbb;
rom[85915] = 12'hbbb;
rom[85916] = 12'hccc;
rom[85917] = 12'hddd;
rom[85918] = 12'hddd;
rom[85919] = 12'heee;
rom[85920] = 12'heee;
rom[85921] = 12'heee;
rom[85922] = 12'heee;
rom[85923] = 12'heee;
rom[85924] = 12'hddd;
rom[85925] = 12'hddd;
rom[85926] = 12'hccc;
rom[85927] = 12'hccc;
rom[85928] = 12'hbbb;
rom[85929] = 12'hbbb;
rom[85930] = 12'hbbb;
rom[85931] = 12'hbbb;
rom[85932] = 12'hbbb;
rom[85933] = 12'haaa;
rom[85934] = 12'h999;
rom[85935] = 12'h999;
rom[85936] = 12'h888;
rom[85937] = 12'h888;
rom[85938] = 12'h777;
rom[85939] = 12'h777;
rom[85940] = 12'h777;
rom[85941] = 12'h777;
rom[85942] = 12'h666;
rom[85943] = 12'h555;
rom[85944] = 12'h555;
rom[85945] = 12'h555;
rom[85946] = 12'h555;
rom[85947] = 12'h555;
rom[85948] = 12'h444;
rom[85949] = 12'h444;
rom[85950] = 12'h555;
rom[85951] = 12'h555;
rom[85952] = 12'h555;
rom[85953] = 12'h555;
rom[85954] = 12'h555;
rom[85955] = 12'h555;
rom[85956] = 12'h555;
rom[85957] = 12'h555;
rom[85958] = 12'h444;
rom[85959] = 12'h444;
rom[85960] = 12'h444;
rom[85961] = 12'h444;
rom[85962] = 12'h444;
rom[85963] = 12'h444;
rom[85964] = 12'h444;
rom[85965] = 12'h444;
rom[85966] = 12'h444;
rom[85967] = 12'h444;
rom[85968] = 12'h444;
rom[85969] = 12'h444;
rom[85970] = 12'h444;
rom[85971] = 12'h444;
rom[85972] = 12'h444;
rom[85973] = 12'h444;
rom[85974] = 12'h444;
rom[85975] = 12'h444;
rom[85976] = 12'h333;
rom[85977] = 12'h333;
rom[85978] = 12'h333;
rom[85979] = 12'h333;
rom[85980] = 12'h333;
rom[85981] = 12'h333;
rom[85982] = 12'h333;
rom[85983] = 12'h333;
rom[85984] = 12'h222;
rom[85985] = 12'h222;
rom[85986] = 12'h222;
rom[85987] = 12'h222;
rom[85988] = 12'h222;
rom[85989] = 12'h222;
rom[85990] = 12'h222;
rom[85991] = 12'h222;
rom[85992] = 12'h222;
rom[85993] = 12'h222;
rom[85994] = 12'h222;
rom[85995] = 12'h222;
rom[85996] = 12'h222;
rom[85997] = 12'h222;
rom[85998] = 12'h222;
rom[85999] = 12'h222;
rom[86000] = 12'hfff;
rom[86001] = 12'hfff;
rom[86002] = 12'hfff;
rom[86003] = 12'hfff;
rom[86004] = 12'hfff;
rom[86005] = 12'hfff;
rom[86006] = 12'hfff;
rom[86007] = 12'hfff;
rom[86008] = 12'hfff;
rom[86009] = 12'hfff;
rom[86010] = 12'hfff;
rom[86011] = 12'hfff;
rom[86012] = 12'hfff;
rom[86013] = 12'hfff;
rom[86014] = 12'hfff;
rom[86015] = 12'hfff;
rom[86016] = 12'hfff;
rom[86017] = 12'hfff;
rom[86018] = 12'hfff;
rom[86019] = 12'hfff;
rom[86020] = 12'hfff;
rom[86021] = 12'hfff;
rom[86022] = 12'hfff;
rom[86023] = 12'hfff;
rom[86024] = 12'hfff;
rom[86025] = 12'hfff;
rom[86026] = 12'hfff;
rom[86027] = 12'hfff;
rom[86028] = 12'hfff;
rom[86029] = 12'hfff;
rom[86030] = 12'hfff;
rom[86031] = 12'hfff;
rom[86032] = 12'hfff;
rom[86033] = 12'hfff;
rom[86034] = 12'hfff;
rom[86035] = 12'hfff;
rom[86036] = 12'hfff;
rom[86037] = 12'hfff;
rom[86038] = 12'hfff;
rom[86039] = 12'hfff;
rom[86040] = 12'hfff;
rom[86041] = 12'hfff;
rom[86042] = 12'hfff;
rom[86043] = 12'hfff;
rom[86044] = 12'hfff;
rom[86045] = 12'hfff;
rom[86046] = 12'hfff;
rom[86047] = 12'hfff;
rom[86048] = 12'hfff;
rom[86049] = 12'hfff;
rom[86050] = 12'hfff;
rom[86051] = 12'hfff;
rom[86052] = 12'hfff;
rom[86053] = 12'hfff;
rom[86054] = 12'hfff;
rom[86055] = 12'hfff;
rom[86056] = 12'hfff;
rom[86057] = 12'hfff;
rom[86058] = 12'hfff;
rom[86059] = 12'hfff;
rom[86060] = 12'hfff;
rom[86061] = 12'hfff;
rom[86062] = 12'hfff;
rom[86063] = 12'hfff;
rom[86064] = 12'hfff;
rom[86065] = 12'hfff;
rom[86066] = 12'hfff;
rom[86067] = 12'hfff;
rom[86068] = 12'hfff;
rom[86069] = 12'hfff;
rom[86070] = 12'hfff;
rom[86071] = 12'hfff;
rom[86072] = 12'hfff;
rom[86073] = 12'hfff;
rom[86074] = 12'hfff;
rom[86075] = 12'hfff;
rom[86076] = 12'hfff;
rom[86077] = 12'hfff;
rom[86078] = 12'hfff;
rom[86079] = 12'hfff;
rom[86080] = 12'hfff;
rom[86081] = 12'hfff;
rom[86082] = 12'hfff;
rom[86083] = 12'hfff;
rom[86084] = 12'hfff;
rom[86085] = 12'hfff;
rom[86086] = 12'hfff;
rom[86087] = 12'hfff;
rom[86088] = 12'hfff;
rom[86089] = 12'hfff;
rom[86090] = 12'hfff;
rom[86091] = 12'hfff;
rom[86092] = 12'hfff;
rom[86093] = 12'hfff;
rom[86094] = 12'hfff;
rom[86095] = 12'hfff;
rom[86096] = 12'hfff;
rom[86097] = 12'hfff;
rom[86098] = 12'hfff;
rom[86099] = 12'hfff;
rom[86100] = 12'hfff;
rom[86101] = 12'hfff;
rom[86102] = 12'hfff;
rom[86103] = 12'hfff;
rom[86104] = 12'hfff;
rom[86105] = 12'hfff;
rom[86106] = 12'hfff;
rom[86107] = 12'hfff;
rom[86108] = 12'hfff;
rom[86109] = 12'hfff;
rom[86110] = 12'hfff;
rom[86111] = 12'hfff;
rom[86112] = 12'hfff;
rom[86113] = 12'hfff;
rom[86114] = 12'hfff;
rom[86115] = 12'hfff;
rom[86116] = 12'hfff;
rom[86117] = 12'hfff;
rom[86118] = 12'hfff;
rom[86119] = 12'hfff;
rom[86120] = 12'hfff;
rom[86121] = 12'hfff;
rom[86122] = 12'hfff;
rom[86123] = 12'hfff;
rom[86124] = 12'hfff;
rom[86125] = 12'heee;
rom[86126] = 12'heee;
rom[86127] = 12'heee;
rom[86128] = 12'hddd;
rom[86129] = 12'hddd;
rom[86130] = 12'hddd;
rom[86131] = 12'hddd;
rom[86132] = 12'hccc;
rom[86133] = 12'hccc;
rom[86134] = 12'hccc;
rom[86135] = 12'hccc;
rom[86136] = 12'hccc;
rom[86137] = 12'hbbb;
rom[86138] = 12'hbbb;
rom[86139] = 12'hbbb;
rom[86140] = 12'haaa;
rom[86141] = 12'haaa;
rom[86142] = 12'haaa;
rom[86143] = 12'haaa;
rom[86144] = 12'h999;
rom[86145] = 12'haaa;
rom[86146] = 12'haaa;
rom[86147] = 12'hbbb;
rom[86148] = 12'hbbb;
rom[86149] = 12'hbbb;
rom[86150] = 12'hbbb;
rom[86151] = 12'hccc;
rom[86152] = 12'hccc;
rom[86153] = 12'hbbb;
rom[86154] = 12'hbbb;
rom[86155] = 12'hbbb;
rom[86156] = 12'hbbb;
rom[86157] = 12'haaa;
rom[86158] = 12'haaa;
rom[86159] = 12'h999;
rom[86160] = 12'h888;
rom[86161] = 12'h888;
rom[86162] = 12'h777;
rom[86163] = 12'h777;
rom[86164] = 12'h777;
rom[86165] = 12'h666;
rom[86166] = 12'h666;
rom[86167] = 12'h666;
rom[86168] = 12'h666;
rom[86169] = 12'h555;
rom[86170] = 12'h555;
rom[86171] = 12'h555;
rom[86172] = 12'h555;
rom[86173] = 12'h555;
rom[86174] = 12'h555;
rom[86175] = 12'h555;
rom[86176] = 12'h555;
rom[86177] = 12'h555;
rom[86178] = 12'h555;
rom[86179] = 12'h555;
rom[86180] = 12'h555;
rom[86181] = 12'h555;
rom[86182] = 12'h555;
rom[86183] = 12'h555;
rom[86184] = 12'h555;
rom[86185] = 12'h555;
rom[86186] = 12'h555;
rom[86187] = 12'h555;
rom[86188] = 12'h555;
rom[86189] = 12'h555;
rom[86190] = 12'h555;
rom[86191] = 12'h555;
rom[86192] = 12'h555;
rom[86193] = 12'h444;
rom[86194] = 12'h444;
rom[86195] = 12'h444;
rom[86196] = 12'h444;
rom[86197] = 12'h444;
rom[86198] = 12'h444;
rom[86199] = 12'h444;
rom[86200] = 12'h444;
rom[86201] = 12'h555;
rom[86202] = 12'h555;
rom[86203] = 12'h666;
rom[86204] = 12'h666;
rom[86205] = 12'h555;
rom[86206] = 12'h555;
rom[86207] = 12'h555;
rom[86208] = 12'h555;
rom[86209] = 12'h555;
rom[86210] = 12'h555;
rom[86211] = 12'h444;
rom[86212] = 12'h555;
rom[86213] = 12'h666;
rom[86214] = 12'h777;
rom[86215] = 12'h666;
rom[86216] = 12'h888;
rom[86217] = 12'h777;
rom[86218] = 12'h666;
rom[86219] = 12'h555;
rom[86220] = 12'h444;
rom[86221] = 12'h444;
rom[86222] = 12'h333;
rom[86223] = 12'h333;
rom[86224] = 12'h222;
rom[86225] = 12'h222;
rom[86226] = 12'h222;
rom[86227] = 12'h222;
rom[86228] = 12'h222;
rom[86229] = 12'h222;
rom[86230] = 12'h111;
rom[86231] = 12'h111;
rom[86232] = 12'h111;
rom[86233] = 12'h111;
rom[86234] = 12'h111;
rom[86235] = 12'h  0;
rom[86236] = 12'h  0;
rom[86237] = 12'h  0;
rom[86238] = 12'h  0;
rom[86239] = 12'h  0;
rom[86240] = 12'h  0;
rom[86241] = 12'h  0;
rom[86242] = 12'h  0;
rom[86243] = 12'h  0;
rom[86244] = 12'h  0;
rom[86245] = 12'h  0;
rom[86246] = 12'h  0;
rom[86247] = 12'h  0;
rom[86248] = 12'h  0;
rom[86249] = 12'h  0;
rom[86250] = 12'h  0;
rom[86251] = 12'h  0;
rom[86252] = 12'h  0;
rom[86253] = 12'h  0;
rom[86254] = 12'h  0;
rom[86255] = 12'h  0;
rom[86256] = 12'h  0;
rom[86257] = 12'h  0;
rom[86258] = 12'h  0;
rom[86259] = 12'h  0;
rom[86260] = 12'h  0;
rom[86261] = 12'h111;
rom[86262] = 12'h111;
rom[86263] = 12'h111;
rom[86264] = 12'h111;
rom[86265] = 12'h111;
rom[86266] = 12'h111;
rom[86267] = 12'h111;
rom[86268] = 12'h111;
rom[86269] = 12'h222;
rom[86270] = 12'h222;
rom[86271] = 12'h222;
rom[86272] = 12'h222;
rom[86273] = 12'h222;
rom[86274] = 12'h333;
rom[86275] = 12'h333;
rom[86276] = 12'h333;
rom[86277] = 12'h333;
rom[86278] = 12'h444;
rom[86279] = 12'h444;
rom[86280] = 12'h666;
rom[86281] = 12'h888;
rom[86282] = 12'h999;
rom[86283] = 12'h999;
rom[86284] = 12'h888;
rom[86285] = 12'h777;
rom[86286] = 12'h777;
rom[86287] = 12'h777;
rom[86288] = 12'h666;
rom[86289] = 12'h666;
rom[86290] = 12'h666;
rom[86291] = 12'h666;
rom[86292] = 12'h666;
rom[86293] = 12'h666;
rom[86294] = 12'h666;
rom[86295] = 12'h666;
rom[86296] = 12'h666;
rom[86297] = 12'h777;
rom[86298] = 12'h777;
rom[86299] = 12'h777;
rom[86300] = 12'h777;
rom[86301] = 12'h777;
rom[86302] = 12'h888;
rom[86303] = 12'h999;
rom[86304] = 12'haaa;
rom[86305] = 12'hbbb;
rom[86306] = 12'hbbb;
rom[86307] = 12'haaa;
rom[86308] = 12'h999;
rom[86309] = 12'h888;
rom[86310] = 12'h888;
rom[86311] = 12'h888;
rom[86312] = 12'h777;
rom[86313] = 12'h777;
rom[86314] = 12'h888;
rom[86315] = 12'h999;
rom[86316] = 12'haaa;
rom[86317] = 12'haaa;
rom[86318] = 12'hbbb;
rom[86319] = 12'hccc;
rom[86320] = 12'hddd;
rom[86321] = 12'hddd;
rom[86322] = 12'heee;
rom[86323] = 12'heee;
rom[86324] = 12'hfff;
rom[86325] = 12'hfff;
rom[86326] = 12'hfff;
rom[86327] = 12'hfff;
rom[86328] = 12'hfff;
rom[86329] = 12'hfff;
rom[86330] = 12'heee;
rom[86331] = 12'heee;
rom[86332] = 12'heee;
rom[86333] = 12'hddd;
rom[86334] = 12'hccc;
rom[86335] = 12'hccc;
rom[86336] = 12'hbbb;
rom[86337] = 12'haaa;
rom[86338] = 12'haaa;
rom[86339] = 12'h999;
rom[86340] = 12'h999;
rom[86341] = 12'h888;
rom[86342] = 12'h777;
rom[86343] = 12'h777;
rom[86344] = 12'h666;
rom[86345] = 12'h666;
rom[86346] = 12'h666;
rom[86347] = 12'h666;
rom[86348] = 12'h555;
rom[86349] = 12'h555;
rom[86350] = 12'h555;
rom[86351] = 12'h555;
rom[86352] = 12'h555;
rom[86353] = 12'h555;
rom[86354] = 12'h555;
rom[86355] = 12'h555;
rom[86356] = 12'h555;
rom[86357] = 12'h555;
rom[86358] = 12'h555;
rom[86359] = 12'h555;
rom[86360] = 12'h555;
rom[86361] = 12'h555;
rom[86362] = 12'h555;
rom[86363] = 12'h555;
rom[86364] = 12'h555;
rom[86365] = 12'h444;
rom[86366] = 12'h444;
rom[86367] = 12'h555;
rom[86368] = 12'h444;
rom[86369] = 12'h444;
rom[86370] = 12'h444;
rom[86371] = 12'h444;
rom[86372] = 12'h444;
rom[86373] = 12'h444;
rom[86374] = 12'h444;
rom[86375] = 12'h444;
rom[86376] = 12'h333;
rom[86377] = 12'h333;
rom[86378] = 12'h333;
rom[86379] = 12'h333;
rom[86380] = 12'h333;
rom[86381] = 12'h333;
rom[86382] = 12'h333;
rom[86383] = 12'h333;
rom[86384] = 12'h222;
rom[86385] = 12'h222;
rom[86386] = 12'h222;
rom[86387] = 12'h222;
rom[86388] = 12'h222;
rom[86389] = 12'h222;
rom[86390] = 12'h222;
rom[86391] = 12'h222;
rom[86392] = 12'h222;
rom[86393] = 12'h222;
rom[86394] = 12'h222;
rom[86395] = 12'h222;
rom[86396] = 12'h222;
rom[86397] = 12'h222;
rom[86398] = 12'h222;
rom[86399] = 12'h222;
rom[86400] = 12'hfff;
rom[86401] = 12'hfff;
rom[86402] = 12'hfff;
rom[86403] = 12'hfff;
rom[86404] = 12'hfff;
rom[86405] = 12'hfff;
rom[86406] = 12'hfff;
rom[86407] = 12'hfff;
rom[86408] = 12'hfff;
rom[86409] = 12'hfff;
rom[86410] = 12'hfff;
rom[86411] = 12'hfff;
rom[86412] = 12'hfff;
rom[86413] = 12'hfff;
rom[86414] = 12'hfff;
rom[86415] = 12'hfff;
rom[86416] = 12'hfff;
rom[86417] = 12'hfff;
rom[86418] = 12'hfff;
rom[86419] = 12'hfff;
rom[86420] = 12'hfff;
rom[86421] = 12'hfff;
rom[86422] = 12'hfff;
rom[86423] = 12'hfff;
rom[86424] = 12'hfff;
rom[86425] = 12'hfff;
rom[86426] = 12'hfff;
rom[86427] = 12'hfff;
rom[86428] = 12'hfff;
rom[86429] = 12'hfff;
rom[86430] = 12'hfff;
rom[86431] = 12'hfff;
rom[86432] = 12'hfff;
rom[86433] = 12'hfff;
rom[86434] = 12'hfff;
rom[86435] = 12'hfff;
rom[86436] = 12'hfff;
rom[86437] = 12'hfff;
rom[86438] = 12'hfff;
rom[86439] = 12'hfff;
rom[86440] = 12'hfff;
rom[86441] = 12'hfff;
rom[86442] = 12'hfff;
rom[86443] = 12'hfff;
rom[86444] = 12'hfff;
rom[86445] = 12'hfff;
rom[86446] = 12'hfff;
rom[86447] = 12'hfff;
rom[86448] = 12'hfff;
rom[86449] = 12'hfff;
rom[86450] = 12'hfff;
rom[86451] = 12'hfff;
rom[86452] = 12'hfff;
rom[86453] = 12'hfff;
rom[86454] = 12'hfff;
rom[86455] = 12'hfff;
rom[86456] = 12'hfff;
rom[86457] = 12'hfff;
rom[86458] = 12'hfff;
rom[86459] = 12'hfff;
rom[86460] = 12'hfff;
rom[86461] = 12'hfff;
rom[86462] = 12'hfff;
rom[86463] = 12'hfff;
rom[86464] = 12'hfff;
rom[86465] = 12'hfff;
rom[86466] = 12'hfff;
rom[86467] = 12'hfff;
rom[86468] = 12'hfff;
rom[86469] = 12'hfff;
rom[86470] = 12'hfff;
rom[86471] = 12'hfff;
rom[86472] = 12'hfff;
rom[86473] = 12'hfff;
rom[86474] = 12'hfff;
rom[86475] = 12'hfff;
rom[86476] = 12'hfff;
rom[86477] = 12'hfff;
rom[86478] = 12'hfff;
rom[86479] = 12'hfff;
rom[86480] = 12'hfff;
rom[86481] = 12'hfff;
rom[86482] = 12'hfff;
rom[86483] = 12'hfff;
rom[86484] = 12'hfff;
rom[86485] = 12'hfff;
rom[86486] = 12'hfff;
rom[86487] = 12'hfff;
rom[86488] = 12'hfff;
rom[86489] = 12'hfff;
rom[86490] = 12'hfff;
rom[86491] = 12'hfff;
rom[86492] = 12'hfff;
rom[86493] = 12'hfff;
rom[86494] = 12'hfff;
rom[86495] = 12'hfff;
rom[86496] = 12'hfff;
rom[86497] = 12'hfff;
rom[86498] = 12'hfff;
rom[86499] = 12'hfff;
rom[86500] = 12'hfff;
rom[86501] = 12'hfff;
rom[86502] = 12'hfff;
rom[86503] = 12'hfff;
rom[86504] = 12'hfff;
rom[86505] = 12'hfff;
rom[86506] = 12'hfff;
rom[86507] = 12'hfff;
rom[86508] = 12'hfff;
rom[86509] = 12'hfff;
rom[86510] = 12'hfff;
rom[86511] = 12'hfff;
rom[86512] = 12'hfff;
rom[86513] = 12'hfff;
rom[86514] = 12'hfff;
rom[86515] = 12'hfff;
rom[86516] = 12'hfff;
rom[86517] = 12'hfff;
rom[86518] = 12'hfff;
rom[86519] = 12'hfff;
rom[86520] = 12'hfff;
rom[86521] = 12'hfff;
rom[86522] = 12'hfff;
rom[86523] = 12'hfff;
rom[86524] = 12'hfff;
rom[86525] = 12'hfff;
rom[86526] = 12'heee;
rom[86527] = 12'heee;
rom[86528] = 12'hddd;
rom[86529] = 12'hddd;
rom[86530] = 12'hddd;
rom[86531] = 12'hddd;
rom[86532] = 12'hccc;
rom[86533] = 12'hccc;
rom[86534] = 12'hccc;
rom[86535] = 12'hccc;
rom[86536] = 12'hbbb;
rom[86537] = 12'hbbb;
rom[86538] = 12'hbbb;
rom[86539] = 12'hbbb;
rom[86540] = 12'haaa;
rom[86541] = 12'haaa;
rom[86542] = 12'h999;
rom[86543] = 12'h999;
rom[86544] = 12'h999;
rom[86545] = 12'h999;
rom[86546] = 12'h999;
rom[86547] = 12'h999;
rom[86548] = 12'haaa;
rom[86549] = 12'haaa;
rom[86550] = 12'haaa;
rom[86551] = 12'hbbb;
rom[86552] = 12'hbbb;
rom[86553] = 12'hbbb;
rom[86554] = 12'hbbb;
rom[86555] = 12'hbbb;
rom[86556] = 12'hbbb;
rom[86557] = 12'hbbb;
rom[86558] = 12'haaa;
rom[86559] = 12'haaa;
rom[86560] = 12'haaa;
rom[86561] = 12'h999;
rom[86562] = 12'h999;
rom[86563] = 12'h888;
rom[86564] = 12'h888;
rom[86565] = 12'h777;
rom[86566] = 12'h777;
rom[86567] = 12'h777;
rom[86568] = 12'h666;
rom[86569] = 12'h666;
rom[86570] = 12'h666;
rom[86571] = 12'h666;
rom[86572] = 12'h666;
rom[86573] = 12'h666;
rom[86574] = 12'h666;
rom[86575] = 12'h666;
rom[86576] = 12'h666;
rom[86577] = 12'h666;
rom[86578] = 12'h666;
rom[86579] = 12'h666;
rom[86580] = 12'h666;
rom[86581] = 12'h666;
rom[86582] = 12'h666;
rom[86583] = 12'h666;
rom[86584] = 12'h666;
rom[86585] = 12'h666;
rom[86586] = 12'h666;
rom[86587] = 12'h666;
rom[86588] = 12'h666;
rom[86589] = 12'h666;
rom[86590] = 12'h555;
rom[86591] = 12'h555;
rom[86592] = 12'h555;
rom[86593] = 12'h555;
rom[86594] = 12'h444;
rom[86595] = 12'h444;
rom[86596] = 12'h444;
rom[86597] = 12'h444;
rom[86598] = 12'h444;
rom[86599] = 12'h444;
rom[86600] = 12'h555;
rom[86601] = 12'h555;
rom[86602] = 12'h666;
rom[86603] = 12'h666;
rom[86604] = 12'h666;
rom[86605] = 12'h666;
rom[86606] = 12'h555;
rom[86607] = 12'h555;
rom[86608] = 12'h555;
rom[86609] = 12'h555;
rom[86610] = 12'h444;
rom[86611] = 12'h444;
rom[86612] = 12'h444;
rom[86613] = 12'h555;
rom[86614] = 12'h555;
rom[86615] = 12'h666;
rom[86616] = 12'h777;
rom[86617] = 12'h777;
rom[86618] = 12'h777;
rom[86619] = 12'h777;
rom[86620] = 12'h666;
rom[86621] = 12'h444;
rom[86622] = 12'h333;
rom[86623] = 12'h333;
rom[86624] = 12'h333;
rom[86625] = 12'h222;
rom[86626] = 12'h222;
rom[86627] = 12'h222;
rom[86628] = 12'h222;
rom[86629] = 12'h222;
rom[86630] = 12'h222;
rom[86631] = 12'h222;
rom[86632] = 12'h111;
rom[86633] = 12'h111;
rom[86634] = 12'h111;
rom[86635] = 12'h  0;
rom[86636] = 12'h  0;
rom[86637] = 12'h  0;
rom[86638] = 12'h  0;
rom[86639] = 12'h  0;
rom[86640] = 12'h  0;
rom[86641] = 12'h  0;
rom[86642] = 12'h  0;
rom[86643] = 12'h  0;
rom[86644] = 12'h  0;
rom[86645] = 12'h  0;
rom[86646] = 12'h  0;
rom[86647] = 12'h  0;
rom[86648] = 12'h  0;
rom[86649] = 12'h  0;
rom[86650] = 12'h  0;
rom[86651] = 12'h  0;
rom[86652] = 12'h  0;
rom[86653] = 12'h  0;
rom[86654] = 12'h  0;
rom[86655] = 12'h  0;
rom[86656] = 12'h  0;
rom[86657] = 12'h  0;
rom[86658] = 12'h  0;
rom[86659] = 12'h  0;
rom[86660] = 12'h  0;
rom[86661] = 12'h  0;
rom[86662] = 12'h  0;
rom[86663] = 12'h  0;
rom[86664] = 12'h111;
rom[86665] = 12'h111;
rom[86666] = 12'h111;
rom[86667] = 12'h111;
rom[86668] = 12'h111;
rom[86669] = 12'h111;
rom[86670] = 12'h222;
rom[86671] = 12'h222;
rom[86672] = 12'h222;
rom[86673] = 12'h222;
rom[86674] = 12'h222;
rom[86675] = 12'h333;
rom[86676] = 12'h333;
rom[86677] = 12'h333;
rom[86678] = 12'h444;
rom[86679] = 12'h444;
rom[86680] = 12'h666;
rom[86681] = 12'h888;
rom[86682] = 12'h999;
rom[86683] = 12'h999;
rom[86684] = 12'h888;
rom[86685] = 12'h777;
rom[86686] = 12'h777;
rom[86687] = 12'h777;
rom[86688] = 12'h777;
rom[86689] = 12'h777;
rom[86690] = 12'h666;
rom[86691] = 12'h666;
rom[86692] = 12'h666;
rom[86693] = 12'h666;
rom[86694] = 12'h666;
rom[86695] = 12'h666;
rom[86696] = 12'h777;
rom[86697] = 12'h777;
rom[86698] = 12'h777;
rom[86699] = 12'h777;
rom[86700] = 12'h888;
rom[86701] = 12'h888;
rom[86702] = 12'h888;
rom[86703] = 12'h999;
rom[86704] = 12'hbbb;
rom[86705] = 12'hbbb;
rom[86706] = 12'hbbb;
rom[86707] = 12'haaa;
rom[86708] = 12'h999;
rom[86709] = 12'h999;
rom[86710] = 12'h999;
rom[86711] = 12'h999;
rom[86712] = 12'h888;
rom[86713] = 12'h888;
rom[86714] = 12'h888;
rom[86715] = 12'h888;
rom[86716] = 12'h888;
rom[86717] = 12'h999;
rom[86718] = 12'h999;
rom[86719] = 12'h999;
rom[86720] = 12'haaa;
rom[86721] = 12'haaa;
rom[86722] = 12'hbbb;
rom[86723] = 12'hbbb;
rom[86724] = 12'hccc;
rom[86725] = 12'hddd;
rom[86726] = 12'heee;
rom[86727] = 12'heee;
rom[86728] = 12'hfff;
rom[86729] = 12'hfff;
rom[86730] = 12'hfff;
rom[86731] = 12'hfff;
rom[86732] = 12'hfff;
rom[86733] = 12'hfff;
rom[86734] = 12'hfff;
rom[86735] = 12'hfff;
rom[86736] = 12'hfff;
rom[86737] = 12'hfff;
rom[86738] = 12'heee;
rom[86739] = 12'heee;
rom[86740] = 12'hddd;
rom[86741] = 12'hddd;
rom[86742] = 12'hccc;
rom[86743] = 12'hccc;
rom[86744] = 12'hbbb;
rom[86745] = 12'hbbb;
rom[86746] = 12'haaa;
rom[86747] = 12'haaa;
rom[86748] = 12'haaa;
rom[86749] = 12'h999;
rom[86750] = 12'h888;
rom[86751] = 12'h888;
rom[86752] = 12'h777;
rom[86753] = 12'h777;
rom[86754] = 12'h777;
rom[86755] = 12'h777;
rom[86756] = 12'h777;
rom[86757] = 12'h666;
rom[86758] = 12'h666;
rom[86759] = 12'h555;
rom[86760] = 12'h555;
rom[86761] = 12'h555;
rom[86762] = 12'h555;
rom[86763] = 12'h555;
rom[86764] = 12'h555;
rom[86765] = 12'h555;
rom[86766] = 12'h555;
rom[86767] = 12'h555;
rom[86768] = 12'h555;
rom[86769] = 12'h555;
rom[86770] = 12'h555;
rom[86771] = 12'h555;
rom[86772] = 12'h555;
rom[86773] = 12'h555;
rom[86774] = 12'h444;
rom[86775] = 12'h444;
rom[86776] = 12'h444;
rom[86777] = 12'h444;
rom[86778] = 12'h444;
rom[86779] = 12'h444;
rom[86780] = 12'h444;
rom[86781] = 12'h333;
rom[86782] = 12'h333;
rom[86783] = 12'h333;
rom[86784] = 12'h333;
rom[86785] = 12'h333;
rom[86786] = 12'h333;
rom[86787] = 12'h333;
rom[86788] = 12'h333;
rom[86789] = 12'h333;
rom[86790] = 12'h222;
rom[86791] = 12'h222;
rom[86792] = 12'h222;
rom[86793] = 12'h222;
rom[86794] = 12'h222;
rom[86795] = 12'h222;
rom[86796] = 12'h222;
rom[86797] = 12'h222;
rom[86798] = 12'h222;
rom[86799] = 12'h222;
rom[86800] = 12'hfff;
rom[86801] = 12'hfff;
rom[86802] = 12'hfff;
rom[86803] = 12'hfff;
rom[86804] = 12'hfff;
rom[86805] = 12'hfff;
rom[86806] = 12'hfff;
rom[86807] = 12'hfff;
rom[86808] = 12'hfff;
rom[86809] = 12'hfff;
rom[86810] = 12'hfff;
rom[86811] = 12'hfff;
rom[86812] = 12'hfff;
rom[86813] = 12'hfff;
rom[86814] = 12'hfff;
rom[86815] = 12'hfff;
rom[86816] = 12'hfff;
rom[86817] = 12'hfff;
rom[86818] = 12'hfff;
rom[86819] = 12'hfff;
rom[86820] = 12'hfff;
rom[86821] = 12'hfff;
rom[86822] = 12'hfff;
rom[86823] = 12'hfff;
rom[86824] = 12'hfff;
rom[86825] = 12'hfff;
rom[86826] = 12'hfff;
rom[86827] = 12'hfff;
rom[86828] = 12'hfff;
rom[86829] = 12'hfff;
rom[86830] = 12'hfff;
rom[86831] = 12'hfff;
rom[86832] = 12'hfff;
rom[86833] = 12'hfff;
rom[86834] = 12'hfff;
rom[86835] = 12'hfff;
rom[86836] = 12'hfff;
rom[86837] = 12'hfff;
rom[86838] = 12'hfff;
rom[86839] = 12'hfff;
rom[86840] = 12'hfff;
rom[86841] = 12'hfff;
rom[86842] = 12'hfff;
rom[86843] = 12'hfff;
rom[86844] = 12'hfff;
rom[86845] = 12'hfff;
rom[86846] = 12'hfff;
rom[86847] = 12'hfff;
rom[86848] = 12'hfff;
rom[86849] = 12'hfff;
rom[86850] = 12'hfff;
rom[86851] = 12'hfff;
rom[86852] = 12'hfff;
rom[86853] = 12'hfff;
rom[86854] = 12'hfff;
rom[86855] = 12'hfff;
rom[86856] = 12'hfff;
rom[86857] = 12'hfff;
rom[86858] = 12'hfff;
rom[86859] = 12'hfff;
rom[86860] = 12'hfff;
rom[86861] = 12'hfff;
rom[86862] = 12'hfff;
rom[86863] = 12'hfff;
rom[86864] = 12'hfff;
rom[86865] = 12'hfff;
rom[86866] = 12'hfff;
rom[86867] = 12'hfff;
rom[86868] = 12'hfff;
rom[86869] = 12'hfff;
rom[86870] = 12'hfff;
rom[86871] = 12'hfff;
rom[86872] = 12'hfff;
rom[86873] = 12'hfff;
rom[86874] = 12'hfff;
rom[86875] = 12'hfff;
rom[86876] = 12'hfff;
rom[86877] = 12'hfff;
rom[86878] = 12'hfff;
rom[86879] = 12'hfff;
rom[86880] = 12'hfff;
rom[86881] = 12'hfff;
rom[86882] = 12'hfff;
rom[86883] = 12'hfff;
rom[86884] = 12'hfff;
rom[86885] = 12'hfff;
rom[86886] = 12'hfff;
rom[86887] = 12'hfff;
rom[86888] = 12'hfff;
rom[86889] = 12'hfff;
rom[86890] = 12'hfff;
rom[86891] = 12'hfff;
rom[86892] = 12'hfff;
rom[86893] = 12'hfff;
rom[86894] = 12'hfff;
rom[86895] = 12'hfff;
rom[86896] = 12'hfff;
rom[86897] = 12'hfff;
rom[86898] = 12'hfff;
rom[86899] = 12'hfff;
rom[86900] = 12'hfff;
rom[86901] = 12'hfff;
rom[86902] = 12'hfff;
rom[86903] = 12'hfff;
rom[86904] = 12'hfff;
rom[86905] = 12'hfff;
rom[86906] = 12'hfff;
rom[86907] = 12'hfff;
rom[86908] = 12'hfff;
rom[86909] = 12'hfff;
rom[86910] = 12'hfff;
rom[86911] = 12'hfff;
rom[86912] = 12'hfff;
rom[86913] = 12'hfff;
rom[86914] = 12'hfff;
rom[86915] = 12'hfff;
rom[86916] = 12'hfff;
rom[86917] = 12'hfff;
rom[86918] = 12'hfff;
rom[86919] = 12'hfff;
rom[86920] = 12'hfff;
rom[86921] = 12'hfff;
rom[86922] = 12'hfff;
rom[86923] = 12'hfff;
rom[86924] = 12'hfff;
rom[86925] = 12'hfff;
rom[86926] = 12'heee;
rom[86927] = 12'heee;
rom[86928] = 12'heee;
rom[86929] = 12'hddd;
rom[86930] = 12'hddd;
rom[86931] = 12'hddd;
rom[86932] = 12'hccc;
rom[86933] = 12'hccc;
rom[86934] = 12'hccc;
rom[86935] = 12'hccc;
rom[86936] = 12'hccc;
rom[86937] = 12'hbbb;
rom[86938] = 12'hbbb;
rom[86939] = 12'hbbb;
rom[86940] = 12'haaa;
rom[86941] = 12'haaa;
rom[86942] = 12'haaa;
rom[86943] = 12'h999;
rom[86944] = 12'h999;
rom[86945] = 12'h999;
rom[86946] = 12'h999;
rom[86947] = 12'h999;
rom[86948] = 12'h999;
rom[86949] = 12'h999;
rom[86950] = 12'h999;
rom[86951] = 12'h999;
rom[86952] = 12'haaa;
rom[86953] = 12'haaa;
rom[86954] = 12'haaa;
rom[86955] = 12'haaa;
rom[86956] = 12'haaa;
rom[86957] = 12'haaa;
rom[86958] = 12'haaa;
rom[86959] = 12'haaa;
rom[86960] = 12'haaa;
rom[86961] = 12'haaa;
rom[86962] = 12'h999;
rom[86963] = 12'h999;
rom[86964] = 12'h888;
rom[86965] = 12'h888;
rom[86966] = 12'h888;
rom[86967] = 12'h777;
rom[86968] = 12'h777;
rom[86969] = 12'h777;
rom[86970] = 12'h777;
rom[86971] = 12'h777;
rom[86972] = 12'h777;
rom[86973] = 12'h777;
rom[86974] = 12'h777;
rom[86975] = 12'h666;
rom[86976] = 12'h666;
rom[86977] = 12'h666;
rom[86978] = 12'h666;
rom[86979] = 12'h666;
rom[86980] = 12'h666;
rom[86981] = 12'h666;
rom[86982] = 12'h666;
rom[86983] = 12'h666;
rom[86984] = 12'h555;
rom[86985] = 12'h555;
rom[86986] = 12'h666;
rom[86987] = 12'h666;
rom[86988] = 12'h666;
rom[86989] = 12'h555;
rom[86990] = 12'h555;
rom[86991] = 12'h555;
rom[86992] = 12'h555;
rom[86993] = 12'h555;
rom[86994] = 12'h555;
rom[86995] = 12'h555;
rom[86996] = 12'h555;
rom[86997] = 12'h555;
rom[86998] = 12'h555;
rom[86999] = 12'h555;
rom[87000] = 12'h555;
rom[87001] = 12'h555;
rom[87002] = 12'h666;
rom[87003] = 12'h666;
rom[87004] = 12'h666;
rom[87005] = 12'h555;
rom[87006] = 12'h555;
rom[87007] = 12'h555;
rom[87008] = 12'h555;
rom[87009] = 12'h555;
rom[87010] = 12'h444;
rom[87011] = 12'h444;
rom[87012] = 12'h444;
rom[87013] = 12'h444;
rom[87014] = 12'h555;
rom[87015] = 12'h555;
rom[87016] = 12'h666;
rom[87017] = 12'h777;
rom[87018] = 12'h777;
rom[87019] = 12'h777;
rom[87020] = 12'h666;
rom[87021] = 12'h555;
rom[87022] = 12'h444;
rom[87023] = 12'h444;
rom[87024] = 12'h333;
rom[87025] = 12'h222;
rom[87026] = 12'h222;
rom[87027] = 12'h222;
rom[87028] = 12'h222;
rom[87029] = 12'h222;
rom[87030] = 12'h222;
rom[87031] = 12'h222;
rom[87032] = 12'h111;
rom[87033] = 12'h111;
rom[87034] = 12'h111;
rom[87035] = 12'h  0;
rom[87036] = 12'h  0;
rom[87037] = 12'h  0;
rom[87038] = 12'h  0;
rom[87039] = 12'h  0;
rom[87040] = 12'h  0;
rom[87041] = 12'h  0;
rom[87042] = 12'h  0;
rom[87043] = 12'h  0;
rom[87044] = 12'h  0;
rom[87045] = 12'h  0;
rom[87046] = 12'h  0;
rom[87047] = 12'h  0;
rom[87048] = 12'h  0;
rom[87049] = 12'h  0;
rom[87050] = 12'h  0;
rom[87051] = 12'h  0;
rom[87052] = 12'h  0;
rom[87053] = 12'h  0;
rom[87054] = 12'h  0;
rom[87055] = 12'h  0;
rom[87056] = 12'h  0;
rom[87057] = 12'h  0;
rom[87058] = 12'h  0;
rom[87059] = 12'h  0;
rom[87060] = 12'h  0;
rom[87061] = 12'h  0;
rom[87062] = 12'h  0;
rom[87063] = 12'h  0;
rom[87064] = 12'h  0;
rom[87065] = 12'h  0;
rom[87066] = 12'h  0;
rom[87067] = 12'h111;
rom[87068] = 12'h111;
rom[87069] = 12'h111;
rom[87070] = 12'h111;
rom[87071] = 12'h111;
rom[87072] = 12'h222;
rom[87073] = 12'h222;
rom[87074] = 12'h222;
rom[87075] = 12'h333;
rom[87076] = 12'h333;
rom[87077] = 12'h333;
rom[87078] = 12'h444;
rom[87079] = 12'h444;
rom[87080] = 12'h666;
rom[87081] = 12'h888;
rom[87082] = 12'h999;
rom[87083] = 12'h999;
rom[87084] = 12'h888;
rom[87085] = 12'h777;
rom[87086] = 12'h777;
rom[87087] = 12'h777;
rom[87088] = 12'h777;
rom[87089] = 12'h777;
rom[87090] = 12'h777;
rom[87091] = 12'h666;
rom[87092] = 12'h666;
rom[87093] = 12'h666;
rom[87094] = 12'h666;
rom[87095] = 12'h666;
rom[87096] = 12'h666;
rom[87097] = 12'h666;
rom[87098] = 12'h777;
rom[87099] = 12'h777;
rom[87100] = 12'h777;
rom[87101] = 12'h888;
rom[87102] = 12'h999;
rom[87103] = 12'haaa;
rom[87104] = 12'hbbb;
rom[87105] = 12'hbbb;
rom[87106] = 12'hbbb;
rom[87107] = 12'haaa;
rom[87108] = 12'h999;
rom[87109] = 12'h999;
rom[87110] = 12'h999;
rom[87111] = 12'h999;
rom[87112] = 12'haaa;
rom[87113] = 12'haaa;
rom[87114] = 12'haaa;
rom[87115] = 12'haaa;
rom[87116] = 12'haaa;
rom[87117] = 12'haaa;
rom[87118] = 12'haaa;
rom[87119] = 12'haaa;
rom[87120] = 12'haaa;
rom[87121] = 12'haaa;
rom[87122] = 12'haaa;
rom[87123] = 12'haaa;
rom[87124] = 12'haaa;
rom[87125] = 12'haaa;
rom[87126] = 12'hbbb;
rom[87127] = 12'hbbb;
rom[87128] = 12'hccc;
rom[87129] = 12'hddd;
rom[87130] = 12'hddd;
rom[87131] = 12'heee;
rom[87132] = 12'heee;
rom[87133] = 12'hfff;
rom[87134] = 12'hfff;
rom[87135] = 12'hfff;
rom[87136] = 12'hfff;
rom[87137] = 12'hfff;
rom[87138] = 12'hfff;
rom[87139] = 12'heee;
rom[87140] = 12'heee;
rom[87141] = 12'hddd;
rom[87142] = 12'hddd;
rom[87143] = 12'hddd;
rom[87144] = 12'hccc;
rom[87145] = 12'hccc;
rom[87146] = 12'hccc;
rom[87147] = 12'hccc;
rom[87148] = 12'hccc;
rom[87149] = 12'hccc;
rom[87150] = 12'hbbb;
rom[87151] = 12'hbbb;
rom[87152] = 12'hbbb;
rom[87153] = 12'hbbb;
rom[87154] = 12'haaa;
rom[87155] = 12'haaa;
rom[87156] = 12'haaa;
rom[87157] = 12'haaa;
rom[87158] = 12'h999;
rom[87159] = 12'h888;
rom[87160] = 12'h888;
rom[87161] = 12'h888;
rom[87162] = 12'h888;
rom[87163] = 12'h777;
rom[87164] = 12'h777;
rom[87165] = 12'h666;
rom[87166] = 12'h666;
rom[87167] = 12'h666;
rom[87168] = 12'h555;
rom[87169] = 12'h555;
rom[87170] = 12'h555;
rom[87171] = 12'h555;
rom[87172] = 12'h555;
rom[87173] = 12'h555;
rom[87174] = 12'h555;
rom[87175] = 12'h555;
rom[87176] = 12'h555;
rom[87177] = 12'h444;
rom[87178] = 12'h444;
rom[87179] = 12'h444;
rom[87180] = 12'h444;
rom[87181] = 12'h444;
rom[87182] = 12'h333;
rom[87183] = 12'h333;
rom[87184] = 12'h333;
rom[87185] = 12'h333;
rom[87186] = 12'h333;
rom[87187] = 12'h333;
rom[87188] = 12'h333;
rom[87189] = 12'h333;
rom[87190] = 12'h333;
rom[87191] = 12'h222;
rom[87192] = 12'h222;
rom[87193] = 12'h222;
rom[87194] = 12'h222;
rom[87195] = 12'h222;
rom[87196] = 12'h222;
rom[87197] = 12'h222;
rom[87198] = 12'h222;
rom[87199] = 12'h222;
rom[87200] = 12'hfff;
rom[87201] = 12'hfff;
rom[87202] = 12'hfff;
rom[87203] = 12'hfff;
rom[87204] = 12'hfff;
rom[87205] = 12'hfff;
rom[87206] = 12'hfff;
rom[87207] = 12'hfff;
rom[87208] = 12'hfff;
rom[87209] = 12'hfff;
rom[87210] = 12'hfff;
rom[87211] = 12'hfff;
rom[87212] = 12'hfff;
rom[87213] = 12'hfff;
rom[87214] = 12'hfff;
rom[87215] = 12'hfff;
rom[87216] = 12'hfff;
rom[87217] = 12'hfff;
rom[87218] = 12'hfff;
rom[87219] = 12'hfff;
rom[87220] = 12'hfff;
rom[87221] = 12'hfff;
rom[87222] = 12'hfff;
rom[87223] = 12'hfff;
rom[87224] = 12'hfff;
rom[87225] = 12'hfff;
rom[87226] = 12'hfff;
rom[87227] = 12'hfff;
rom[87228] = 12'hfff;
rom[87229] = 12'hfff;
rom[87230] = 12'hfff;
rom[87231] = 12'hfff;
rom[87232] = 12'hfff;
rom[87233] = 12'hfff;
rom[87234] = 12'hfff;
rom[87235] = 12'hfff;
rom[87236] = 12'hfff;
rom[87237] = 12'hfff;
rom[87238] = 12'hfff;
rom[87239] = 12'hfff;
rom[87240] = 12'hfff;
rom[87241] = 12'hfff;
rom[87242] = 12'hfff;
rom[87243] = 12'hfff;
rom[87244] = 12'hfff;
rom[87245] = 12'hfff;
rom[87246] = 12'hfff;
rom[87247] = 12'hfff;
rom[87248] = 12'hfff;
rom[87249] = 12'hfff;
rom[87250] = 12'hfff;
rom[87251] = 12'hfff;
rom[87252] = 12'hfff;
rom[87253] = 12'hfff;
rom[87254] = 12'hfff;
rom[87255] = 12'hfff;
rom[87256] = 12'hfff;
rom[87257] = 12'hfff;
rom[87258] = 12'hfff;
rom[87259] = 12'hfff;
rom[87260] = 12'hfff;
rom[87261] = 12'hfff;
rom[87262] = 12'hfff;
rom[87263] = 12'hfff;
rom[87264] = 12'hfff;
rom[87265] = 12'hfff;
rom[87266] = 12'hfff;
rom[87267] = 12'hfff;
rom[87268] = 12'hfff;
rom[87269] = 12'hfff;
rom[87270] = 12'hfff;
rom[87271] = 12'hfff;
rom[87272] = 12'hfff;
rom[87273] = 12'hfff;
rom[87274] = 12'hfff;
rom[87275] = 12'hfff;
rom[87276] = 12'hfff;
rom[87277] = 12'hfff;
rom[87278] = 12'hfff;
rom[87279] = 12'hfff;
rom[87280] = 12'hfff;
rom[87281] = 12'hfff;
rom[87282] = 12'hfff;
rom[87283] = 12'hfff;
rom[87284] = 12'hfff;
rom[87285] = 12'hfff;
rom[87286] = 12'hfff;
rom[87287] = 12'hfff;
rom[87288] = 12'hfff;
rom[87289] = 12'hfff;
rom[87290] = 12'hfff;
rom[87291] = 12'hfff;
rom[87292] = 12'hfff;
rom[87293] = 12'hfff;
rom[87294] = 12'hfff;
rom[87295] = 12'hfff;
rom[87296] = 12'hfff;
rom[87297] = 12'hfff;
rom[87298] = 12'hfff;
rom[87299] = 12'hfff;
rom[87300] = 12'hfff;
rom[87301] = 12'hfff;
rom[87302] = 12'hfff;
rom[87303] = 12'hfff;
rom[87304] = 12'hfff;
rom[87305] = 12'hfff;
rom[87306] = 12'hfff;
rom[87307] = 12'hfff;
rom[87308] = 12'hfff;
rom[87309] = 12'hfff;
rom[87310] = 12'hfff;
rom[87311] = 12'hfff;
rom[87312] = 12'hfff;
rom[87313] = 12'hfff;
rom[87314] = 12'hfff;
rom[87315] = 12'hfff;
rom[87316] = 12'hfff;
rom[87317] = 12'hfff;
rom[87318] = 12'hfff;
rom[87319] = 12'hfff;
rom[87320] = 12'hfff;
rom[87321] = 12'hfff;
rom[87322] = 12'hfff;
rom[87323] = 12'hfff;
rom[87324] = 12'hfff;
rom[87325] = 12'hfff;
rom[87326] = 12'heee;
rom[87327] = 12'heee;
rom[87328] = 12'heee;
rom[87329] = 12'hddd;
rom[87330] = 12'hddd;
rom[87331] = 12'hddd;
rom[87332] = 12'hccc;
rom[87333] = 12'hccc;
rom[87334] = 12'hccc;
rom[87335] = 12'hccc;
rom[87336] = 12'hccc;
rom[87337] = 12'hbbb;
rom[87338] = 12'hbbb;
rom[87339] = 12'hbbb;
rom[87340] = 12'hbbb;
rom[87341] = 12'haaa;
rom[87342] = 12'haaa;
rom[87343] = 12'haaa;
rom[87344] = 12'haaa;
rom[87345] = 12'h999;
rom[87346] = 12'h999;
rom[87347] = 12'h999;
rom[87348] = 12'h888;
rom[87349] = 12'h888;
rom[87350] = 12'h888;
rom[87351] = 12'h888;
rom[87352] = 12'h888;
rom[87353] = 12'h888;
rom[87354] = 12'h999;
rom[87355] = 12'h999;
rom[87356] = 12'h999;
rom[87357] = 12'h999;
rom[87358] = 12'haaa;
rom[87359] = 12'haaa;
rom[87360] = 12'haaa;
rom[87361] = 12'haaa;
rom[87362] = 12'haaa;
rom[87363] = 12'h999;
rom[87364] = 12'h999;
rom[87365] = 12'h999;
rom[87366] = 12'h888;
rom[87367] = 12'h888;
rom[87368] = 12'h888;
rom[87369] = 12'h777;
rom[87370] = 12'h777;
rom[87371] = 12'h777;
rom[87372] = 12'h777;
rom[87373] = 12'h777;
rom[87374] = 12'h777;
rom[87375] = 12'h777;
rom[87376] = 12'h666;
rom[87377] = 12'h666;
rom[87378] = 12'h666;
rom[87379] = 12'h666;
rom[87380] = 12'h666;
rom[87381] = 12'h666;
rom[87382] = 12'h666;
rom[87383] = 12'h666;
rom[87384] = 12'h555;
rom[87385] = 12'h555;
rom[87386] = 12'h555;
rom[87387] = 12'h555;
rom[87388] = 12'h666;
rom[87389] = 12'h555;
rom[87390] = 12'h555;
rom[87391] = 12'h555;
rom[87392] = 12'h555;
rom[87393] = 12'h555;
rom[87394] = 12'h555;
rom[87395] = 12'h555;
rom[87396] = 12'h555;
rom[87397] = 12'h555;
rom[87398] = 12'h555;
rom[87399] = 12'h555;
rom[87400] = 12'h555;
rom[87401] = 12'h555;
rom[87402] = 12'h666;
rom[87403] = 12'h666;
rom[87404] = 12'h555;
rom[87405] = 12'h555;
rom[87406] = 12'h555;
rom[87407] = 12'h555;
rom[87408] = 12'h555;
rom[87409] = 12'h555;
rom[87410] = 12'h444;
rom[87411] = 12'h444;
rom[87412] = 12'h444;
rom[87413] = 12'h444;
rom[87414] = 12'h555;
rom[87415] = 12'h555;
rom[87416] = 12'h555;
rom[87417] = 12'h666;
rom[87418] = 12'h777;
rom[87419] = 12'h777;
rom[87420] = 12'h777;
rom[87421] = 12'h666;
rom[87422] = 12'h555;
rom[87423] = 12'h555;
rom[87424] = 12'h333;
rom[87425] = 12'h333;
rom[87426] = 12'h222;
rom[87427] = 12'h222;
rom[87428] = 12'h222;
rom[87429] = 12'h333;
rom[87430] = 12'h222;
rom[87431] = 12'h222;
rom[87432] = 12'h111;
rom[87433] = 12'h111;
rom[87434] = 12'h111;
rom[87435] = 12'h111;
rom[87436] = 12'h  0;
rom[87437] = 12'h  0;
rom[87438] = 12'h  0;
rom[87439] = 12'h  0;
rom[87440] = 12'h  0;
rom[87441] = 12'h  0;
rom[87442] = 12'h  0;
rom[87443] = 12'h  0;
rom[87444] = 12'h  0;
rom[87445] = 12'h  0;
rom[87446] = 12'h  0;
rom[87447] = 12'h  0;
rom[87448] = 12'h  0;
rom[87449] = 12'h  0;
rom[87450] = 12'h  0;
rom[87451] = 12'h  0;
rom[87452] = 12'h  0;
rom[87453] = 12'h  0;
rom[87454] = 12'h  0;
rom[87455] = 12'h  0;
rom[87456] = 12'h  0;
rom[87457] = 12'h  0;
rom[87458] = 12'h  0;
rom[87459] = 12'h  0;
rom[87460] = 12'h  0;
rom[87461] = 12'h  0;
rom[87462] = 12'h  0;
rom[87463] = 12'h  0;
rom[87464] = 12'h  0;
rom[87465] = 12'h  0;
rom[87466] = 12'h  0;
rom[87467] = 12'h  0;
rom[87468] = 12'h  0;
rom[87469] = 12'h111;
rom[87470] = 12'h111;
rom[87471] = 12'h111;
rom[87472] = 12'h222;
rom[87473] = 12'h222;
rom[87474] = 12'h222;
rom[87475] = 12'h222;
rom[87476] = 12'h333;
rom[87477] = 12'h333;
rom[87478] = 12'h444;
rom[87479] = 12'h444;
rom[87480] = 12'h666;
rom[87481] = 12'h888;
rom[87482] = 12'h999;
rom[87483] = 12'h999;
rom[87484] = 12'h888;
rom[87485] = 12'h777;
rom[87486] = 12'h777;
rom[87487] = 12'h777;
rom[87488] = 12'h777;
rom[87489] = 12'h777;
rom[87490] = 12'h777;
rom[87491] = 12'h777;
rom[87492] = 12'h777;
rom[87493] = 12'h777;
rom[87494] = 12'h777;
rom[87495] = 12'h666;
rom[87496] = 12'h777;
rom[87497] = 12'h777;
rom[87498] = 12'h777;
rom[87499] = 12'h777;
rom[87500] = 12'h777;
rom[87501] = 12'h888;
rom[87502] = 12'h999;
rom[87503] = 12'haaa;
rom[87504] = 12'hbbb;
rom[87505] = 12'hbbb;
rom[87506] = 12'haaa;
rom[87507] = 12'h999;
rom[87508] = 12'h999;
rom[87509] = 12'h999;
rom[87510] = 12'haaa;
rom[87511] = 12'haaa;
rom[87512] = 12'haaa;
rom[87513] = 12'haaa;
rom[87514] = 12'hbbb;
rom[87515] = 12'hbbb;
rom[87516] = 12'hccc;
rom[87517] = 12'hccc;
rom[87518] = 12'hbbb;
rom[87519] = 12'hbbb;
rom[87520] = 12'hbbb;
rom[87521] = 12'hbbb;
rom[87522] = 12'hbbb;
rom[87523] = 12'hbbb;
rom[87524] = 12'haaa;
rom[87525] = 12'haaa;
rom[87526] = 12'haaa;
rom[87527] = 12'haaa;
rom[87528] = 12'hbbb;
rom[87529] = 12'hbbb;
rom[87530] = 12'hbbb;
rom[87531] = 12'hccc;
rom[87532] = 12'hccc;
rom[87533] = 12'hddd;
rom[87534] = 12'hddd;
rom[87535] = 12'heee;
rom[87536] = 12'hfff;
rom[87537] = 12'hfff;
rom[87538] = 12'hfff;
rom[87539] = 12'hfff;
rom[87540] = 12'hfff;
rom[87541] = 12'heee;
rom[87542] = 12'heee;
rom[87543] = 12'hddd;
rom[87544] = 12'hccc;
rom[87545] = 12'hccc;
rom[87546] = 12'hccc;
rom[87547] = 12'hccc;
rom[87548] = 12'hccc;
rom[87549] = 12'hccc;
rom[87550] = 12'hccc;
rom[87551] = 12'hccc;
rom[87552] = 12'hccc;
rom[87553] = 12'hccc;
rom[87554] = 12'hccc;
rom[87555] = 12'hccc;
rom[87556] = 12'hccc;
rom[87557] = 12'hccc;
rom[87558] = 12'hbbb;
rom[87559] = 12'hbbb;
rom[87560] = 12'hbbb;
rom[87561] = 12'hbbb;
rom[87562] = 12'hbbb;
rom[87563] = 12'haaa;
rom[87564] = 12'haaa;
rom[87565] = 12'h999;
rom[87566] = 12'h999;
rom[87567] = 12'h999;
rom[87568] = 12'h888;
rom[87569] = 12'h888;
rom[87570] = 12'h777;
rom[87571] = 12'h777;
rom[87572] = 12'h666;
rom[87573] = 12'h666;
rom[87574] = 12'h666;
rom[87575] = 12'h666;
rom[87576] = 12'h555;
rom[87577] = 12'h555;
rom[87578] = 12'h555;
rom[87579] = 12'h555;
rom[87580] = 12'h444;
rom[87581] = 12'h444;
rom[87582] = 12'h444;
rom[87583] = 12'h444;
rom[87584] = 12'h444;
rom[87585] = 12'h333;
rom[87586] = 12'h333;
rom[87587] = 12'h333;
rom[87588] = 12'h333;
rom[87589] = 12'h333;
rom[87590] = 12'h333;
rom[87591] = 12'h333;
rom[87592] = 12'h222;
rom[87593] = 12'h222;
rom[87594] = 12'h222;
rom[87595] = 12'h222;
rom[87596] = 12'h222;
rom[87597] = 12'h222;
rom[87598] = 12'h222;
rom[87599] = 12'h111;
rom[87600] = 12'hfff;
rom[87601] = 12'hfff;
rom[87602] = 12'hfff;
rom[87603] = 12'hfff;
rom[87604] = 12'hfff;
rom[87605] = 12'hfff;
rom[87606] = 12'hfff;
rom[87607] = 12'hfff;
rom[87608] = 12'hfff;
rom[87609] = 12'hfff;
rom[87610] = 12'hfff;
rom[87611] = 12'hfff;
rom[87612] = 12'hfff;
rom[87613] = 12'hfff;
rom[87614] = 12'hfff;
rom[87615] = 12'hfff;
rom[87616] = 12'hfff;
rom[87617] = 12'hfff;
rom[87618] = 12'hfff;
rom[87619] = 12'hfff;
rom[87620] = 12'hfff;
rom[87621] = 12'hfff;
rom[87622] = 12'hfff;
rom[87623] = 12'hfff;
rom[87624] = 12'hfff;
rom[87625] = 12'hfff;
rom[87626] = 12'hfff;
rom[87627] = 12'hfff;
rom[87628] = 12'hfff;
rom[87629] = 12'hfff;
rom[87630] = 12'hfff;
rom[87631] = 12'hfff;
rom[87632] = 12'hfff;
rom[87633] = 12'hfff;
rom[87634] = 12'hfff;
rom[87635] = 12'hfff;
rom[87636] = 12'hfff;
rom[87637] = 12'hfff;
rom[87638] = 12'hfff;
rom[87639] = 12'hfff;
rom[87640] = 12'hfff;
rom[87641] = 12'hfff;
rom[87642] = 12'hfff;
rom[87643] = 12'hfff;
rom[87644] = 12'hfff;
rom[87645] = 12'hfff;
rom[87646] = 12'hfff;
rom[87647] = 12'hfff;
rom[87648] = 12'hfff;
rom[87649] = 12'hfff;
rom[87650] = 12'hfff;
rom[87651] = 12'hfff;
rom[87652] = 12'hfff;
rom[87653] = 12'hfff;
rom[87654] = 12'hfff;
rom[87655] = 12'hfff;
rom[87656] = 12'hfff;
rom[87657] = 12'hfff;
rom[87658] = 12'hfff;
rom[87659] = 12'hfff;
rom[87660] = 12'hfff;
rom[87661] = 12'hfff;
rom[87662] = 12'hfff;
rom[87663] = 12'hfff;
rom[87664] = 12'hfff;
rom[87665] = 12'hfff;
rom[87666] = 12'hfff;
rom[87667] = 12'hfff;
rom[87668] = 12'hfff;
rom[87669] = 12'hfff;
rom[87670] = 12'hfff;
rom[87671] = 12'hfff;
rom[87672] = 12'hfff;
rom[87673] = 12'hfff;
rom[87674] = 12'hfff;
rom[87675] = 12'hfff;
rom[87676] = 12'hfff;
rom[87677] = 12'hfff;
rom[87678] = 12'hfff;
rom[87679] = 12'hfff;
rom[87680] = 12'hfff;
rom[87681] = 12'hfff;
rom[87682] = 12'hfff;
rom[87683] = 12'hfff;
rom[87684] = 12'hfff;
rom[87685] = 12'hfff;
rom[87686] = 12'hfff;
rom[87687] = 12'hfff;
rom[87688] = 12'hfff;
rom[87689] = 12'hfff;
rom[87690] = 12'hfff;
rom[87691] = 12'hfff;
rom[87692] = 12'hfff;
rom[87693] = 12'hfff;
rom[87694] = 12'hfff;
rom[87695] = 12'hfff;
rom[87696] = 12'hfff;
rom[87697] = 12'hfff;
rom[87698] = 12'hfff;
rom[87699] = 12'hfff;
rom[87700] = 12'hfff;
rom[87701] = 12'hfff;
rom[87702] = 12'hfff;
rom[87703] = 12'hfff;
rom[87704] = 12'hfff;
rom[87705] = 12'hfff;
rom[87706] = 12'hfff;
rom[87707] = 12'hfff;
rom[87708] = 12'hfff;
rom[87709] = 12'hfff;
rom[87710] = 12'hfff;
rom[87711] = 12'hfff;
rom[87712] = 12'hfff;
rom[87713] = 12'hfff;
rom[87714] = 12'hfff;
rom[87715] = 12'hfff;
rom[87716] = 12'hfff;
rom[87717] = 12'hfff;
rom[87718] = 12'hfff;
rom[87719] = 12'hfff;
rom[87720] = 12'hfff;
rom[87721] = 12'hfff;
rom[87722] = 12'hfff;
rom[87723] = 12'hfff;
rom[87724] = 12'hfff;
rom[87725] = 12'hfff;
rom[87726] = 12'heee;
rom[87727] = 12'heee;
rom[87728] = 12'heee;
rom[87729] = 12'hddd;
rom[87730] = 12'hddd;
rom[87731] = 12'hddd;
rom[87732] = 12'hccc;
rom[87733] = 12'hccc;
rom[87734] = 12'hccc;
rom[87735] = 12'hccc;
rom[87736] = 12'hccc;
rom[87737] = 12'hbbb;
rom[87738] = 12'hbbb;
rom[87739] = 12'hbbb;
rom[87740] = 12'hbbb;
rom[87741] = 12'hbbb;
rom[87742] = 12'haaa;
rom[87743] = 12'haaa;
rom[87744] = 12'haaa;
rom[87745] = 12'h999;
rom[87746] = 12'h999;
rom[87747] = 12'h999;
rom[87748] = 12'h888;
rom[87749] = 12'h888;
rom[87750] = 12'h888;
rom[87751] = 12'h888;
rom[87752] = 12'h888;
rom[87753] = 12'h888;
rom[87754] = 12'h888;
rom[87755] = 12'h888;
rom[87756] = 12'h888;
rom[87757] = 12'h999;
rom[87758] = 12'h999;
rom[87759] = 12'h999;
rom[87760] = 12'h999;
rom[87761] = 12'h999;
rom[87762] = 12'h999;
rom[87763] = 12'h999;
rom[87764] = 12'h999;
rom[87765] = 12'h999;
rom[87766] = 12'h999;
rom[87767] = 12'h888;
rom[87768] = 12'h888;
rom[87769] = 12'h888;
rom[87770] = 12'h777;
rom[87771] = 12'h777;
rom[87772] = 12'h777;
rom[87773] = 12'h777;
rom[87774] = 12'h777;
rom[87775] = 12'h777;
rom[87776] = 12'h666;
rom[87777] = 12'h666;
rom[87778] = 12'h666;
rom[87779] = 12'h666;
rom[87780] = 12'h666;
rom[87781] = 12'h666;
rom[87782] = 12'h555;
rom[87783] = 12'h555;
rom[87784] = 12'h555;
rom[87785] = 12'h555;
rom[87786] = 12'h555;
rom[87787] = 12'h666;
rom[87788] = 12'h666;
rom[87789] = 12'h666;
rom[87790] = 12'h666;
rom[87791] = 12'h666;
rom[87792] = 12'h555;
rom[87793] = 12'h555;
rom[87794] = 12'h555;
rom[87795] = 12'h555;
rom[87796] = 12'h555;
rom[87797] = 12'h555;
rom[87798] = 12'h555;
rom[87799] = 12'h555;
rom[87800] = 12'h666;
rom[87801] = 12'h666;
rom[87802] = 12'h666;
rom[87803] = 12'h666;
rom[87804] = 12'h555;
rom[87805] = 12'h555;
rom[87806] = 12'h555;
rom[87807] = 12'h555;
rom[87808] = 12'h555;
rom[87809] = 12'h555;
rom[87810] = 12'h444;
rom[87811] = 12'h444;
rom[87812] = 12'h444;
rom[87813] = 12'h444;
rom[87814] = 12'h444;
rom[87815] = 12'h444;
rom[87816] = 12'h555;
rom[87817] = 12'h555;
rom[87818] = 12'h666;
rom[87819] = 12'h777;
rom[87820] = 12'h777;
rom[87821] = 12'h666;
rom[87822] = 12'h666;
rom[87823] = 12'h555;
rom[87824] = 12'h444;
rom[87825] = 12'h333;
rom[87826] = 12'h333;
rom[87827] = 12'h222;
rom[87828] = 12'h333;
rom[87829] = 12'h333;
rom[87830] = 12'h222;
rom[87831] = 12'h222;
rom[87832] = 12'h222;
rom[87833] = 12'h111;
rom[87834] = 12'h111;
rom[87835] = 12'h111;
rom[87836] = 12'h  0;
rom[87837] = 12'h  0;
rom[87838] = 12'h  0;
rom[87839] = 12'h  0;
rom[87840] = 12'h  0;
rom[87841] = 12'h  0;
rom[87842] = 12'h  0;
rom[87843] = 12'h  0;
rom[87844] = 12'h  0;
rom[87845] = 12'h  0;
rom[87846] = 12'h  0;
rom[87847] = 12'h  0;
rom[87848] = 12'h  0;
rom[87849] = 12'h  0;
rom[87850] = 12'h  0;
rom[87851] = 12'h  0;
rom[87852] = 12'h  0;
rom[87853] = 12'h  0;
rom[87854] = 12'h  0;
rom[87855] = 12'h  0;
rom[87856] = 12'h  0;
rom[87857] = 12'h  0;
rom[87858] = 12'h  0;
rom[87859] = 12'h  0;
rom[87860] = 12'h  0;
rom[87861] = 12'h  0;
rom[87862] = 12'h  0;
rom[87863] = 12'h  0;
rom[87864] = 12'h  0;
rom[87865] = 12'h  0;
rom[87866] = 12'h  0;
rom[87867] = 12'h  0;
rom[87868] = 12'h  0;
rom[87869] = 12'h111;
rom[87870] = 12'h111;
rom[87871] = 12'h111;
rom[87872] = 12'h111;
rom[87873] = 12'h111;
rom[87874] = 12'h222;
rom[87875] = 12'h222;
rom[87876] = 12'h222;
rom[87877] = 12'h333;
rom[87878] = 12'h444;
rom[87879] = 12'h555;
rom[87880] = 12'h777;
rom[87881] = 12'h888;
rom[87882] = 12'h999;
rom[87883] = 12'h999;
rom[87884] = 12'h888;
rom[87885] = 12'h777;
rom[87886] = 12'h777;
rom[87887] = 12'h777;
rom[87888] = 12'h666;
rom[87889] = 12'h777;
rom[87890] = 12'h777;
rom[87891] = 12'h777;
rom[87892] = 12'h777;
rom[87893] = 12'h777;
rom[87894] = 12'h777;
rom[87895] = 12'h777;
rom[87896] = 12'h777;
rom[87897] = 12'h777;
rom[87898] = 12'h777;
rom[87899] = 12'h777;
rom[87900] = 12'h888;
rom[87901] = 12'h999;
rom[87902] = 12'haaa;
rom[87903] = 12'hbbb;
rom[87904] = 12'hbbb;
rom[87905] = 12'hbbb;
rom[87906] = 12'haaa;
rom[87907] = 12'h999;
rom[87908] = 12'h999;
rom[87909] = 12'h999;
rom[87910] = 12'h999;
rom[87911] = 12'h999;
rom[87912] = 12'h999;
rom[87913] = 12'h999;
rom[87914] = 12'h999;
rom[87915] = 12'h999;
rom[87916] = 12'h999;
rom[87917] = 12'haaa;
rom[87918] = 12'haaa;
rom[87919] = 12'haaa;
rom[87920] = 12'haaa;
rom[87921] = 12'hbbb;
rom[87922] = 12'hbbb;
rom[87923] = 12'hbbb;
rom[87924] = 12'hbbb;
rom[87925] = 12'hbbb;
rom[87926] = 12'hbbb;
rom[87927] = 12'hbbb;
rom[87928] = 12'haaa;
rom[87929] = 12'haaa;
rom[87930] = 12'haaa;
rom[87931] = 12'haaa;
rom[87932] = 12'hbbb;
rom[87933] = 12'hbbb;
rom[87934] = 12'hbbb;
rom[87935] = 12'hbbb;
rom[87936] = 12'hccc;
rom[87937] = 12'hddd;
rom[87938] = 12'heee;
rom[87939] = 12'heee;
rom[87940] = 12'hfff;
rom[87941] = 12'heee;
rom[87942] = 12'heee;
rom[87943] = 12'heee;
rom[87944] = 12'hddd;
rom[87945] = 12'hccc;
rom[87946] = 12'hbbb;
rom[87947] = 12'haaa;
rom[87948] = 12'h999;
rom[87949] = 12'h999;
rom[87950] = 12'h999;
rom[87951] = 12'h999;
rom[87952] = 12'haaa;
rom[87953] = 12'h999;
rom[87954] = 12'h999;
rom[87955] = 12'haaa;
rom[87956] = 12'haaa;
rom[87957] = 12'haaa;
rom[87958] = 12'haaa;
rom[87959] = 12'hbbb;
rom[87960] = 12'hbbb;
rom[87961] = 12'hbbb;
rom[87962] = 12'hbbb;
rom[87963] = 12'hbbb;
rom[87964] = 12'hbbb;
rom[87965] = 12'hbbb;
rom[87966] = 12'hbbb;
rom[87967] = 12'hbbb;
rom[87968] = 12'hbbb;
rom[87969] = 12'haaa;
rom[87970] = 12'haaa;
rom[87971] = 12'haaa;
rom[87972] = 12'h999;
rom[87973] = 12'h999;
rom[87974] = 12'h888;
rom[87975] = 12'h888;
rom[87976] = 12'h888;
rom[87977] = 12'h777;
rom[87978] = 12'h666;
rom[87979] = 12'h666;
rom[87980] = 12'h555;
rom[87981] = 12'h555;
rom[87982] = 12'h555;
rom[87983] = 12'h555;
rom[87984] = 12'h444;
rom[87985] = 12'h444;
rom[87986] = 12'h444;
rom[87987] = 12'h333;
rom[87988] = 12'h333;
rom[87989] = 12'h333;
rom[87990] = 12'h333;
rom[87991] = 12'h333;
rom[87992] = 12'h222;
rom[87993] = 12'h222;
rom[87994] = 12'h222;
rom[87995] = 12'h222;
rom[87996] = 12'h222;
rom[87997] = 12'h222;
rom[87998] = 12'h222;
rom[87999] = 12'h222;
rom[88000] = 12'hfff;
rom[88001] = 12'hfff;
rom[88002] = 12'hfff;
rom[88003] = 12'hfff;
rom[88004] = 12'hfff;
rom[88005] = 12'hfff;
rom[88006] = 12'hfff;
rom[88007] = 12'hfff;
rom[88008] = 12'hfff;
rom[88009] = 12'hfff;
rom[88010] = 12'hfff;
rom[88011] = 12'hfff;
rom[88012] = 12'hfff;
rom[88013] = 12'hfff;
rom[88014] = 12'hfff;
rom[88015] = 12'hfff;
rom[88016] = 12'hfff;
rom[88017] = 12'hfff;
rom[88018] = 12'hfff;
rom[88019] = 12'hfff;
rom[88020] = 12'hfff;
rom[88021] = 12'hfff;
rom[88022] = 12'hfff;
rom[88023] = 12'hfff;
rom[88024] = 12'hfff;
rom[88025] = 12'hfff;
rom[88026] = 12'hfff;
rom[88027] = 12'hfff;
rom[88028] = 12'hfff;
rom[88029] = 12'hfff;
rom[88030] = 12'hfff;
rom[88031] = 12'hfff;
rom[88032] = 12'hfff;
rom[88033] = 12'hfff;
rom[88034] = 12'hfff;
rom[88035] = 12'hfff;
rom[88036] = 12'hfff;
rom[88037] = 12'hfff;
rom[88038] = 12'hfff;
rom[88039] = 12'hfff;
rom[88040] = 12'hfff;
rom[88041] = 12'hfff;
rom[88042] = 12'hfff;
rom[88043] = 12'hfff;
rom[88044] = 12'hfff;
rom[88045] = 12'hfff;
rom[88046] = 12'hfff;
rom[88047] = 12'hfff;
rom[88048] = 12'hfff;
rom[88049] = 12'hfff;
rom[88050] = 12'hfff;
rom[88051] = 12'hfff;
rom[88052] = 12'hfff;
rom[88053] = 12'hfff;
rom[88054] = 12'hfff;
rom[88055] = 12'hfff;
rom[88056] = 12'hfff;
rom[88057] = 12'hfff;
rom[88058] = 12'hfff;
rom[88059] = 12'hfff;
rom[88060] = 12'hfff;
rom[88061] = 12'hfff;
rom[88062] = 12'hfff;
rom[88063] = 12'hfff;
rom[88064] = 12'hfff;
rom[88065] = 12'hfff;
rom[88066] = 12'hfff;
rom[88067] = 12'hfff;
rom[88068] = 12'hfff;
rom[88069] = 12'hfff;
rom[88070] = 12'hfff;
rom[88071] = 12'hfff;
rom[88072] = 12'hfff;
rom[88073] = 12'hfff;
rom[88074] = 12'hfff;
rom[88075] = 12'hfff;
rom[88076] = 12'hfff;
rom[88077] = 12'hfff;
rom[88078] = 12'hfff;
rom[88079] = 12'hfff;
rom[88080] = 12'hfff;
rom[88081] = 12'hfff;
rom[88082] = 12'hfff;
rom[88083] = 12'hfff;
rom[88084] = 12'hfff;
rom[88085] = 12'hfff;
rom[88086] = 12'hfff;
rom[88087] = 12'hfff;
rom[88088] = 12'hfff;
rom[88089] = 12'hfff;
rom[88090] = 12'hfff;
rom[88091] = 12'hfff;
rom[88092] = 12'hfff;
rom[88093] = 12'hfff;
rom[88094] = 12'hfff;
rom[88095] = 12'hfff;
rom[88096] = 12'hfff;
rom[88097] = 12'hfff;
rom[88098] = 12'hfff;
rom[88099] = 12'hfff;
rom[88100] = 12'hfff;
rom[88101] = 12'hfff;
rom[88102] = 12'hfff;
rom[88103] = 12'hfff;
rom[88104] = 12'hfff;
rom[88105] = 12'hfff;
rom[88106] = 12'hfff;
rom[88107] = 12'hfff;
rom[88108] = 12'hfff;
rom[88109] = 12'hfff;
rom[88110] = 12'hfff;
rom[88111] = 12'hfff;
rom[88112] = 12'hfff;
rom[88113] = 12'hfff;
rom[88114] = 12'hfff;
rom[88115] = 12'hfff;
rom[88116] = 12'hfff;
rom[88117] = 12'hfff;
rom[88118] = 12'hfff;
rom[88119] = 12'hfff;
rom[88120] = 12'hfff;
rom[88121] = 12'hfff;
rom[88122] = 12'hfff;
rom[88123] = 12'hfff;
rom[88124] = 12'hfff;
rom[88125] = 12'hfff;
rom[88126] = 12'hfff;
rom[88127] = 12'hfff;
rom[88128] = 12'heee;
rom[88129] = 12'heee;
rom[88130] = 12'hddd;
rom[88131] = 12'hddd;
rom[88132] = 12'hddd;
rom[88133] = 12'hccc;
rom[88134] = 12'hccc;
rom[88135] = 12'hccc;
rom[88136] = 12'hccc;
rom[88137] = 12'hbbb;
rom[88138] = 12'hbbb;
rom[88139] = 12'hbbb;
rom[88140] = 12'hbbb;
rom[88141] = 12'haaa;
rom[88142] = 12'haaa;
rom[88143] = 12'haaa;
rom[88144] = 12'h999;
rom[88145] = 12'h999;
rom[88146] = 12'h999;
rom[88147] = 12'h999;
rom[88148] = 12'h888;
rom[88149] = 12'h888;
rom[88150] = 12'h888;
rom[88151] = 12'h999;
rom[88152] = 12'h888;
rom[88153] = 12'h888;
rom[88154] = 12'h777;
rom[88155] = 12'h777;
rom[88156] = 12'h777;
rom[88157] = 12'h888;
rom[88158] = 12'h888;
rom[88159] = 12'h888;
rom[88160] = 12'h888;
rom[88161] = 12'h999;
rom[88162] = 12'h999;
rom[88163] = 12'h999;
rom[88164] = 12'h999;
rom[88165] = 12'h999;
rom[88166] = 12'h999;
rom[88167] = 12'h999;
rom[88168] = 12'h888;
rom[88169] = 12'h888;
rom[88170] = 12'h888;
rom[88171] = 12'h777;
rom[88172] = 12'h777;
rom[88173] = 12'h777;
rom[88174] = 12'h777;
rom[88175] = 12'h777;
rom[88176] = 12'h666;
rom[88177] = 12'h666;
rom[88178] = 12'h666;
rom[88179] = 12'h666;
rom[88180] = 12'h666;
rom[88181] = 12'h666;
rom[88182] = 12'h555;
rom[88183] = 12'h555;
rom[88184] = 12'h666;
rom[88185] = 12'h666;
rom[88186] = 12'h666;
rom[88187] = 12'h666;
rom[88188] = 12'h666;
rom[88189] = 12'h666;
rom[88190] = 12'h666;
rom[88191] = 12'h666;
rom[88192] = 12'h666;
rom[88193] = 12'h555;
rom[88194] = 12'h555;
rom[88195] = 12'h555;
rom[88196] = 12'h555;
rom[88197] = 12'h555;
rom[88198] = 12'h555;
rom[88199] = 12'h555;
rom[88200] = 12'h666;
rom[88201] = 12'h666;
rom[88202] = 12'h666;
rom[88203] = 12'h555;
rom[88204] = 12'h555;
rom[88205] = 12'h555;
rom[88206] = 12'h555;
rom[88207] = 12'h555;
rom[88208] = 12'h555;
rom[88209] = 12'h444;
rom[88210] = 12'h444;
rom[88211] = 12'h444;
rom[88212] = 12'h444;
rom[88213] = 12'h444;
rom[88214] = 12'h444;
rom[88215] = 12'h444;
rom[88216] = 12'h555;
rom[88217] = 12'h555;
rom[88218] = 12'h666;
rom[88219] = 12'h666;
rom[88220] = 12'h777;
rom[88221] = 12'h777;
rom[88222] = 12'h666;
rom[88223] = 12'h666;
rom[88224] = 12'h444;
rom[88225] = 12'h444;
rom[88226] = 12'h333;
rom[88227] = 12'h333;
rom[88228] = 12'h333;
rom[88229] = 12'h333;
rom[88230] = 12'h333;
rom[88231] = 12'h222;
rom[88232] = 12'h222;
rom[88233] = 12'h222;
rom[88234] = 12'h111;
rom[88235] = 12'h111;
rom[88236] = 12'h111;
rom[88237] = 12'h111;
rom[88238] = 12'h  0;
rom[88239] = 12'h  0;
rom[88240] = 12'h  0;
rom[88241] = 12'h  0;
rom[88242] = 12'h  0;
rom[88243] = 12'h  0;
rom[88244] = 12'h  0;
rom[88245] = 12'h  0;
rom[88246] = 12'h  0;
rom[88247] = 12'h  0;
rom[88248] = 12'h  0;
rom[88249] = 12'h  0;
rom[88250] = 12'h  0;
rom[88251] = 12'h  0;
rom[88252] = 12'h  0;
rom[88253] = 12'h  0;
rom[88254] = 12'h  0;
rom[88255] = 12'h  0;
rom[88256] = 12'h  0;
rom[88257] = 12'h  0;
rom[88258] = 12'h  0;
rom[88259] = 12'h  0;
rom[88260] = 12'h  0;
rom[88261] = 12'h  0;
rom[88262] = 12'h  0;
rom[88263] = 12'h  0;
rom[88264] = 12'h  0;
rom[88265] = 12'h  0;
rom[88266] = 12'h  0;
rom[88267] = 12'h  0;
rom[88268] = 12'h  0;
rom[88269] = 12'h111;
rom[88270] = 12'h111;
rom[88271] = 12'h111;
rom[88272] = 12'h111;
rom[88273] = 12'h111;
rom[88274] = 12'h222;
rom[88275] = 12'h222;
rom[88276] = 12'h333;
rom[88277] = 12'h333;
rom[88278] = 12'h444;
rom[88279] = 12'h555;
rom[88280] = 12'h777;
rom[88281] = 12'h888;
rom[88282] = 12'h999;
rom[88283] = 12'h888;
rom[88284] = 12'h888;
rom[88285] = 12'h777;
rom[88286] = 12'h777;
rom[88287] = 12'h777;
rom[88288] = 12'h666;
rom[88289] = 12'h777;
rom[88290] = 12'h777;
rom[88291] = 12'h888;
rom[88292] = 12'h888;
rom[88293] = 12'h888;
rom[88294] = 12'h777;
rom[88295] = 12'h777;
rom[88296] = 12'h777;
rom[88297] = 12'h777;
rom[88298] = 12'h777;
rom[88299] = 12'h777;
rom[88300] = 12'h888;
rom[88301] = 12'h999;
rom[88302] = 12'hbbb;
rom[88303] = 12'hccc;
rom[88304] = 12'hbbb;
rom[88305] = 12'haaa;
rom[88306] = 12'h999;
rom[88307] = 12'h999;
rom[88308] = 12'h888;
rom[88309] = 12'h888;
rom[88310] = 12'h888;
rom[88311] = 12'h888;
rom[88312] = 12'h777;
rom[88313] = 12'h777;
rom[88314] = 12'h666;
rom[88315] = 12'h666;
rom[88316] = 12'h666;
rom[88317] = 12'h666;
rom[88318] = 12'h777;
rom[88319] = 12'h777;
rom[88320] = 12'h777;
rom[88321] = 12'h888;
rom[88322] = 12'h888;
rom[88323] = 12'h999;
rom[88324] = 12'h999;
rom[88325] = 12'h999;
rom[88326] = 12'h999;
rom[88327] = 12'h999;
rom[88328] = 12'h999;
rom[88329] = 12'h999;
rom[88330] = 12'haaa;
rom[88331] = 12'haaa;
rom[88332] = 12'haaa;
rom[88333] = 12'haaa;
rom[88334] = 12'haaa;
rom[88335] = 12'hbbb;
rom[88336] = 12'hbbb;
rom[88337] = 12'hbbb;
rom[88338] = 12'hccc;
rom[88339] = 12'hddd;
rom[88340] = 12'heee;
rom[88341] = 12'heee;
rom[88342] = 12'heee;
rom[88343] = 12'heee;
rom[88344] = 12'heee;
rom[88345] = 12'heee;
rom[88346] = 12'hddd;
rom[88347] = 12'hbbb;
rom[88348] = 12'haaa;
rom[88349] = 12'h999;
rom[88350] = 12'h888;
rom[88351] = 12'h888;
rom[88352] = 12'h777;
rom[88353] = 12'h777;
rom[88354] = 12'h777;
rom[88355] = 12'h777;
rom[88356] = 12'h777;
rom[88357] = 12'h777;
rom[88358] = 12'h777;
rom[88359] = 12'h777;
rom[88360] = 12'h777;
rom[88361] = 12'h888;
rom[88362] = 12'h888;
rom[88363] = 12'h888;
rom[88364] = 12'h999;
rom[88365] = 12'h999;
rom[88366] = 12'h999;
rom[88367] = 12'haaa;
rom[88368] = 12'haaa;
rom[88369] = 12'haaa;
rom[88370] = 12'hbbb;
rom[88371] = 12'haaa;
rom[88372] = 12'haaa;
rom[88373] = 12'haaa;
rom[88374] = 12'haaa;
rom[88375] = 12'haaa;
rom[88376] = 12'haaa;
rom[88377] = 12'haaa;
rom[88378] = 12'h999;
rom[88379] = 12'h888;
rom[88380] = 12'h777;
rom[88381] = 12'h777;
rom[88382] = 12'h666;
rom[88383] = 12'h666;
rom[88384] = 12'h666;
rom[88385] = 12'h666;
rom[88386] = 12'h555;
rom[88387] = 12'h555;
rom[88388] = 12'h444;
rom[88389] = 12'h444;
rom[88390] = 12'h333;
rom[88391] = 12'h333;
rom[88392] = 12'h333;
rom[88393] = 12'h333;
rom[88394] = 12'h333;
rom[88395] = 12'h333;
rom[88396] = 12'h333;
rom[88397] = 12'h222;
rom[88398] = 12'h222;
rom[88399] = 12'h222;
rom[88400] = 12'hfff;
rom[88401] = 12'hfff;
rom[88402] = 12'hfff;
rom[88403] = 12'hfff;
rom[88404] = 12'hfff;
rom[88405] = 12'hfff;
rom[88406] = 12'hfff;
rom[88407] = 12'hfff;
rom[88408] = 12'hfff;
rom[88409] = 12'hfff;
rom[88410] = 12'hfff;
rom[88411] = 12'hfff;
rom[88412] = 12'hfff;
rom[88413] = 12'hfff;
rom[88414] = 12'hfff;
rom[88415] = 12'hfff;
rom[88416] = 12'hfff;
rom[88417] = 12'hfff;
rom[88418] = 12'hfff;
rom[88419] = 12'hfff;
rom[88420] = 12'hfff;
rom[88421] = 12'hfff;
rom[88422] = 12'hfff;
rom[88423] = 12'hfff;
rom[88424] = 12'hfff;
rom[88425] = 12'hfff;
rom[88426] = 12'hfff;
rom[88427] = 12'hfff;
rom[88428] = 12'hfff;
rom[88429] = 12'hfff;
rom[88430] = 12'hfff;
rom[88431] = 12'hfff;
rom[88432] = 12'hfff;
rom[88433] = 12'hfff;
rom[88434] = 12'hfff;
rom[88435] = 12'hfff;
rom[88436] = 12'hfff;
rom[88437] = 12'hfff;
rom[88438] = 12'hfff;
rom[88439] = 12'hfff;
rom[88440] = 12'hfff;
rom[88441] = 12'hfff;
rom[88442] = 12'hfff;
rom[88443] = 12'hfff;
rom[88444] = 12'hfff;
rom[88445] = 12'hfff;
rom[88446] = 12'hfff;
rom[88447] = 12'hfff;
rom[88448] = 12'hfff;
rom[88449] = 12'hfff;
rom[88450] = 12'hfff;
rom[88451] = 12'hfff;
rom[88452] = 12'hfff;
rom[88453] = 12'hfff;
rom[88454] = 12'hfff;
rom[88455] = 12'hfff;
rom[88456] = 12'hfff;
rom[88457] = 12'hfff;
rom[88458] = 12'hfff;
rom[88459] = 12'hfff;
rom[88460] = 12'hfff;
rom[88461] = 12'hfff;
rom[88462] = 12'hfff;
rom[88463] = 12'hfff;
rom[88464] = 12'hfff;
rom[88465] = 12'hfff;
rom[88466] = 12'hfff;
rom[88467] = 12'hfff;
rom[88468] = 12'hfff;
rom[88469] = 12'hfff;
rom[88470] = 12'hfff;
rom[88471] = 12'hfff;
rom[88472] = 12'hfff;
rom[88473] = 12'hfff;
rom[88474] = 12'hfff;
rom[88475] = 12'hfff;
rom[88476] = 12'hfff;
rom[88477] = 12'hfff;
rom[88478] = 12'hfff;
rom[88479] = 12'hfff;
rom[88480] = 12'hfff;
rom[88481] = 12'hfff;
rom[88482] = 12'hfff;
rom[88483] = 12'hfff;
rom[88484] = 12'hfff;
rom[88485] = 12'hfff;
rom[88486] = 12'hfff;
rom[88487] = 12'hfff;
rom[88488] = 12'hfff;
rom[88489] = 12'hfff;
rom[88490] = 12'hfff;
rom[88491] = 12'hfff;
rom[88492] = 12'hfff;
rom[88493] = 12'hfff;
rom[88494] = 12'hfff;
rom[88495] = 12'hfff;
rom[88496] = 12'hfff;
rom[88497] = 12'hfff;
rom[88498] = 12'hfff;
rom[88499] = 12'hfff;
rom[88500] = 12'hfff;
rom[88501] = 12'hfff;
rom[88502] = 12'hfff;
rom[88503] = 12'hfff;
rom[88504] = 12'hfff;
rom[88505] = 12'hfff;
rom[88506] = 12'hfff;
rom[88507] = 12'hfff;
rom[88508] = 12'hfff;
rom[88509] = 12'hfff;
rom[88510] = 12'hfff;
rom[88511] = 12'hfff;
rom[88512] = 12'hfff;
rom[88513] = 12'hfff;
rom[88514] = 12'hfff;
rom[88515] = 12'hfff;
rom[88516] = 12'hfff;
rom[88517] = 12'hfff;
rom[88518] = 12'hfff;
rom[88519] = 12'hfff;
rom[88520] = 12'hfff;
rom[88521] = 12'hfff;
rom[88522] = 12'hfff;
rom[88523] = 12'hfff;
rom[88524] = 12'hfff;
rom[88525] = 12'hfff;
rom[88526] = 12'hfff;
rom[88527] = 12'hfff;
rom[88528] = 12'heee;
rom[88529] = 12'heee;
rom[88530] = 12'hddd;
rom[88531] = 12'hddd;
rom[88532] = 12'hddd;
rom[88533] = 12'hddd;
rom[88534] = 12'hccc;
rom[88535] = 12'hccc;
rom[88536] = 12'hccc;
rom[88537] = 12'hccc;
rom[88538] = 12'hbbb;
rom[88539] = 12'hbbb;
rom[88540] = 12'hbbb;
rom[88541] = 12'haaa;
rom[88542] = 12'haaa;
rom[88543] = 12'h999;
rom[88544] = 12'h999;
rom[88545] = 12'h999;
rom[88546] = 12'h999;
rom[88547] = 12'h888;
rom[88548] = 12'h888;
rom[88549] = 12'h888;
rom[88550] = 12'h888;
rom[88551] = 12'h888;
rom[88552] = 12'h888;
rom[88553] = 12'h888;
rom[88554] = 12'h777;
rom[88555] = 12'h777;
rom[88556] = 12'h777;
rom[88557] = 12'h777;
rom[88558] = 12'h777;
rom[88559] = 12'h777;
rom[88560] = 12'h888;
rom[88561] = 12'h888;
rom[88562] = 12'h888;
rom[88563] = 12'h888;
rom[88564] = 12'h999;
rom[88565] = 12'h999;
rom[88566] = 12'h999;
rom[88567] = 12'h999;
rom[88568] = 12'h888;
rom[88569] = 12'h888;
rom[88570] = 12'h888;
rom[88571] = 12'h888;
rom[88572] = 12'h888;
rom[88573] = 12'h777;
rom[88574] = 12'h777;
rom[88575] = 12'h777;
rom[88576] = 12'h777;
rom[88577] = 12'h666;
rom[88578] = 12'h666;
rom[88579] = 12'h666;
rom[88580] = 12'h666;
rom[88581] = 12'h666;
rom[88582] = 12'h666;
rom[88583] = 12'h666;
rom[88584] = 12'h666;
rom[88585] = 12'h666;
rom[88586] = 12'h666;
rom[88587] = 12'h666;
rom[88588] = 12'h666;
rom[88589] = 12'h666;
rom[88590] = 12'h666;
rom[88591] = 12'h666;
rom[88592] = 12'h666;
rom[88593] = 12'h666;
rom[88594] = 12'h555;
rom[88595] = 12'h555;
rom[88596] = 12'h555;
rom[88597] = 12'h555;
rom[88598] = 12'h555;
rom[88599] = 12'h555;
rom[88600] = 12'h666;
rom[88601] = 12'h666;
rom[88602] = 12'h666;
rom[88603] = 12'h555;
rom[88604] = 12'h555;
rom[88605] = 12'h555;
rom[88606] = 12'h555;
rom[88607] = 12'h555;
rom[88608] = 12'h555;
rom[88609] = 12'h444;
rom[88610] = 12'h444;
rom[88611] = 12'h444;
rom[88612] = 12'h444;
rom[88613] = 12'h444;
rom[88614] = 12'h444;
rom[88615] = 12'h444;
rom[88616] = 12'h444;
rom[88617] = 12'h555;
rom[88618] = 12'h555;
rom[88619] = 12'h666;
rom[88620] = 12'h666;
rom[88621] = 12'h777;
rom[88622] = 12'h777;
rom[88623] = 12'h777;
rom[88624] = 12'h666;
rom[88625] = 12'h555;
rom[88626] = 12'h444;
rom[88627] = 12'h333;
rom[88628] = 12'h333;
rom[88629] = 12'h333;
rom[88630] = 12'h333;
rom[88631] = 12'h333;
rom[88632] = 12'h222;
rom[88633] = 12'h222;
rom[88634] = 12'h222;
rom[88635] = 12'h111;
rom[88636] = 12'h111;
rom[88637] = 12'h111;
rom[88638] = 12'h111;
rom[88639] = 12'h  0;
rom[88640] = 12'h  0;
rom[88641] = 12'h  0;
rom[88642] = 12'h  0;
rom[88643] = 12'h  0;
rom[88644] = 12'h  0;
rom[88645] = 12'h  0;
rom[88646] = 12'h  0;
rom[88647] = 12'h  0;
rom[88648] = 12'h  0;
rom[88649] = 12'h  0;
rom[88650] = 12'h  0;
rom[88651] = 12'h  0;
rom[88652] = 12'h  0;
rom[88653] = 12'h  0;
rom[88654] = 12'h  0;
rom[88655] = 12'h  0;
rom[88656] = 12'h  0;
rom[88657] = 12'h  0;
rom[88658] = 12'h  0;
rom[88659] = 12'h  0;
rom[88660] = 12'h  0;
rom[88661] = 12'h  0;
rom[88662] = 12'h  0;
rom[88663] = 12'h  0;
rom[88664] = 12'h  0;
rom[88665] = 12'h  0;
rom[88666] = 12'h  0;
rom[88667] = 12'h  0;
rom[88668] = 12'h111;
rom[88669] = 12'h111;
rom[88670] = 12'h111;
rom[88671] = 12'h111;
rom[88672] = 12'h111;
rom[88673] = 12'h111;
rom[88674] = 12'h222;
rom[88675] = 12'h222;
rom[88676] = 12'h333;
rom[88677] = 12'h333;
rom[88678] = 12'h444;
rom[88679] = 12'h555;
rom[88680] = 12'h777;
rom[88681] = 12'h888;
rom[88682] = 12'h999;
rom[88683] = 12'h888;
rom[88684] = 12'h888;
rom[88685] = 12'h777;
rom[88686] = 12'h777;
rom[88687] = 12'h777;
rom[88688] = 12'h666;
rom[88689] = 12'h777;
rom[88690] = 12'h777;
rom[88691] = 12'h777;
rom[88692] = 12'h888;
rom[88693] = 12'h888;
rom[88694] = 12'h888;
rom[88695] = 12'h888;
rom[88696] = 12'h777;
rom[88697] = 12'h777;
rom[88698] = 12'h777;
rom[88699] = 12'h888;
rom[88700] = 12'h999;
rom[88701] = 12'haaa;
rom[88702] = 12'hbbb;
rom[88703] = 12'hccc;
rom[88704] = 12'hbbb;
rom[88705] = 12'haaa;
rom[88706] = 12'h999;
rom[88707] = 12'h888;
rom[88708] = 12'h888;
rom[88709] = 12'h777;
rom[88710] = 12'h777;
rom[88711] = 12'h666;
rom[88712] = 12'h666;
rom[88713] = 12'h666;
rom[88714] = 12'h666;
rom[88715] = 12'h555;
rom[88716] = 12'h555;
rom[88717] = 12'h555;
rom[88718] = 12'h555;
rom[88719] = 12'h555;
rom[88720] = 12'h555;
rom[88721] = 12'h555;
rom[88722] = 12'h555;
rom[88723] = 12'h666;
rom[88724] = 12'h666;
rom[88725] = 12'h666;
rom[88726] = 12'h777;
rom[88727] = 12'h777;
rom[88728] = 12'h777;
rom[88729] = 12'h777;
rom[88730] = 12'h777;
rom[88731] = 12'h777;
rom[88732] = 12'h777;
rom[88733] = 12'h888;
rom[88734] = 12'h888;
rom[88735] = 12'h888;
rom[88736] = 12'h999;
rom[88737] = 12'h999;
rom[88738] = 12'haaa;
rom[88739] = 12'haaa;
rom[88740] = 12'hbbb;
rom[88741] = 12'hccc;
rom[88742] = 12'hddd;
rom[88743] = 12'hddd;
rom[88744] = 12'heee;
rom[88745] = 12'hfff;
rom[88746] = 12'hfff;
rom[88747] = 12'heee;
rom[88748] = 12'hddd;
rom[88749] = 12'hccc;
rom[88750] = 12'hbbb;
rom[88751] = 12'haaa;
rom[88752] = 12'h888;
rom[88753] = 12'h888;
rom[88754] = 12'h777;
rom[88755] = 12'h666;
rom[88756] = 12'h555;
rom[88757] = 12'h555;
rom[88758] = 12'h555;
rom[88759] = 12'h555;
rom[88760] = 12'h555;
rom[88761] = 12'h555;
rom[88762] = 12'h555;
rom[88763] = 12'h555;
rom[88764] = 12'h555;
rom[88765] = 12'h666;
rom[88766] = 12'h666;
rom[88767] = 12'h666;
rom[88768] = 12'h777;
rom[88769] = 12'h777;
rom[88770] = 12'h777;
rom[88771] = 12'h888;
rom[88772] = 12'h888;
rom[88773] = 12'h999;
rom[88774] = 12'h999;
rom[88775] = 12'h999;
rom[88776] = 12'haaa;
rom[88777] = 12'haaa;
rom[88778] = 12'haaa;
rom[88779] = 12'haaa;
rom[88780] = 12'haaa;
rom[88781] = 12'h999;
rom[88782] = 12'h999;
rom[88783] = 12'h999;
rom[88784] = 12'h888;
rom[88785] = 12'h888;
rom[88786] = 12'h777;
rom[88787] = 12'h666;
rom[88788] = 12'h666;
rom[88789] = 12'h555;
rom[88790] = 12'h555;
rom[88791] = 12'h555;
rom[88792] = 12'h444;
rom[88793] = 12'h444;
rom[88794] = 12'h333;
rom[88795] = 12'h333;
rom[88796] = 12'h333;
rom[88797] = 12'h333;
rom[88798] = 12'h222;
rom[88799] = 12'h222;
rom[88800] = 12'hfff;
rom[88801] = 12'hfff;
rom[88802] = 12'hfff;
rom[88803] = 12'hfff;
rom[88804] = 12'hfff;
rom[88805] = 12'hfff;
rom[88806] = 12'hfff;
rom[88807] = 12'hfff;
rom[88808] = 12'hfff;
rom[88809] = 12'hfff;
rom[88810] = 12'hfff;
rom[88811] = 12'hfff;
rom[88812] = 12'hfff;
rom[88813] = 12'hfff;
rom[88814] = 12'hfff;
rom[88815] = 12'hfff;
rom[88816] = 12'hfff;
rom[88817] = 12'hfff;
rom[88818] = 12'hfff;
rom[88819] = 12'hfff;
rom[88820] = 12'hfff;
rom[88821] = 12'hfff;
rom[88822] = 12'hfff;
rom[88823] = 12'hfff;
rom[88824] = 12'hfff;
rom[88825] = 12'hfff;
rom[88826] = 12'hfff;
rom[88827] = 12'hfff;
rom[88828] = 12'hfff;
rom[88829] = 12'hfff;
rom[88830] = 12'hfff;
rom[88831] = 12'hfff;
rom[88832] = 12'hfff;
rom[88833] = 12'hfff;
rom[88834] = 12'hfff;
rom[88835] = 12'hfff;
rom[88836] = 12'hfff;
rom[88837] = 12'hfff;
rom[88838] = 12'hfff;
rom[88839] = 12'hfff;
rom[88840] = 12'hfff;
rom[88841] = 12'hfff;
rom[88842] = 12'hfff;
rom[88843] = 12'hfff;
rom[88844] = 12'hfff;
rom[88845] = 12'hfff;
rom[88846] = 12'hfff;
rom[88847] = 12'hfff;
rom[88848] = 12'hfff;
rom[88849] = 12'hfff;
rom[88850] = 12'hfff;
rom[88851] = 12'hfff;
rom[88852] = 12'hfff;
rom[88853] = 12'hfff;
rom[88854] = 12'hfff;
rom[88855] = 12'hfff;
rom[88856] = 12'hfff;
rom[88857] = 12'hfff;
rom[88858] = 12'hfff;
rom[88859] = 12'hfff;
rom[88860] = 12'hfff;
rom[88861] = 12'hfff;
rom[88862] = 12'hfff;
rom[88863] = 12'hfff;
rom[88864] = 12'hfff;
rom[88865] = 12'hfff;
rom[88866] = 12'hfff;
rom[88867] = 12'hfff;
rom[88868] = 12'hfff;
rom[88869] = 12'hfff;
rom[88870] = 12'hfff;
rom[88871] = 12'hfff;
rom[88872] = 12'hfff;
rom[88873] = 12'hfff;
rom[88874] = 12'hfff;
rom[88875] = 12'hfff;
rom[88876] = 12'hfff;
rom[88877] = 12'hfff;
rom[88878] = 12'hfff;
rom[88879] = 12'hfff;
rom[88880] = 12'hfff;
rom[88881] = 12'hfff;
rom[88882] = 12'hfff;
rom[88883] = 12'hfff;
rom[88884] = 12'hfff;
rom[88885] = 12'hfff;
rom[88886] = 12'hfff;
rom[88887] = 12'hfff;
rom[88888] = 12'hfff;
rom[88889] = 12'hfff;
rom[88890] = 12'hfff;
rom[88891] = 12'hfff;
rom[88892] = 12'hfff;
rom[88893] = 12'hfff;
rom[88894] = 12'hfff;
rom[88895] = 12'hfff;
rom[88896] = 12'hfff;
rom[88897] = 12'hfff;
rom[88898] = 12'hfff;
rom[88899] = 12'hfff;
rom[88900] = 12'hfff;
rom[88901] = 12'hfff;
rom[88902] = 12'hfff;
rom[88903] = 12'hfff;
rom[88904] = 12'hfff;
rom[88905] = 12'hfff;
rom[88906] = 12'hfff;
rom[88907] = 12'hfff;
rom[88908] = 12'hfff;
rom[88909] = 12'hfff;
rom[88910] = 12'hfff;
rom[88911] = 12'hfff;
rom[88912] = 12'hfff;
rom[88913] = 12'hfff;
rom[88914] = 12'hfff;
rom[88915] = 12'hfff;
rom[88916] = 12'hfff;
rom[88917] = 12'hfff;
rom[88918] = 12'hfff;
rom[88919] = 12'hfff;
rom[88920] = 12'hfff;
rom[88921] = 12'hfff;
rom[88922] = 12'hfff;
rom[88923] = 12'hfff;
rom[88924] = 12'hfff;
rom[88925] = 12'hfff;
rom[88926] = 12'hfff;
rom[88927] = 12'hfff;
rom[88928] = 12'heee;
rom[88929] = 12'heee;
rom[88930] = 12'heee;
rom[88931] = 12'hddd;
rom[88932] = 12'hddd;
rom[88933] = 12'hddd;
rom[88934] = 12'hccc;
rom[88935] = 12'hccc;
rom[88936] = 12'hccc;
rom[88937] = 12'hccc;
rom[88938] = 12'hbbb;
rom[88939] = 12'hbbb;
rom[88940] = 12'hbbb;
rom[88941] = 12'haaa;
rom[88942] = 12'haaa;
rom[88943] = 12'haaa;
rom[88944] = 12'h999;
rom[88945] = 12'h999;
rom[88946] = 12'h999;
rom[88947] = 12'h888;
rom[88948] = 12'h888;
rom[88949] = 12'h888;
rom[88950] = 12'h888;
rom[88951] = 12'h888;
rom[88952] = 12'h888;
rom[88953] = 12'h888;
rom[88954] = 12'h888;
rom[88955] = 12'h777;
rom[88956] = 12'h777;
rom[88957] = 12'h777;
rom[88958] = 12'h777;
rom[88959] = 12'h777;
rom[88960] = 12'h777;
rom[88961] = 12'h777;
rom[88962] = 12'h777;
rom[88963] = 12'h888;
rom[88964] = 12'h888;
rom[88965] = 12'h888;
rom[88966] = 12'h888;
rom[88967] = 12'h888;
rom[88968] = 12'h888;
rom[88969] = 12'h888;
rom[88970] = 12'h888;
rom[88971] = 12'h888;
rom[88972] = 12'h888;
rom[88973] = 12'h888;
rom[88974] = 12'h777;
rom[88975] = 12'h777;
rom[88976] = 12'h777;
rom[88977] = 12'h777;
rom[88978] = 12'h666;
rom[88979] = 12'h666;
rom[88980] = 12'h666;
rom[88981] = 12'h666;
rom[88982] = 12'h666;
rom[88983] = 12'h666;
rom[88984] = 12'h666;
rom[88985] = 12'h666;
rom[88986] = 12'h666;
rom[88987] = 12'h666;
rom[88988] = 12'h666;
rom[88989] = 12'h666;
rom[88990] = 12'h666;
rom[88991] = 12'h666;
rom[88992] = 12'h666;
rom[88993] = 12'h666;
rom[88994] = 12'h666;
rom[88995] = 12'h666;
rom[88996] = 12'h555;
rom[88997] = 12'h555;
rom[88998] = 12'h555;
rom[88999] = 12'h555;
rom[89000] = 12'h666;
rom[89001] = 12'h666;
rom[89002] = 12'h555;
rom[89003] = 12'h555;
rom[89004] = 12'h555;
rom[89005] = 12'h555;
rom[89006] = 12'h555;
rom[89007] = 12'h555;
rom[89008] = 12'h555;
rom[89009] = 12'h444;
rom[89010] = 12'h444;
rom[89011] = 12'h444;
rom[89012] = 12'h444;
rom[89013] = 12'h444;
rom[89014] = 12'h444;
rom[89015] = 12'h333;
rom[89016] = 12'h444;
rom[89017] = 12'h444;
rom[89018] = 12'h444;
rom[89019] = 12'h555;
rom[89020] = 12'h555;
rom[89021] = 12'h666;
rom[89022] = 12'h777;
rom[89023] = 12'h777;
rom[89024] = 12'h777;
rom[89025] = 12'h666;
rom[89026] = 12'h555;
rom[89027] = 12'h444;
rom[89028] = 12'h444;
rom[89029] = 12'h333;
rom[89030] = 12'h333;
rom[89031] = 12'h333;
rom[89032] = 12'h333;
rom[89033] = 12'h222;
rom[89034] = 12'h222;
rom[89035] = 12'h111;
rom[89036] = 12'h111;
rom[89037] = 12'h111;
rom[89038] = 12'h111;
rom[89039] = 12'h111;
rom[89040] = 12'h111;
rom[89041] = 12'h111;
rom[89042] = 12'h111;
rom[89043] = 12'h111;
rom[89044] = 12'h  0;
rom[89045] = 12'h  0;
rom[89046] = 12'h  0;
rom[89047] = 12'h  0;
rom[89048] = 12'h  0;
rom[89049] = 12'h  0;
rom[89050] = 12'h  0;
rom[89051] = 12'h  0;
rom[89052] = 12'h  0;
rom[89053] = 12'h  0;
rom[89054] = 12'h  0;
rom[89055] = 12'h  0;
rom[89056] = 12'h  0;
rom[89057] = 12'h  0;
rom[89058] = 12'h  0;
rom[89059] = 12'h  0;
rom[89060] = 12'h  0;
rom[89061] = 12'h  0;
rom[89062] = 12'h  0;
rom[89063] = 12'h  0;
rom[89064] = 12'h111;
rom[89065] = 12'h111;
rom[89066] = 12'h111;
rom[89067] = 12'h111;
rom[89068] = 12'h111;
rom[89069] = 12'h111;
rom[89070] = 12'h111;
rom[89071] = 12'h111;
rom[89072] = 12'h111;
rom[89073] = 12'h111;
rom[89074] = 12'h222;
rom[89075] = 12'h222;
rom[89076] = 12'h333;
rom[89077] = 12'h333;
rom[89078] = 12'h444;
rom[89079] = 12'h666;
rom[89080] = 12'h777;
rom[89081] = 12'h888;
rom[89082] = 12'h999;
rom[89083] = 12'h888;
rom[89084] = 12'h888;
rom[89085] = 12'h777;
rom[89086] = 12'h777;
rom[89087] = 12'h777;
rom[89088] = 12'h777;
rom[89089] = 12'h777;
rom[89090] = 12'h777;
rom[89091] = 12'h777;
rom[89092] = 12'h777;
rom[89093] = 12'h888;
rom[89094] = 12'h888;
rom[89095] = 12'h888;
rom[89096] = 12'h888;
rom[89097] = 12'h888;
rom[89098] = 12'h777;
rom[89099] = 12'h888;
rom[89100] = 12'haaa;
rom[89101] = 12'hbbb;
rom[89102] = 12'hccc;
rom[89103] = 12'hccc;
rom[89104] = 12'hbbb;
rom[89105] = 12'h999;
rom[89106] = 12'h888;
rom[89107] = 12'h888;
rom[89108] = 12'h777;
rom[89109] = 12'h777;
rom[89110] = 12'h666;
rom[89111] = 12'h666;
rom[89112] = 12'h555;
rom[89113] = 12'h555;
rom[89114] = 12'h555;
rom[89115] = 12'h555;
rom[89116] = 12'h555;
rom[89117] = 12'h555;
rom[89118] = 12'h444;
rom[89119] = 12'h444;
rom[89120] = 12'h444;
rom[89121] = 12'h444;
rom[89122] = 12'h444;
rom[89123] = 12'h444;
rom[89124] = 12'h444;
rom[89125] = 12'h555;
rom[89126] = 12'h555;
rom[89127] = 12'h555;
rom[89128] = 12'h555;
rom[89129] = 12'h555;
rom[89130] = 12'h555;
rom[89131] = 12'h555;
rom[89132] = 12'h555;
rom[89133] = 12'h555;
rom[89134] = 12'h555;
rom[89135] = 12'h555;
rom[89136] = 12'h666;
rom[89137] = 12'h666;
rom[89138] = 12'h777;
rom[89139] = 12'h777;
rom[89140] = 12'h777;
rom[89141] = 12'h888;
rom[89142] = 12'h999;
rom[89143] = 12'haaa;
rom[89144] = 12'hbbb;
rom[89145] = 12'hccc;
rom[89146] = 12'hddd;
rom[89147] = 12'heee;
rom[89148] = 12'hfff;
rom[89149] = 12'hfff;
rom[89150] = 12'heee;
rom[89151] = 12'hddd;
rom[89152] = 12'hbbb;
rom[89153] = 12'haaa;
rom[89154] = 12'h999;
rom[89155] = 12'h888;
rom[89156] = 12'h777;
rom[89157] = 12'h666;
rom[89158] = 12'h555;
rom[89159] = 12'h555;
rom[89160] = 12'h555;
rom[89161] = 12'h555;
rom[89162] = 12'h444;
rom[89163] = 12'h444;
rom[89164] = 12'h444;
rom[89165] = 12'h444;
rom[89166] = 12'h444;
rom[89167] = 12'h444;
rom[89168] = 12'h444;
rom[89169] = 12'h444;
rom[89170] = 12'h444;
rom[89171] = 12'h555;
rom[89172] = 12'h555;
rom[89173] = 12'h555;
rom[89174] = 12'h666;
rom[89175] = 12'h666;
rom[89176] = 12'h777;
rom[89177] = 12'h777;
rom[89178] = 12'h888;
rom[89179] = 12'h999;
rom[89180] = 12'h999;
rom[89181] = 12'h999;
rom[89182] = 12'h999;
rom[89183] = 12'h999;
rom[89184] = 12'h999;
rom[89185] = 12'h999;
rom[89186] = 12'h888;
rom[89187] = 12'h888;
rom[89188] = 12'h888;
rom[89189] = 12'h888;
rom[89190] = 12'h777;
rom[89191] = 12'h777;
rom[89192] = 12'h666;
rom[89193] = 12'h666;
rom[89194] = 12'h555;
rom[89195] = 12'h555;
rom[89196] = 12'h444;
rom[89197] = 12'h444;
rom[89198] = 12'h444;
rom[89199] = 12'h444;
rom[89200] = 12'hfff;
rom[89201] = 12'hfff;
rom[89202] = 12'hfff;
rom[89203] = 12'hfff;
rom[89204] = 12'hfff;
rom[89205] = 12'hfff;
rom[89206] = 12'hfff;
rom[89207] = 12'hfff;
rom[89208] = 12'hfff;
rom[89209] = 12'hfff;
rom[89210] = 12'hfff;
rom[89211] = 12'hfff;
rom[89212] = 12'hfff;
rom[89213] = 12'hfff;
rom[89214] = 12'hfff;
rom[89215] = 12'hfff;
rom[89216] = 12'hfff;
rom[89217] = 12'hfff;
rom[89218] = 12'hfff;
rom[89219] = 12'hfff;
rom[89220] = 12'hfff;
rom[89221] = 12'hfff;
rom[89222] = 12'hfff;
rom[89223] = 12'hfff;
rom[89224] = 12'hfff;
rom[89225] = 12'hfff;
rom[89226] = 12'hfff;
rom[89227] = 12'hfff;
rom[89228] = 12'hfff;
rom[89229] = 12'hfff;
rom[89230] = 12'hfff;
rom[89231] = 12'hfff;
rom[89232] = 12'hfff;
rom[89233] = 12'hfff;
rom[89234] = 12'hfff;
rom[89235] = 12'hfff;
rom[89236] = 12'hfff;
rom[89237] = 12'hfff;
rom[89238] = 12'hfff;
rom[89239] = 12'hfff;
rom[89240] = 12'hfff;
rom[89241] = 12'hfff;
rom[89242] = 12'hfff;
rom[89243] = 12'hfff;
rom[89244] = 12'hfff;
rom[89245] = 12'hfff;
rom[89246] = 12'hfff;
rom[89247] = 12'hfff;
rom[89248] = 12'hfff;
rom[89249] = 12'hfff;
rom[89250] = 12'hfff;
rom[89251] = 12'hfff;
rom[89252] = 12'hfff;
rom[89253] = 12'hfff;
rom[89254] = 12'hfff;
rom[89255] = 12'hfff;
rom[89256] = 12'hfff;
rom[89257] = 12'hfff;
rom[89258] = 12'hfff;
rom[89259] = 12'hfff;
rom[89260] = 12'hfff;
rom[89261] = 12'hfff;
rom[89262] = 12'hfff;
rom[89263] = 12'hfff;
rom[89264] = 12'hfff;
rom[89265] = 12'hfff;
rom[89266] = 12'hfff;
rom[89267] = 12'hfff;
rom[89268] = 12'hfff;
rom[89269] = 12'hfff;
rom[89270] = 12'hfff;
rom[89271] = 12'hfff;
rom[89272] = 12'hfff;
rom[89273] = 12'hfff;
rom[89274] = 12'hfff;
rom[89275] = 12'hfff;
rom[89276] = 12'hfff;
rom[89277] = 12'hfff;
rom[89278] = 12'hfff;
rom[89279] = 12'hfff;
rom[89280] = 12'hfff;
rom[89281] = 12'hfff;
rom[89282] = 12'hfff;
rom[89283] = 12'hfff;
rom[89284] = 12'hfff;
rom[89285] = 12'hfff;
rom[89286] = 12'hfff;
rom[89287] = 12'hfff;
rom[89288] = 12'hfff;
rom[89289] = 12'hfff;
rom[89290] = 12'hfff;
rom[89291] = 12'hfff;
rom[89292] = 12'hfff;
rom[89293] = 12'hfff;
rom[89294] = 12'hfff;
rom[89295] = 12'hfff;
rom[89296] = 12'hfff;
rom[89297] = 12'hfff;
rom[89298] = 12'hfff;
rom[89299] = 12'hfff;
rom[89300] = 12'hfff;
rom[89301] = 12'hfff;
rom[89302] = 12'hfff;
rom[89303] = 12'hfff;
rom[89304] = 12'hfff;
rom[89305] = 12'hfff;
rom[89306] = 12'hfff;
rom[89307] = 12'hfff;
rom[89308] = 12'hfff;
rom[89309] = 12'hfff;
rom[89310] = 12'hfff;
rom[89311] = 12'hfff;
rom[89312] = 12'hfff;
rom[89313] = 12'hfff;
rom[89314] = 12'hfff;
rom[89315] = 12'hfff;
rom[89316] = 12'hfff;
rom[89317] = 12'hfff;
rom[89318] = 12'hfff;
rom[89319] = 12'hfff;
rom[89320] = 12'hfff;
rom[89321] = 12'hfff;
rom[89322] = 12'hfff;
rom[89323] = 12'hfff;
rom[89324] = 12'hfff;
rom[89325] = 12'hfff;
rom[89326] = 12'hfff;
rom[89327] = 12'hfff;
rom[89328] = 12'heee;
rom[89329] = 12'heee;
rom[89330] = 12'heee;
rom[89331] = 12'hddd;
rom[89332] = 12'hddd;
rom[89333] = 12'hddd;
rom[89334] = 12'hddd;
rom[89335] = 12'hccc;
rom[89336] = 12'hccc;
rom[89337] = 12'hccc;
rom[89338] = 12'hbbb;
rom[89339] = 12'hbbb;
rom[89340] = 12'hbbb;
rom[89341] = 12'hbbb;
rom[89342] = 12'haaa;
rom[89343] = 12'haaa;
rom[89344] = 12'h999;
rom[89345] = 12'h999;
rom[89346] = 12'h999;
rom[89347] = 12'h999;
rom[89348] = 12'h888;
rom[89349] = 12'h888;
rom[89350] = 12'h888;
rom[89351] = 12'h888;
rom[89352] = 12'h888;
rom[89353] = 12'h888;
rom[89354] = 12'h888;
rom[89355] = 12'h888;
rom[89356] = 12'h888;
rom[89357] = 12'h888;
rom[89358] = 12'h777;
rom[89359] = 12'h777;
rom[89360] = 12'h777;
rom[89361] = 12'h777;
rom[89362] = 12'h777;
rom[89363] = 12'h777;
rom[89364] = 12'h777;
rom[89365] = 12'h777;
rom[89366] = 12'h888;
rom[89367] = 12'h888;
rom[89368] = 12'h888;
rom[89369] = 12'h888;
rom[89370] = 12'h888;
rom[89371] = 12'h888;
rom[89372] = 12'h888;
rom[89373] = 12'h888;
rom[89374] = 12'h777;
rom[89375] = 12'h777;
rom[89376] = 12'h777;
rom[89377] = 12'h777;
rom[89378] = 12'h666;
rom[89379] = 12'h666;
rom[89380] = 12'h666;
rom[89381] = 12'h666;
rom[89382] = 12'h666;
rom[89383] = 12'h666;
rom[89384] = 12'h666;
rom[89385] = 12'h666;
rom[89386] = 12'h666;
rom[89387] = 12'h666;
rom[89388] = 12'h666;
rom[89389] = 12'h666;
rom[89390] = 12'h666;
rom[89391] = 12'h666;
rom[89392] = 12'h666;
rom[89393] = 12'h666;
rom[89394] = 12'h666;
rom[89395] = 12'h666;
rom[89396] = 12'h666;
rom[89397] = 12'h666;
rom[89398] = 12'h666;
rom[89399] = 12'h666;
rom[89400] = 12'h555;
rom[89401] = 12'h555;
rom[89402] = 12'h555;
rom[89403] = 12'h555;
rom[89404] = 12'h555;
rom[89405] = 12'h555;
rom[89406] = 12'h555;
rom[89407] = 12'h555;
rom[89408] = 12'h555;
rom[89409] = 12'h444;
rom[89410] = 12'h444;
rom[89411] = 12'h444;
rom[89412] = 12'h444;
rom[89413] = 12'h444;
rom[89414] = 12'h444;
rom[89415] = 12'h333;
rom[89416] = 12'h333;
rom[89417] = 12'h333;
rom[89418] = 12'h333;
rom[89419] = 12'h333;
rom[89420] = 12'h444;
rom[89421] = 12'h666;
rom[89422] = 12'h666;
rom[89423] = 12'h777;
rom[89424] = 12'h888;
rom[89425] = 12'h777;
rom[89426] = 12'h555;
rom[89427] = 12'h444;
rom[89428] = 12'h444;
rom[89429] = 12'h444;
rom[89430] = 12'h333;
rom[89431] = 12'h333;
rom[89432] = 12'h333;
rom[89433] = 12'h222;
rom[89434] = 12'h222;
rom[89435] = 12'h111;
rom[89436] = 12'h111;
rom[89437] = 12'h111;
rom[89438] = 12'h111;
rom[89439] = 12'h111;
rom[89440] = 12'h111;
rom[89441] = 12'h111;
rom[89442] = 12'h111;
rom[89443] = 12'h111;
rom[89444] = 12'h111;
rom[89445] = 12'h  0;
rom[89446] = 12'h  0;
rom[89447] = 12'h  0;
rom[89448] = 12'h  0;
rom[89449] = 12'h  0;
rom[89450] = 12'h  0;
rom[89451] = 12'h  0;
rom[89452] = 12'h  0;
rom[89453] = 12'h  0;
rom[89454] = 12'h  0;
rom[89455] = 12'h  0;
rom[89456] = 12'h  0;
rom[89457] = 12'h  0;
rom[89458] = 12'h  0;
rom[89459] = 12'h  0;
rom[89460] = 12'h  0;
rom[89461] = 12'h  0;
rom[89462] = 12'h  0;
rom[89463] = 12'h111;
rom[89464] = 12'h111;
rom[89465] = 12'h111;
rom[89466] = 12'h111;
rom[89467] = 12'h111;
rom[89468] = 12'h111;
rom[89469] = 12'h111;
rom[89470] = 12'h111;
rom[89471] = 12'h111;
rom[89472] = 12'h111;
rom[89473] = 12'h222;
rom[89474] = 12'h222;
rom[89475] = 12'h333;
rom[89476] = 12'h333;
rom[89477] = 12'h333;
rom[89478] = 12'h555;
rom[89479] = 12'h666;
rom[89480] = 12'h777;
rom[89481] = 12'h888;
rom[89482] = 12'h888;
rom[89483] = 12'h888;
rom[89484] = 12'h888;
rom[89485] = 12'h777;
rom[89486] = 12'h777;
rom[89487] = 12'h777;
rom[89488] = 12'h777;
rom[89489] = 12'h777;
rom[89490] = 12'h777;
rom[89491] = 12'h777;
rom[89492] = 12'h777;
rom[89493] = 12'h888;
rom[89494] = 12'h888;
rom[89495] = 12'h999;
rom[89496] = 12'h888;
rom[89497] = 12'h888;
rom[89498] = 12'h888;
rom[89499] = 12'h999;
rom[89500] = 12'haaa;
rom[89501] = 12'hccc;
rom[89502] = 12'hccc;
rom[89503] = 12'hccc;
rom[89504] = 12'haaa;
rom[89505] = 12'h999;
rom[89506] = 12'h888;
rom[89507] = 12'h777;
rom[89508] = 12'h777;
rom[89509] = 12'h666;
rom[89510] = 12'h666;
rom[89511] = 12'h555;
rom[89512] = 12'h555;
rom[89513] = 12'h555;
rom[89514] = 12'h444;
rom[89515] = 12'h444;
rom[89516] = 12'h444;
rom[89517] = 12'h444;
rom[89518] = 12'h444;
rom[89519] = 12'h444;
rom[89520] = 12'h444;
rom[89521] = 12'h444;
rom[89522] = 12'h444;
rom[89523] = 12'h444;
rom[89524] = 12'h444;
rom[89525] = 12'h444;
rom[89526] = 12'h555;
rom[89527] = 12'h555;
rom[89528] = 12'h444;
rom[89529] = 12'h444;
rom[89530] = 12'h444;
rom[89531] = 12'h444;
rom[89532] = 12'h444;
rom[89533] = 12'h444;
rom[89534] = 12'h444;
rom[89535] = 12'h444;
rom[89536] = 12'h444;
rom[89537] = 12'h444;
rom[89538] = 12'h555;
rom[89539] = 12'h555;
rom[89540] = 12'h555;
rom[89541] = 12'h666;
rom[89542] = 12'h777;
rom[89543] = 12'h777;
rom[89544] = 12'h888;
rom[89545] = 12'h999;
rom[89546] = 12'hbbb;
rom[89547] = 12'hccc;
rom[89548] = 12'heee;
rom[89549] = 12'hfff;
rom[89550] = 12'hfff;
rom[89551] = 12'hfff;
rom[89552] = 12'hddd;
rom[89553] = 12'hccc;
rom[89554] = 12'hbbb;
rom[89555] = 12'h999;
rom[89556] = 12'h888;
rom[89557] = 12'h777;
rom[89558] = 12'h777;
rom[89559] = 12'h666;
rom[89560] = 12'h666;
rom[89561] = 12'h666;
rom[89562] = 12'h555;
rom[89563] = 12'h555;
rom[89564] = 12'h555;
rom[89565] = 12'h444;
rom[89566] = 12'h444;
rom[89567] = 12'h444;
rom[89568] = 12'h444;
rom[89569] = 12'h444;
rom[89570] = 12'h444;
rom[89571] = 12'h444;
rom[89572] = 12'h333;
rom[89573] = 12'h333;
rom[89574] = 12'h444;
rom[89575] = 12'h444;
rom[89576] = 12'h444;
rom[89577] = 12'h555;
rom[89578] = 12'h555;
rom[89579] = 12'h666;
rom[89580] = 12'h666;
rom[89581] = 12'h777;
rom[89582] = 12'h888;
rom[89583] = 12'h888;
rom[89584] = 12'h999;
rom[89585] = 12'h999;
rom[89586] = 12'h999;
rom[89587] = 12'h999;
rom[89588] = 12'h999;
rom[89589] = 12'h999;
rom[89590] = 12'h999;
rom[89591] = 12'h999;
rom[89592] = 12'h888;
rom[89593] = 12'h888;
rom[89594] = 12'h888;
rom[89595] = 12'h777;
rom[89596] = 12'h777;
rom[89597] = 12'h666;
rom[89598] = 12'h666;
rom[89599] = 12'h666;
rom[89600] = 12'hfff;
rom[89601] = 12'hfff;
rom[89602] = 12'hfff;
rom[89603] = 12'hfff;
rom[89604] = 12'hfff;
rom[89605] = 12'hfff;
rom[89606] = 12'hfff;
rom[89607] = 12'hfff;
rom[89608] = 12'hfff;
rom[89609] = 12'hfff;
rom[89610] = 12'hfff;
rom[89611] = 12'hfff;
rom[89612] = 12'hfff;
rom[89613] = 12'hfff;
rom[89614] = 12'hfff;
rom[89615] = 12'hfff;
rom[89616] = 12'hfff;
rom[89617] = 12'hfff;
rom[89618] = 12'hfff;
rom[89619] = 12'hfff;
rom[89620] = 12'hfff;
rom[89621] = 12'hfff;
rom[89622] = 12'hfff;
rom[89623] = 12'hfff;
rom[89624] = 12'hfff;
rom[89625] = 12'hfff;
rom[89626] = 12'hfff;
rom[89627] = 12'hfff;
rom[89628] = 12'hfff;
rom[89629] = 12'hfff;
rom[89630] = 12'hfff;
rom[89631] = 12'hfff;
rom[89632] = 12'hfff;
rom[89633] = 12'hfff;
rom[89634] = 12'hfff;
rom[89635] = 12'hfff;
rom[89636] = 12'hfff;
rom[89637] = 12'hfff;
rom[89638] = 12'hfff;
rom[89639] = 12'hfff;
rom[89640] = 12'hfff;
rom[89641] = 12'hfff;
rom[89642] = 12'hfff;
rom[89643] = 12'hfff;
rom[89644] = 12'hfff;
rom[89645] = 12'hfff;
rom[89646] = 12'hfff;
rom[89647] = 12'hfff;
rom[89648] = 12'hfff;
rom[89649] = 12'hfff;
rom[89650] = 12'hfff;
rom[89651] = 12'hfff;
rom[89652] = 12'hfff;
rom[89653] = 12'hfff;
rom[89654] = 12'hfff;
rom[89655] = 12'hfff;
rom[89656] = 12'hfff;
rom[89657] = 12'hfff;
rom[89658] = 12'hfff;
rom[89659] = 12'hfff;
rom[89660] = 12'hfff;
rom[89661] = 12'hfff;
rom[89662] = 12'hfff;
rom[89663] = 12'hfff;
rom[89664] = 12'hfff;
rom[89665] = 12'hfff;
rom[89666] = 12'hfff;
rom[89667] = 12'hfff;
rom[89668] = 12'hfff;
rom[89669] = 12'hfff;
rom[89670] = 12'hfff;
rom[89671] = 12'hfff;
rom[89672] = 12'hfff;
rom[89673] = 12'hfff;
rom[89674] = 12'hfff;
rom[89675] = 12'hfff;
rom[89676] = 12'hfff;
rom[89677] = 12'hfff;
rom[89678] = 12'hfff;
rom[89679] = 12'hfff;
rom[89680] = 12'hfff;
rom[89681] = 12'hfff;
rom[89682] = 12'hfff;
rom[89683] = 12'hfff;
rom[89684] = 12'hfff;
rom[89685] = 12'hfff;
rom[89686] = 12'hfff;
rom[89687] = 12'hfff;
rom[89688] = 12'hfff;
rom[89689] = 12'hfff;
rom[89690] = 12'hfff;
rom[89691] = 12'hfff;
rom[89692] = 12'hfff;
rom[89693] = 12'hfff;
rom[89694] = 12'hfff;
rom[89695] = 12'hfff;
rom[89696] = 12'hfff;
rom[89697] = 12'hfff;
rom[89698] = 12'hfff;
rom[89699] = 12'hfff;
rom[89700] = 12'hfff;
rom[89701] = 12'hfff;
rom[89702] = 12'hfff;
rom[89703] = 12'hfff;
rom[89704] = 12'hfff;
rom[89705] = 12'hfff;
rom[89706] = 12'hfff;
rom[89707] = 12'hfff;
rom[89708] = 12'hfff;
rom[89709] = 12'hfff;
rom[89710] = 12'hfff;
rom[89711] = 12'hfff;
rom[89712] = 12'hfff;
rom[89713] = 12'hfff;
rom[89714] = 12'hfff;
rom[89715] = 12'hfff;
rom[89716] = 12'hfff;
rom[89717] = 12'hfff;
rom[89718] = 12'hfff;
rom[89719] = 12'hfff;
rom[89720] = 12'hfff;
rom[89721] = 12'hfff;
rom[89722] = 12'hfff;
rom[89723] = 12'hfff;
rom[89724] = 12'hfff;
rom[89725] = 12'hfff;
rom[89726] = 12'hfff;
rom[89727] = 12'hfff;
rom[89728] = 12'hfff;
rom[89729] = 12'hfff;
rom[89730] = 12'heee;
rom[89731] = 12'heee;
rom[89732] = 12'heee;
rom[89733] = 12'hddd;
rom[89734] = 12'hddd;
rom[89735] = 12'hddd;
rom[89736] = 12'hccc;
rom[89737] = 12'hccc;
rom[89738] = 12'hccc;
rom[89739] = 12'hbbb;
rom[89740] = 12'hbbb;
rom[89741] = 12'hbbb;
rom[89742] = 12'haaa;
rom[89743] = 12'haaa;
rom[89744] = 12'haaa;
rom[89745] = 12'h999;
rom[89746] = 12'h999;
rom[89747] = 12'h888;
rom[89748] = 12'h888;
rom[89749] = 12'h999;
rom[89750] = 12'h999;
rom[89751] = 12'h999;
rom[89752] = 12'h888;
rom[89753] = 12'h888;
rom[89754] = 12'h888;
rom[89755] = 12'h888;
rom[89756] = 12'h888;
rom[89757] = 12'h777;
rom[89758] = 12'h777;
rom[89759] = 12'h777;
rom[89760] = 12'h777;
rom[89761] = 12'h777;
rom[89762] = 12'h777;
rom[89763] = 12'h777;
rom[89764] = 12'h777;
rom[89765] = 12'h777;
rom[89766] = 12'h777;
rom[89767] = 12'h777;
rom[89768] = 12'h888;
rom[89769] = 12'h888;
rom[89770] = 12'h888;
rom[89771] = 12'h888;
rom[89772] = 12'h888;
rom[89773] = 12'h888;
rom[89774] = 12'h888;
rom[89775] = 12'h888;
rom[89776] = 12'h777;
rom[89777] = 12'h777;
rom[89778] = 12'h777;
rom[89779] = 12'h777;
rom[89780] = 12'h777;
rom[89781] = 12'h777;
rom[89782] = 12'h666;
rom[89783] = 12'h666;
rom[89784] = 12'h666;
rom[89785] = 12'h666;
rom[89786] = 12'h666;
rom[89787] = 12'h666;
rom[89788] = 12'h666;
rom[89789] = 12'h666;
rom[89790] = 12'h666;
rom[89791] = 12'h666;
rom[89792] = 12'h666;
rom[89793] = 12'h666;
rom[89794] = 12'h666;
rom[89795] = 12'h666;
rom[89796] = 12'h666;
rom[89797] = 12'h666;
rom[89798] = 12'h666;
rom[89799] = 12'h666;
rom[89800] = 12'h666;
rom[89801] = 12'h555;
rom[89802] = 12'h555;
rom[89803] = 12'h555;
rom[89804] = 12'h555;
rom[89805] = 12'h555;
rom[89806] = 12'h555;
rom[89807] = 12'h555;
rom[89808] = 12'h555;
rom[89809] = 12'h444;
rom[89810] = 12'h444;
rom[89811] = 12'h444;
rom[89812] = 12'h444;
rom[89813] = 12'h444;
rom[89814] = 12'h333;
rom[89815] = 12'h333;
rom[89816] = 12'h333;
rom[89817] = 12'h333;
rom[89818] = 12'h222;
rom[89819] = 12'h222;
rom[89820] = 12'h222;
rom[89821] = 12'h333;
rom[89822] = 12'h444;
rom[89823] = 12'h555;
rom[89824] = 12'h777;
rom[89825] = 12'h777;
rom[89826] = 12'h777;
rom[89827] = 12'h666;
rom[89828] = 12'h555;
rom[89829] = 12'h444;
rom[89830] = 12'h444;
rom[89831] = 12'h444;
rom[89832] = 12'h333;
rom[89833] = 12'h333;
rom[89834] = 12'h333;
rom[89835] = 12'h222;
rom[89836] = 12'h222;
rom[89837] = 12'h111;
rom[89838] = 12'h111;
rom[89839] = 12'h111;
rom[89840] = 12'h111;
rom[89841] = 12'h111;
rom[89842] = 12'h111;
rom[89843] = 12'h111;
rom[89844] = 12'h  0;
rom[89845] = 12'h  0;
rom[89846] = 12'h  0;
rom[89847] = 12'h  0;
rom[89848] = 12'h  0;
rom[89849] = 12'h  0;
rom[89850] = 12'h  0;
rom[89851] = 12'h  0;
rom[89852] = 12'h  0;
rom[89853] = 12'h  0;
rom[89854] = 12'h  0;
rom[89855] = 12'h  0;
rom[89856] = 12'h  0;
rom[89857] = 12'h  0;
rom[89858] = 12'h  0;
rom[89859] = 12'h  0;
rom[89860] = 12'h  0;
rom[89861] = 12'h  0;
rom[89862] = 12'h  0;
rom[89863] = 12'h111;
rom[89864] = 12'h111;
rom[89865] = 12'h111;
rom[89866] = 12'h111;
rom[89867] = 12'h111;
rom[89868] = 12'h111;
rom[89869] = 12'h111;
rom[89870] = 12'h111;
rom[89871] = 12'h222;
rom[89872] = 12'h222;
rom[89873] = 12'h222;
rom[89874] = 12'h222;
rom[89875] = 12'h333;
rom[89876] = 12'h333;
rom[89877] = 12'h444;
rom[89878] = 12'h555;
rom[89879] = 12'h666;
rom[89880] = 12'h888;
rom[89881] = 12'h888;
rom[89882] = 12'h888;
rom[89883] = 12'h888;
rom[89884] = 12'h888;
rom[89885] = 12'h777;
rom[89886] = 12'h777;
rom[89887] = 12'h777;
rom[89888] = 12'h777;
rom[89889] = 12'h777;
rom[89890] = 12'h777;
rom[89891] = 12'h888;
rom[89892] = 12'h888;
rom[89893] = 12'h888;
rom[89894] = 12'h888;
rom[89895] = 12'h999;
rom[89896] = 12'h999;
rom[89897] = 12'h888;
rom[89898] = 12'h888;
rom[89899] = 12'haaa;
rom[89900] = 12'hbbb;
rom[89901] = 12'hccc;
rom[89902] = 12'hccc;
rom[89903] = 12'hbbb;
rom[89904] = 12'haaa;
rom[89905] = 12'h999;
rom[89906] = 12'h888;
rom[89907] = 12'h777;
rom[89908] = 12'h777;
rom[89909] = 12'h666;
rom[89910] = 12'h666;
rom[89911] = 12'h555;
rom[89912] = 12'h555;
rom[89913] = 12'h555;
rom[89914] = 12'h444;
rom[89915] = 12'h444;
rom[89916] = 12'h444;
rom[89917] = 12'h444;
rom[89918] = 12'h444;
rom[89919] = 12'h444;
rom[89920] = 12'h444;
rom[89921] = 12'h444;
rom[89922] = 12'h444;
rom[89923] = 12'h444;
rom[89924] = 12'h444;
rom[89925] = 12'h444;
rom[89926] = 12'h444;
rom[89927] = 12'h444;
rom[89928] = 12'h444;
rom[89929] = 12'h444;
rom[89930] = 12'h444;
rom[89931] = 12'h444;
rom[89932] = 12'h444;
rom[89933] = 12'h444;
rom[89934] = 12'h444;
rom[89935] = 12'h444;
rom[89936] = 12'h444;
rom[89937] = 12'h444;
rom[89938] = 12'h444;
rom[89939] = 12'h444;
rom[89940] = 12'h444;
rom[89941] = 12'h444;
rom[89942] = 12'h444;
rom[89943] = 12'h444;
rom[89944] = 12'h555;
rom[89945] = 12'h666;
rom[89946] = 12'h777;
rom[89947] = 12'h888;
rom[89948] = 12'haaa;
rom[89949] = 12'hbbb;
rom[89950] = 12'hddd;
rom[89951] = 12'hfff;
rom[89952] = 12'hfff;
rom[89953] = 12'hfff;
rom[89954] = 12'hfff;
rom[89955] = 12'hddd;
rom[89956] = 12'hbbb;
rom[89957] = 12'h999;
rom[89958] = 12'h888;
rom[89959] = 12'h777;
rom[89960] = 12'h666;
rom[89961] = 12'h666;
rom[89962] = 12'h666;
rom[89963] = 12'h666;
rom[89964] = 12'h555;
rom[89965] = 12'h555;
rom[89966] = 12'h444;
rom[89967] = 12'h555;
rom[89968] = 12'h444;
rom[89969] = 12'h333;
rom[89970] = 12'h333;
rom[89971] = 12'h333;
rom[89972] = 12'h444;
rom[89973] = 12'h444;
rom[89974] = 12'h333;
rom[89975] = 12'h333;
rom[89976] = 12'h333;
rom[89977] = 12'h333;
rom[89978] = 12'h333;
rom[89979] = 12'h333;
rom[89980] = 12'h444;
rom[89981] = 12'h444;
rom[89982] = 12'h444;
rom[89983] = 12'h555;
rom[89984] = 12'h555;
rom[89985] = 12'h666;
rom[89986] = 12'h666;
rom[89987] = 12'h777;
rom[89988] = 12'h777;
rom[89989] = 12'h888;
rom[89990] = 12'h888;
rom[89991] = 12'h888;
rom[89992] = 12'h999;
rom[89993] = 12'h999;
rom[89994] = 12'h999;
rom[89995] = 12'h999;
rom[89996] = 12'h888;
rom[89997] = 12'h888;
rom[89998] = 12'h888;
rom[89999] = 12'h888;
rom[90000] = 12'hfff;
rom[90001] = 12'hfff;
rom[90002] = 12'hfff;
rom[90003] = 12'hfff;
rom[90004] = 12'hfff;
rom[90005] = 12'hfff;
rom[90006] = 12'hfff;
rom[90007] = 12'hfff;
rom[90008] = 12'hfff;
rom[90009] = 12'hfff;
rom[90010] = 12'hfff;
rom[90011] = 12'hfff;
rom[90012] = 12'hfff;
rom[90013] = 12'hfff;
rom[90014] = 12'hfff;
rom[90015] = 12'hfff;
rom[90016] = 12'hfff;
rom[90017] = 12'hfff;
rom[90018] = 12'hfff;
rom[90019] = 12'hfff;
rom[90020] = 12'hfff;
rom[90021] = 12'hfff;
rom[90022] = 12'hfff;
rom[90023] = 12'hfff;
rom[90024] = 12'hfff;
rom[90025] = 12'hfff;
rom[90026] = 12'hfff;
rom[90027] = 12'hfff;
rom[90028] = 12'hfff;
rom[90029] = 12'hfff;
rom[90030] = 12'hfff;
rom[90031] = 12'hfff;
rom[90032] = 12'hfff;
rom[90033] = 12'hfff;
rom[90034] = 12'hfff;
rom[90035] = 12'hfff;
rom[90036] = 12'hfff;
rom[90037] = 12'hfff;
rom[90038] = 12'hfff;
rom[90039] = 12'hfff;
rom[90040] = 12'hfff;
rom[90041] = 12'hfff;
rom[90042] = 12'hfff;
rom[90043] = 12'hfff;
rom[90044] = 12'hfff;
rom[90045] = 12'hfff;
rom[90046] = 12'hfff;
rom[90047] = 12'hfff;
rom[90048] = 12'hfff;
rom[90049] = 12'hfff;
rom[90050] = 12'hfff;
rom[90051] = 12'hfff;
rom[90052] = 12'hfff;
rom[90053] = 12'hfff;
rom[90054] = 12'hfff;
rom[90055] = 12'hfff;
rom[90056] = 12'hfff;
rom[90057] = 12'hfff;
rom[90058] = 12'hfff;
rom[90059] = 12'hfff;
rom[90060] = 12'hfff;
rom[90061] = 12'hfff;
rom[90062] = 12'hfff;
rom[90063] = 12'hfff;
rom[90064] = 12'hfff;
rom[90065] = 12'hfff;
rom[90066] = 12'hfff;
rom[90067] = 12'hfff;
rom[90068] = 12'hfff;
rom[90069] = 12'hfff;
rom[90070] = 12'hfff;
rom[90071] = 12'hfff;
rom[90072] = 12'hfff;
rom[90073] = 12'hfff;
rom[90074] = 12'hfff;
rom[90075] = 12'hfff;
rom[90076] = 12'hfff;
rom[90077] = 12'hfff;
rom[90078] = 12'hfff;
rom[90079] = 12'hfff;
rom[90080] = 12'hfff;
rom[90081] = 12'hfff;
rom[90082] = 12'hfff;
rom[90083] = 12'hfff;
rom[90084] = 12'hfff;
rom[90085] = 12'hfff;
rom[90086] = 12'hfff;
rom[90087] = 12'hfff;
rom[90088] = 12'hfff;
rom[90089] = 12'hfff;
rom[90090] = 12'hfff;
rom[90091] = 12'hfff;
rom[90092] = 12'hfff;
rom[90093] = 12'hfff;
rom[90094] = 12'hfff;
rom[90095] = 12'hfff;
rom[90096] = 12'hfff;
rom[90097] = 12'hfff;
rom[90098] = 12'hfff;
rom[90099] = 12'hfff;
rom[90100] = 12'hfff;
rom[90101] = 12'hfff;
rom[90102] = 12'hfff;
rom[90103] = 12'hfff;
rom[90104] = 12'hfff;
rom[90105] = 12'hfff;
rom[90106] = 12'hfff;
rom[90107] = 12'hfff;
rom[90108] = 12'hfff;
rom[90109] = 12'hfff;
rom[90110] = 12'hfff;
rom[90111] = 12'hfff;
rom[90112] = 12'hfff;
rom[90113] = 12'hfff;
rom[90114] = 12'hfff;
rom[90115] = 12'hfff;
rom[90116] = 12'hfff;
rom[90117] = 12'hfff;
rom[90118] = 12'hfff;
rom[90119] = 12'hfff;
rom[90120] = 12'hfff;
rom[90121] = 12'hfff;
rom[90122] = 12'hfff;
rom[90123] = 12'hfff;
rom[90124] = 12'hfff;
rom[90125] = 12'hfff;
rom[90126] = 12'hfff;
rom[90127] = 12'hfff;
rom[90128] = 12'hfff;
rom[90129] = 12'hfff;
rom[90130] = 12'hfff;
rom[90131] = 12'heee;
rom[90132] = 12'heee;
rom[90133] = 12'heee;
rom[90134] = 12'hddd;
rom[90135] = 12'hddd;
rom[90136] = 12'hccc;
rom[90137] = 12'hccc;
rom[90138] = 12'hccc;
rom[90139] = 12'hbbb;
rom[90140] = 12'hbbb;
rom[90141] = 12'hbbb;
rom[90142] = 12'haaa;
rom[90143] = 12'haaa;
rom[90144] = 12'haaa;
rom[90145] = 12'haaa;
rom[90146] = 12'h999;
rom[90147] = 12'h999;
rom[90148] = 12'h999;
rom[90149] = 12'h999;
rom[90150] = 12'h999;
rom[90151] = 12'h999;
rom[90152] = 12'h888;
rom[90153] = 12'h888;
rom[90154] = 12'h888;
rom[90155] = 12'h888;
rom[90156] = 12'h888;
rom[90157] = 12'h777;
rom[90158] = 12'h777;
rom[90159] = 12'h777;
rom[90160] = 12'h777;
rom[90161] = 12'h777;
rom[90162] = 12'h777;
rom[90163] = 12'h777;
rom[90164] = 12'h777;
rom[90165] = 12'h777;
rom[90166] = 12'h777;
rom[90167] = 12'h777;
rom[90168] = 12'h888;
rom[90169] = 12'h888;
rom[90170] = 12'h888;
rom[90171] = 12'h888;
rom[90172] = 12'h888;
rom[90173] = 12'h888;
rom[90174] = 12'h888;
rom[90175] = 12'h888;
rom[90176] = 12'h777;
rom[90177] = 12'h777;
rom[90178] = 12'h777;
rom[90179] = 12'h777;
rom[90180] = 12'h777;
rom[90181] = 12'h777;
rom[90182] = 12'h777;
rom[90183] = 12'h777;
rom[90184] = 12'h666;
rom[90185] = 12'h666;
rom[90186] = 12'h666;
rom[90187] = 12'h666;
rom[90188] = 12'h666;
rom[90189] = 12'h666;
rom[90190] = 12'h666;
rom[90191] = 12'h666;
rom[90192] = 12'h666;
rom[90193] = 12'h666;
rom[90194] = 12'h666;
rom[90195] = 12'h666;
rom[90196] = 12'h666;
rom[90197] = 12'h666;
rom[90198] = 12'h666;
rom[90199] = 12'h666;
rom[90200] = 12'h666;
rom[90201] = 12'h666;
rom[90202] = 12'h555;
rom[90203] = 12'h555;
rom[90204] = 12'h555;
rom[90205] = 12'h555;
rom[90206] = 12'h555;
rom[90207] = 12'h555;
rom[90208] = 12'h555;
rom[90209] = 12'h444;
rom[90210] = 12'h444;
rom[90211] = 12'h444;
rom[90212] = 12'h444;
rom[90213] = 12'h444;
rom[90214] = 12'h333;
rom[90215] = 12'h333;
rom[90216] = 12'h333;
rom[90217] = 12'h222;
rom[90218] = 12'h222;
rom[90219] = 12'h222;
rom[90220] = 12'h222;
rom[90221] = 12'h222;
rom[90222] = 12'h333;
rom[90223] = 12'h444;
rom[90224] = 12'h555;
rom[90225] = 12'h666;
rom[90226] = 12'h777;
rom[90227] = 12'h777;
rom[90228] = 12'h666;
rom[90229] = 12'h555;
rom[90230] = 12'h444;
rom[90231] = 12'h444;
rom[90232] = 12'h444;
rom[90233] = 12'h333;
rom[90234] = 12'h333;
rom[90235] = 12'h222;
rom[90236] = 12'h222;
rom[90237] = 12'h222;
rom[90238] = 12'h111;
rom[90239] = 12'h111;
rom[90240] = 12'h111;
rom[90241] = 12'h111;
rom[90242] = 12'h111;
rom[90243] = 12'h111;
rom[90244] = 12'h111;
rom[90245] = 12'h  0;
rom[90246] = 12'h  0;
rom[90247] = 12'h  0;
rom[90248] = 12'h  0;
rom[90249] = 12'h  0;
rom[90250] = 12'h  0;
rom[90251] = 12'h  0;
rom[90252] = 12'h  0;
rom[90253] = 12'h  0;
rom[90254] = 12'h  0;
rom[90255] = 12'h  0;
rom[90256] = 12'h  0;
rom[90257] = 12'h  0;
rom[90258] = 12'h  0;
rom[90259] = 12'h  0;
rom[90260] = 12'h  0;
rom[90261] = 12'h  0;
rom[90262] = 12'h  0;
rom[90263] = 12'h111;
rom[90264] = 12'h111;
rom[90265] = 12'h111;
rom[90266] = 12'h111;
rom[90267] = 12'h111;
rom[90268] = 12'h111;
rom[90269] = 12'h111;
rom[90270] = 12'h111;
rom[90271] = 12'h222;
rom[90272] = 12'h222;
rom[90273] = 12'h222;
rom[90274] = 12'h333;
rom[90275] = 12'h333;
rom[90276] = 12'h444;
rom[90277] = 12'h555;
rom[90278] = 12'h666;
rom[90279] = 12'h777;
rom[90280] = 12'h888;
rom[90281] = 12'h888;
rom[90282] = 12'h888;
rom[90283] = 12'h888;
rom[90284] = 12'h777;
rom[90285] = 12'h777;
rom[90286] = 12'h777;
rom[90287] = 12'h777;
rom[90288] = 12'h777;
rom[90289] = 12'h777;
rom[90290] = 12'h777;
rom[90291] = 12'h888;
rom[90292] = 12'h888;
rom[90293] = 12'h888;
rom[90294] = 12'h999;
rom[90295] = 12'h999;
rom[90296] = 12'h999;
rom[90297] = 12'h999;
rom[90298] = 12'h999;
rom[90299] = 12'hbbb;
rom[90300] = 12'hccc;
rom[90301] = 12'hddd;
rom[90302] = 12'hccc;
rom[90303] = 12'hbbb;
rom[90304] = 12'h999;
rom[90305] = 12'h888;
rom[90306] = 12'h777;
rom[90307] = 12'h777;
rom[90308] = 12'h777;
rom[90309] = 12'h666;
rom[90310] = 12'h555;
rom[90311] = 12'h555;
rom[90312] = 12'h555;
rom[90313] = 12'h555;
rom[90314] = 12'h444;
rom[90315] = 12'h444;
rom[90316] = 12'h444;
rom[90317] = 12'h444;
rom[90318] = 12'h444;
rom[90319] = 12'h444;
rom[90320] = 12'h444;
rom[90321] = 12'h444;
rom[90322] = 12'h444;
rom[90323] = 12'h444;
rom[90324] = 12'h444;
rom[90325] = 12'h444;
rom[90326] = 12'h444;
rom[90327] = 12'h444;
rom[90328] = 12'h333;
rom[90329] = 12'h444;
rom[90330] = 12'h444;
rom[90331] = 12'h444;
rom[90332] = 12'h444;
rom[90333] = 12'h444;
rom[90334] = 12'h444;
rom[90335] = 12'h444;
rom[90336] = 12'h444;
rom[90337] = 12'h444;
rom[90338] = 12'h444;
rom[90339] = 12'h444;
rom[90340] = 12'h444;
rom[90341] = 12'h444;
rom[90342] = 12'h333;
rom[90343] = 12'h333;
rom[90344] = 12'h333;
rom[90345] = 12'h444;
rom[90346] = 12'h555;
rom[90347] = 12'h555;
rom[90348] = 12'h666;
rom[90349] = 12'h888;
rom[90350] = 12'h999;
rom[90351] = 12'hbbb;
rom[90352] = 12'hddd;
rom[90353] = 12'heee;
rom[90354] = 12'heee;
rom[90355] = 12'heee;
rom[90356] = 12'heee;
rom[90357] = 12'hccc;
rom[90358] = 12'haaa;
rom[90359] = 12'h888;
rom[90360] = 12'h777;
rom[90361] = 12'h666;
rom[90362] = 12'h666;
rom[90363] = 12'h666;
rom[90364] = 12'h555;
rom[90365] = 12'h555;
rom[90366] = 12'h444;
rom[90367] = 12'h444;
rom[90368] = 12'h555;
rom[90369] = 12'h444;
rom[90370] = 12'h444;
rom[90371] = 12'h444;
rom[90372] = 12'h444;
rom[90373] = 12'h444;
rom[90374] = 12'h333;
rom[90375] = 12'h333;
rom[90376] = 12'h333;
rom[90377] = 12'h333;
rom[90378] = 12'h333;
rom[90379] = 12'h333;
rom[90380] = 12'h333;
rom[90381] = 12'h333;
rom[90382] = 12'h333;
rom[90383] = 12'h333;
rom[90384] = 12'h333;
rom[90385] = 12'h444;
rom[90386] = 12'h444;
rom[90387] = 12'h444;
rom[90388] = 12'h555;
rom[90389] = 12'h555;
rom[90390] = 12'h666;
rom[90391] = 12'h666;
rom[90392] = 12'h777;
rom[90393] = 12'h777;
rom[90394] = 12'h777;
rom[90395] = 12'h777;
rom[90396] = 12'h888;
rom[90397] = 12'h888;
rom[90398] = 12'h888;
rom[90399] = 12'h888;
rom[90400] = 12'hfff;
rom[90401] = 12'hfff;
rom[90402] = 12'hfff;
rom[90403] = 12'hfff;
rom[90404] = 12'hfff;
rom[90405] = 12'hfff;
rom[90406] = 12'hfff;
rom[90407] = 12'hfff;
rom[90408] = 12'hfff;
rom[90409] = 12'hfff;
rom[90410] = 12'hfff;
rom[90411] = 12'hfff;
rom[90412] = 12'hfff;
rom[90413] = 12'hfff;
rom[90414] = 12'hfff;
rom[90415] = 12'hfff;
rom[90416] = 12'hfff;
rom[90417] = 12'hfff;
rom[90418] = 12'hfff;
rom[90419] = 12'hfff;
rom[90420] = 12'hfff;
rom[90421] = 12'hfff;
rom[90422] = 12'hfff;
rom[90423] = 12'hfff;
rom[90424] = 12'hfff;
rom[90425] = 12'hfff;
rom[90426] = 12'hfff;
rom[90427] = 12'hfff;
rom[90428] = 12'hfff;
rom[90429] = 12'hfff;
rom[90430] = 12'hfff;
rom[90431] = 12'hfff;
rom[90432] = 12'hfff;
rom[90433] = 12'hfff;
rom[90434] = 12'hfff;
rom[90435] = 12'hfff;
rom[90436] = 12'hfff;
rom[90437] = 12'hfff;
rom[90438] = 12'hfff;
rom[90439] = 12'hfff;
rom[90440] = 12'hfff;
rom[90441] = 12'hfff;
rom[90442] = 12'hfff;
rom[90443] = 12'hfff;
rom[90444] = 12'hfff;
rom[90445] = 12'hfff;
rom[90446] = 12'hfff;
rom[90447] = 12'hfff;
rom[90448] = 12'hfff;
rom[90449] = 12'hfff;
rom[90450] = 12'hfff;
rom[90451] = 12'hfff;
rom[90452] = 12'hfff;
rom[90453] = 12'hfff;
rom[90454] = 12'hfff;
rom[90455] = 12'hfff;
rom[90456] = 12'hfff;
rom[90457] = 12'hfff;
rom[90458] = 12'hfff;
rom[90459] = 12'hfff;
rom[90460] = 12'hfff;
rom[90461] = 12'hfff;
rom[90462] = 12'hfff;
rom[90463] = 12'hfff;
rom[90464] = 12'hfff;
rom[90465] = 12'hfff;
rom[90466] = 12'hfff;
rom[90467] = 12'hfff;
rom[90468] = 12'hfff;
rom[90469] = 12'hfff;
rom[90470] = 12'hfff;
rom[90471] = 12'hfff;
rom[90472] = 12'hfff;
rom[90473] = 12'hfff;
rom[90474] = 12'hfff;
rom[90475] = 12'hfff;
rom[90476] = 12'hfff;
rom[90477] = 12'hfff;
rom[90478] = 12'hfff;
rom[90479] = 12'hfff;
rom[90480] = 12'hfff;
rom[90481] = 12'hfff;
rom[90482] = 12'hfff;
rom[90483] = 12'hfff;
rom[90484] = 12'hfff;
rom[90485] = 12'hfff;
rom[90486] = 12'hfff;
rom[90487] = 12'hfff;
rom[90488] = 12'hfff;
rom[90489] = 12'hfff;
rom[90490] = 12'hfff;
rom[90491] = 12'hfff;
rom[90492] = 12'hfff;
rom[90493] = 12'hfff;
rom[90494] = 12'hfff;
rom[90495] = 12'hfff;
rom[90496] = 12'hfff;
rom[90497] = 12'hfff;
rom[90498] = 12'hfff;
rom[90499] = 12'hfff;
rom[90500] = 12'hfff;
rom[90501] = 12'hfff;
rom[90502] = 12'hfff;
rom[90503] = 12'hfff;
rom[90504] = 12'hfff;
rom[90505] = 12'hfff;
rom[90506] = 12'hfff;
rom[90507] = 12'hfff;
rom[90508] = 12'hfff;
rom[90509] = 12'hfff;
rom[90510] = 12'hfff;
rom[90511] = 12'hfff;
rom[90512] = 12'hfff;
rom[90513] = 12'hfff;
rom[90514] = 12'hfff;
rom[90515] = 12'hfff;
rom[90516] = 12'hfff;
rom[90517] = 12'hfff;
rom[90518] = 12'hfff;
rom[90519] = 12'hfff;
rom[90520] = 12'hfff;
rom[90521] = 12'hfff;
rom[90522] = 12'hfff;
rom[90523] = 12'hfff;
rom[90524] = 12'hfff;
rom[90525] = 12'hfff;
rom[90526] = 12'hfff;
rom[90527] = 12'hfff;
rom[90528] = 12'hfff;
rom[90529] = 12'hfff;
rom[90530] = 12'hfff;
rom[90531] = 12'hfff;
rom[90532] = 12'hfff;
rom[90533] = 12'heee;
rom[90534] = 12'heee;
rom[90535] = 12'heee;
rom[90536] = 12'hddd;
rom[90537] = 12'hddd;
rom[90538] = 12'hccc;
rom[90539] = 12'hccc;
rom[90540] = 12'hccc;
rom[90541] = 12'hbbb;
rom[90542] = 12'hbbb;
rom[90543] = 12'haaa;
rom[90544] = 12'haaa;
rom[90545] = 12'haaa;
rom[90546] = 12'h999;
rom[90547] = 12'h999;
rom[90548] = 12'h999;
rom[90549] = 12'h999;
rom[90550] = 12'h999;
rom[90551] = 12'h999;
rom[90552] = 12'h999;
rom[90553] = 12'h888;
rom[90554] = 12'h888;
rom[90555] = 12'h888;
rom[90556] = 12'h888;
rom[90557] = 12'h888;
rom[90558] = 12'h777;
rom[90559] = 12'h777;
rom[90560] = 12'h777;
rom[90561] = 12'h777;
rom[90562] = 12'h777;
rom[90563] = 12'h777;
rom[90564] = 12'h777;
rom[90565] = 12'h777;
rom[90566] = 12'h777;
rom[90567] = 12'h777;
rom[90568] = 12'h777;
rom[90569] = 12'h777;
rom[90570] = 12'h777;
rom[90571] = 12'h888;
rom[90572] = 12'h888;
rom[90573] = 12'h888;
rom[90574] = 12'h777;
rom[90575] = 12'h777;
rom[90576] = 12'h777;
rom[90577] = 12'h777;
rom[90578] = 12'h777;
rom[90579] = 12'h888;
rom[90580] = 12'h888;
rom[90581] = 12'h888;
rom[90582] = 12'h777;
rom[90583] = 12'h777;
rom[90584] = 12'h777;
rom[90585] = 12'h777;
rom[90586] = 12'h777;
rom[90587] = 12'h777;
rom[90588] = 12'h777;
rom[90589] = 12'h777;
rom[90590] = 12'h777;
rom[90591] = 12'h777;
rom[90592] = 12'h666;
rom[90593] = 12'h666;
rom[90594] = 12'h666;
rom[90595] = 12'h777;
rom[90596] = 12'h666;
rom[90597] = 12'h666;
rom[90598] = 12'h666;
rom[90599] = 12'h666;
rom[90600] = 12'h666;
rom[90601] = 12'h666;
rom[90602] = 12'h666;
rom[90603] = 12'h555;
rom[90604] = 12'h555;
rom[90605] = 12'h555;
rom[90606] = 12'h555;
rom[90607] = 12'h555;
rom[90608] = 12'h555;
rom[90609] = 12'h555;
rom[90610] = 12'h444;
rom[90611] = 12'h444;
rom[90612] = 12'h444;
rom[90613] = 12'h444;
rom[90614] = 12'h333;
rom[90615] = 12'h333;
rom[90616] = 12'h333;
rom[90617] = 12'h222;
rom[90618] = 12'h222;
rom[90619] = 12'h222;
rom[90620] = 12'h222;
rom[90621] = 12'h222;
rom[90622] = 12'h222;
rom[90623] = 12'h222;
rom[90624] = 12'h444;
rom[90625] = 12'h555;
rom[90626] = 12'h777;
rom[90627] = 12'h777;
rom[90628] = 12'h777;
rom[90629] = 12'h666;
rom[90630] = 12'h555;
rom[90631] = 12'h555;
rom[90632] = 12'h444;
rom[90633] = 12'h444;
rom[90634] = 12'h333;
rom[90635] = 12'h333;
rom[90636] = 12'h222;
rom[90637] = 12'h222;
rom[90638] = 12'h222;
rom[90639] = 12'h222;
rom[90640] = 12'h222;
rom[90641] = 12'h111;
rom[90642] = 12'h111;
rom[90643] = 12'h111;
rom[90644] = 12'h111;
rom[90645] = 12'h111;
rom[90646] = 12'h  0;
rom[90647] = 12'h  0;
rom[90648] = 12'h  0;
rom[90649] = 12'h  0;
rom[90650] = 12'h  0;
rom[90651] = 12'h  0;
rom[90652] = 12'h  0;
rom[90653] = 12'h  0;
rom[90654] = 12'h  0;
rom[90655] = 12'h  0;
rom[90656] = 12'h  0;
rom[90657] = 12'h  0;
rom[90658] = 12'h  0;
rom[90659] = 12'h  0;
rom[90660] = 12'h  0;
rom[90661] = 12'h  0;
rom[90662] = 12'h111;
rom[90663] = 12'h111;
rom[90664] = 12'h111;
rom[90665] = 12'h111;
rom[90666] = 12'h111;
rom[90667] = 12'h111;
rom[90668] = 12'h111;
rom[90669] = 12'h111;
rom[90670] = 12'h222;
rom[90671] = 12'h222;
rom[90672] = 12'h222;
rom[90673] = 12'h222;
rom[90674] = 12'h333;
rom[90675] = 12'h444;
rom[90676] = 12'h444;
rom[90677] = 12'h666;
rom[90678] = 12'h777;
rom[90679] = 12'h888;
rom[90680] = 12'h888;
rom[90681] = 12'h888;
rom[90682] = 12'h888;
rom[90683] = 12'h888;
rom[90684] = 12'h777;
rom[90685] = 12'h777;
rom[90686] = 12'h777;
rom[90687] = 12'h777;
rom[90688] = 12'h777;
rom[90689] = 12'h777;
rom[90690] = 12'h777;
rom[90691] = 12'h888;
rom[90692] = 12'h888;
rom[90693] = 12'h888;
rom[90694] = 12'h999;
rom[90695] = 12'h999;
rom[90696] = 12'haaa;
rom[90697] = 12'haaa;
rom[90698] = 12'hbbb;
rom[90699] = 12'hccc;
rom[90700] = 12'hddd;
rom[90701] = 12'hddd;
rom[90702] = 12'hbbb;
rom[90703] = 12'haaa;
rom[90704] = 12'h888;
rom[90705] = 12'h888;
rom[90706] = 12'h888;
rom[90707] = 12'h777;
rom[90708] = 12'h777;
rom[90709] = 12'h666;
rom[90710] = 12'h555;
rom[90711] = 12'h555;
rom[90712] = 12'h444;
rom[90713] = 12'h444;
rom[90714] = 12'h444;
rom[90715] = 12'h444;
rom[90716] = 12'h444;
rom[90717] = 12'h444;
rom[90718] = 12'h444;
rom[90719] = 12'h333;
rom[90720] = 12'h444;
rom[90721] = 12'h444;
rom[90722] = 12'h333;
rom[90723] = 12'h333;
rom[90724] = 12'h333;
rom[90725] = 12'h333;
rom[90726] = 12'h333;
rom[90727] = 12'h333;
rom[90728] = 12'h333;
rom[90729] = 12'h333;
rom[90730] = 12'h333;
rom[90731] = 12'h333;
rom[90732] = 12'h333;
rom[90733] = 12'h333;
rom[90734] = 12'h333;
rom[90735] = 12'h333;
rom[90736] = 12'h333;
rom[90737] = 12'h333;
rom[90738] = 12'h333;
rom[90739] = 12'h333;
rom[90740] = 12'h333;
rom[90741] = 12'h333;
rom[90742] = 12'h333;
rom[90743] = 12'h222;
rom[90744] = 12'h222;
rom[90745] = 12'h333;
rom[90746] = 12'h333;
rom[90747] = 12'h333;
rom[90748] = 12'h444;
rom[90749] = 12'h444;
rom[90750] = 12'h666;
rom[90751] = 12'h777;
rom[90752] = 12'h999;
rom[90753] = 12'haaa;
rom[90754] = 12'hccc;
rom[90755] = 12'heee;
rom[90756] = 12'hfff;
rom[90757] = 12'hfff;
rom[90758] = 12'hddd;
rom[90759] = 12'hccc;
rom[90760] = 12'haaa;
rom[90761] = 12'h888;
rom[90762] = 12'h777;
rom[90763] = 12'h666;
rom[90764] = 12'h555;
rom[90765] = 12'h555;
rom[90766] = 12'h555;
rom[90767] = 12'h555;
rom[90768] = 12'h444;
rom[90769] = 12'h444;
rom[90770] = 12'h444;
rom[90771] = 12'h444;
rom[90772] = 12'h444;
rom[90773] = 12'h444;
rom[90774] = 12'h333;
rom[90775] = 12'h333;
rom[90776] = 12'h333;
rom[90777] = 12'h333;
rom[90778] = 12'h333;
rom[90779] = 12'h333;
rom[90780] = 12'h333;
rom[90781] = 12'h222;
rom[90782] = 12'h222;
rom[90783] = 12'h222;
rom[90784] = 12'h222;
rom[90785] = 12'h222;
rom[90786] = 12'h222;
rom[90787] = 12'h333;
rom[90788] = 12'h333;
rom[90789] = 12'h333;
rom[90790] = 12'h444;
rom[90791] = 12'h444;
rom[90792] = 12'h444;
rom[90793] = 12'h555;
rom[90794] = 12'h555;
rom[90795] = 12'h666;
rom[90796] = 12'h666;
rom[90797] = 12'h666;
rom[90798] = 12'h777;
rom[90799] = 12'h777;
rom[90800] = 12'hfff;
rom[90801] = 12'hfff;
rom[90802] = 12'hfff;
rom[90803] = 12'hfff;
rom[90804] = 12'hfff;
rom[90805] = 12'hfff;
rom[90806] = 12'hfff;
rom[90807] = 12'hfff;
rom[90808] = 12'hfff;
rom[90809] = 12'hfff;
rom[90810] = 12'hfff;
rom[90811] = 12'hfff;
rom[90812] = 12'hfff;
rom[90813] = 12'hfff;
rom[90814] = 12'hfff;
rom[90815] = 12'hfff;
rom[90816] = 12'hfff;
rom[90817] = 12'hfff;
rom[90818] = 12'hfff;
rom[90819] = 12'hfff;
rom[90820] = 12'hfff;
rom[90821] = 12'hfff;
rom[90822] = 12'hfff;
rom[90823] = 12'hfff;
rom[90824] = 12'hfff;
rom[90825] = 12'hfff;
rom[90826] = 12'hfff;
rom[90827] = 12'hfff;
rom[90828] = 12'hfff;
rom[90829] = 12'hfff;
rom[90830] = 12'hfff;
rom[90831] = 12'hfff;
rom[90832] = 12'hfff;
rom[90833] = 12'hfff;
rom[90834] = 12'hfff;
rom[90835] = 12'hfff;
rom[90836] = 12'hfff;
rom[90837] = 12'hfff;
rom[90838] = 12'hfff;
rom[90839] = 12'hfff;
rom[90840] = 12'hfff;
rom[90841] = 12'hfff;
rom[90842] = 12'hfff;
rom[90843] = 12'hfff;
rom[90844] = 12'hfff;
rom[90845] = 12'hfff;
rom[90846] = 12'hfff;
rom[90847] = 12'hfff;
rom[90848] = 12'hfff;
rom[90849] = 12'hfff;
rom[90850] = 12'hfff;
rom[90851] = 12'hfff;
rom[90852] = 12'hfff;
rom[90853] = 12'hfff;
rom[90854] = 12'hfff;
rom[90855] = 12'hfff;
rom[90856] = 12'hfff;
rom[90857] = 12'hfff;
rom[90858] = 12'hfff;
rom[90859] = 12'hfff;
rom[90860] = 12'hfff;
rom[90861] = 12'hfff;
rom[90862] = 12'hfff;
rom[90863] = 12'hfff;
rom[90864] = 12'hfff;
rom[90865] = 12'hfff;
rom[90866] = 12'hfff;
rom[90867] = 12'hfff;
rom[90868] = 12'hfff;
rom[90869] = 12'hfff;
rom[90870] = 12'hfff;
rom[90871] = 12'hfff;
rom[90872] = 12'hfff;
rom[90873] = 12'hfff;
rom[90874] = 12'hfff;
rom[90875] = 12'hfff;
rom[90876] = 12'hfff;
rom[90877] = 12'hfff;
rom[90878] = 12'hfff;
rom[90879] = 12'hfff;
rom[90880] = 12'hfff;
rom[90881] = 12'hfff;
rom[90882] = 12'hfff;
rom[90883] = 12'hfff;
rom[90884] = 12'hfff;
rom[90885] = 12'hfff;
rom[90886] = 12'hfff;
rom[90887] = 12'hfff;
rom[90888] = 12'hfff;
rom[90889] = 12'hfff;
rom[90890] = 12'hfff;
rom[90891] = 12'hfff;
rom[90892] = 12'hfff;
rom[90893] = 12'hfff;
rom[90894] = 12'hfff;
rom[90895] = 12'hfff;
rom[90896] = 12'hfff;
rom[90897] = 12'hfff;
rom[90898] = 12'hfff;
rom[90899] = 12'hfff;
rom[90900] = 12'hfff;
rom[90901] = 12'hfff;
rom[90902] = 12'hfff;
rom[90903] = 12'hfff;
rom[90904] = 12'hfff;
rom[90905] = 12'hfff;
rom[90906] = 12'hfff;
rom[90907] = 12'hfff;
rom[90908] = 12'hfff;
rom[90909] = 12'hfff;
rom[90910] = 12'hfff;
rom[90911] = 12'hfff;
rom[90912] = 12'hfff;
rom[90913] = 12'hfff;
rom[90914] = 12'hfff;
rom[90915] = 12'hfff;
rom[90916] = 12'hfff;
rom[90917] = 12'hfff;
rom[90918] = 12'hfff;
rom[90919] = 12'hfff;
rom[90920] = 12'hfff;
rom[90921] = 12'hfff;
rom[90922] = 12'hfff;
rom[90923] = 12'hfff;
rom[90924] = 12'hfff;
rom[90925] = 12'hfff;
rom[90926] = 12'hfff;
rom[90927] = 12'hfff;
rom[90928] = 12'hfff;
rom[90929] = 12'hfff;
rom[90930] = 12'hfff;
rom[90931] = 12'hfff;
rom[90932] = 12'hfff;
rom[90933] = 12'hfff;
rom[90934] = 12'heee;
rom[90935] = 12'heee;
rom[90936] = 12'heee;
rom[90937] = 12'hddd;
rom[90938] = 12'hddd;
rom[90939] = 12'hddd;
rom[90940] = 12'hccc;
rom[90941] = 12'hccc;
rom[90942] = 12'hbbb;
rom[90943] = 12'hbbb;
rom[90944] = 12'haaa;
rom[90945] = 12'haaa;
rom[90946] = 12'haaa;
rom[90947] = 12'h999;
rom[90948] = 12'h999;
rom[90949] = 12'h999;
rom[90950] = 12'h999;
rom[90951] = 12'h999;
rom[90952] = 12'h999;
rom[90953] = 12'h999;
rom[90954] = 12'h888;
rom[90955] = 12'h888;
rom[90956] = 12'h888;
rom[90957] = 12'h888;
rom[90958] = 12'h888;
rom[90959] = 12'h777;
rom[90960] = 12'h777;
rom[90961] = 12'h777;
rom[90962] = 12'h777;
rom[90963] = 12'h777;
rom[90964] = 12'h777;
rom[90965] = 12'h777;
rom[90966] = 12'h777;
rom[90967] = 12'h777;
rom[90968] = 12'h777;
rom[90969] = 12'h777;
rom[90970] = 12'h777;
rom[90971] = 12'h777;
rom[90972] = 12'h777;
rom[90973] = 12'h777;
rom[90974] = 12'h777;
rom[90975] = 12'h777;
rom[90976] = 12'h777;
rom[90977] = 12'h777;
rom[90978] = 12'h777;
rom[90979] = 12'h888;
rom[90980] = 12'h888;
rom[90981] = 12'h888;
rom[90982] = 12'h888;
rom[90983] = 12'h777;
rom[90984] = 12'h777;
rom[90985] = 12'h777;
rom[90986] = 12'h777;
rom[90987] = 12'h777;
rom[90988] = 12'h777;
rom[90989] = 12'h777;
rom[90990] = 12'h777;
rom[90991] = 12'h777;
rom[90992] = 12'h666;
rom[90993] = 12'h777;
rom[90994] = 12'h777;
rom[90995] = 12'h777;
rom[90996] = 12'h777;
rom[90997] = 12'h777;
rom[90998] = 12'h666;
rom[90999] = 12'h666;
rom[91000] = 12'h666;
rom[91001] = 12'h666;
rom[91002] = 12'h666;
rom[91003] = 12'h666;
rom[91004] = 12'h555;
rom[91005] = 12'h555;
rom[91006] = 12'h555;
rom[91007] = 12'h555;
rom[91008] = 12'h555;
rom[91009] = 12'h555;
rom[91010] = 12'h444;
rom[91011] = 12'h444;
rom[91012] = 12'h444;
rom[91013] = 12'h444;
rom[91014] = 12'h333;
rom[91015] = 12'h333;
rom[91016] = 12'h333;
rom[91017] = 12'h333;
rom[91018] = 12'h222;
rom[91019] = 12'h222;
rom[91020] = 12'h222;
rom[91021] = 12'h222;
rom[91022] = 12'h222;
rom[91023] = 12'h222;
rom[91024] = 12'h333;
rom[91025] = 12'h444;
rom[91026] = 12'h555;
rom[91027] = 12'h777;
rom[91028] = 12'h888;
rom[91029] = 12'h777;
rom[91030] = 12'h666;
rom[91031] = 12'h666;
rom[91032] = 12'h555;
rom[91033] = 12'h444;
rom[91034] = 12'h444;
rom[91035] = 12'h333;
rom[91036] = 12'h333;
rom[91037] = 12'h222;
rom[91038] = 12'h222;
rom[91039] = 12'h222;
rom[91040] = 12'h222;
rom[91041] = 12'h222;
rom[91042] = 12'h111;
rom[91043] = 12'h111;
rom[91044] = 12'h111;
rom[91045] = 12'h111;
rom[91046] = 12'h  0;
rom[91047] = 12'h  0;
rom[91048] = 12'h  0;
rom[91049] = 12'h  0;
rom[91050] = 12'h  0;
rom[91051] = 12'h  0;
rom[91052] = 12'h  0;
rom[91053] = 12'h  0;
rom[91054] = 12'h  0;
rom[91055] = 12'h  0;
rom[91056] = 12'h  0;
rom[91057] = 12'h  0;
rom[91058] = 12'h  0;
rom[91059] = 12'h  0;
rom[91060] = 12'h  0;
rom[91061] = 12'h111;
rom[91062] = 12'h111;
rom[91063] = 12'h111;
rom[91064] = 12'h111;
rom[91065] = 12'h111;
rom[91066] = 12'h111;
rom[91067] = 12'h111;
rom[91068] = 12'h111;
rom[91069] = 12'h222;
rom[91070] = 12'h222;
rom[91071] = 12'h222;
rom[91072] = 12'h222;
rom[91073] = 12'h222;
rom[91074] = 12'h333;
rom[91075] = 12'h444;
rom[91076] = 12'h555;
rom[91077] = 12'h666;
rom[91078] = 12'h888;
rom[91079] = 12'h888;
rom[91080] = 12'h888;
rom[91081] = 12'h888;
rom[91082] = 12'h888;
rom[91083] = 12'h777;
rom[91084] = 12'h777;
rom[91085] = 12'h777;
rom[91086] = 12'h777;
rom[91087] = 12'h777;
rom[91088] = 12'h777;
rom[91089] = 12'h777;
rom[91090] = 12'h777;
rom[91091] = 12'h888;
rom[91092] = 12'h888;
rom[91093] = 12'h888;
rom[91094] = 12'h999;
rom[91095] = 12'h999;
rom[91096] = 12'h999;
rom[91097] = 12'haaa;
rom[91098] = 12'hccc;
rom[91099] = 12'hddd;
rom[91100] = 12'hddd;
rom[91101] = 12'hccc;
rom[91102] = 12'haaa;
rom[91103] = 12'h999;
rom[91104] = 12'h888;
rom[91105] = 12'h888;
rom[91106] = 12'h888;
rom[91107] = 12'h888;
rom[91108] = 12'h777;
rom[91109] = 12'h666;
rom[91110] = 12'h555;
rom[91111] = 12'h555;
rom[91112] = 12'h444;
rom[91113] = 12'h444;
rom[91114] = 12'h444;
rom[91115] = 12'h444;
rom[91116] = 12'h444;
rom[91117] = 12'h444;
rom[91118] = 12'h444;
rom[91119] = 12'h333;
rom[91120] = 12'h333;
rom[91121] = 12'h333;
rom[91122] = 12'h333;
rom[91123] = 12'h333;
rom[91124] = 12'h333;
rom[91125] = 12'h333;
rom[91126] = 12'h333;
rom[91127] = 12'h333;
rom[91128] = 12'h333;
rom[91129] = 12'h333;
rom[91130] = 12'h333;
rom[91131] = 12'h333;
rom[91132] = 12'h333;
rom[91133] = 12'h333;
rom[91134] = 12'h333;
rom[91135] = 12'h333;
rom[91136] = 12'h333;
rom[91137] = 12'h333;
rom[91138] = 12'h333;
rom[91139] = 12'h333;
rom[91140] = 12'h333;
rom[91141] = 12'h333;
rom[91142] = 12'h333;
rom[91143] = 12'h222;
rom[91144] = 12'h333;
rom[91145] = 12'h333;
rom[91146] = 12'h333;
rom[91147] = 12'h333;
rom[91148] = 12'h333;
rom[91149] = 12'h333;
rom[91150] = 12'h444;
rom[91151] = 12'h555;
rom[91152] = 12'h666;
rom[91153] = 12'h777;
rom[91154] = 12'h888;
rom[91155] = 12'hbbb;
rom[91156] = 12'hddd;
rom[91157] = 12'heee;
rom[91158] = 12'hfff;
rom[91159] = 12'hfff;
rom[91160] = 12'hddd;
rom[91161] = 12'hccc;
rom[91162] = 12'h999;
rom[91163] = 12'h777;
rom[91164] = 12'h666;
rom[91165] = 12'h666;
rom[91166] = 12'h666;
rom[91167] = 12'h555;
rom[91168] = 12'h444;
rom[91169] = 12'h444;
rom[91170] = 12'h444;
rom[91171] = 12'h444;
rom[91172] = 12'h444;
rom[91173] = 12'h333;
rom[91174] = 12'h333;
rom[91175] = 12'h333;
rom[91176] = 12'h333;
rom[91177] = 12'h333;
rom[91178] = 12'h333;
rom[91179] = 12'h333;
rom[91180] = 12'h333;
rom[91181] = 12'h222;
rom[91182] = 12'h222;
rom[91183] = 12'h333;
rom[91184] = 12'h222;
rom[91185] = 12'h222;
rom[91186] = 12'h222;
rom[91187] = 12'h222;
rom[91188] = 12'h222;
rom[91189] = 12'h222;
rom[91190] = 12'h333;
rom[91191] = 12'h333;
rom[91192] = 12'h333;
rom[91193] = 12'h333;
rom[91194] = 12'h333;
rom[91195] = 12'h444;
rom[91196] = 12'h444;
rom[91197] = 12'h555;
rom[91198] = 12'h555;
rom[91199] = 12'h555;
rom[91200] = 12'hfff;
rom[91201] = 12'hfff;
rom[91202] = 12'hfff;
rom[91203] = 12'hfff;
rom[91204] = 12'hfff;
rom[91205] = 12'hfff;
rom[91206] = 12'hfff;
rom[91207] = 12'hfff;
rom[91208] = 12'hfff;
rom[91209] = 12'hfff;
rom[91210] = 12'hfff;
rom[91211] = 12'hfff;
rom[91212] = 12'hfff;
rom[91213] = 12'hfff;
rom[91214] = 12'hfff;
rom[91215] = 12'hfff;
rom[91216] = 12'hfff;
rom[91217] = 12'hfff;
rom[91218] = 12'hfff;
rom[91219] = 12'hfff;
rom[91220] = 12'hfff;
rom[91221] = 12'hfff;
rom[91222] = 12'hfff;
rom[91223] = 12'hfff;
rom[91224] = 12'hfff;
rom[91225] = 12'hfff;
rom[91226] = 12'hfff;
rom[91227] = 12'hfff;
rom[91228] = 12'hfff;
rom[91229] = 12'hfff;
rom[91230] = 12'hfff;
rom[91231] = 12'hfff;
rom[91232] = 12'hfff;
rom[91233] = 12'hfff;
rom[91234] = 12'hfff;
rom[91235] = 12'hfff;
rom[91236] = 12'hfff;
rom[91237] = 12'hfff;
rom[91238] = 12'hfff;
rom[91239] = 12'hfff;
rom[91240] = 12'hfff;
rom[91241] = 12'hfff;
rom[91242] = 12'hfff;
rom[91243] = 12'hfff;
rom[91244] = 12'hfff;
rom[91245] = 12'hfff;
rom[91246] = 12'hfff;
rom[91247] = 12'hfff;
rom[91248] = 12'hfff;
rom[91249] = 12'hfff;
rom[91250] = 12'hfff;
rom[91251] = 12'hfff;
rom[91252] = 12'hfff;
rom[91253] = 12'hfff;
rom[91254] = 12'hfff;
rom[91255] = 12'hfff;
rom[91256] = 12'hfff;
rom[91257] = 12'hfff;
rom[91258] = 12'hfff;
rom[91259] = 12'hfff;
rom[91260] = 12'hfff;
rom[91261] = 12'hfff;
rom[91262] = 12'hfff;
rom[91263] = 12'hfff;
rom[91264] = 12'hfff;
rom[91265] = 12'hfff;
rom[91266] = 12'hfff;
rom[91267] = 12'hfff;
rom[91268] = 12'hfff;
rom[91269] = 12'hfff;
rom[91270] = 12'hfff;
rom[91271] = 12'hfff;
rom[91272] = 12'hfff;
rom[91273] = 12'hfff;
rom[91274] = 12'hfff;
rom[91275] = 12'hfff;
rom[91276] = 12'hfff;
rom[91277] = 12'hfff;
rom[91278] = 12'hfff;
rom[91279] = 12'hfff;
rom[91280] = 12'hfff;
rom[91281] = 12'hfff;
rom[91282] = 12'hfff;
rom[91283] = 12'hfff;
rom[91284] = 12'hfff;
rom[91285] = 12'hfff;
rom[91286] = 12'hfff;
rom[91287] = 12'hfff;
rom[91288] = 12'hfff;
rom[91289] = 12'hfff;
rom[91290] = 12'hfff;
rom[91291] = 12'hfff;
rom[91292] = 12'hfff;
rom[91293] = 12'hfff;
rom[91294] = 12'hfff;
rom[91295] = 12'hfff;
rom[91296] = 12'hfff;
rom[91297] = 12'hfff;
rom[91298] = 12'hfff;
rom[91299] = 12'hfff;
rom[91300] = 12'hfff;
rom[91301] = 12'hfff;
rom[91302] = 12'hfff;
rom[91303] = 12'hfff;
rom[91304] = 12'hfff;
rom[91305] = 12'hfff;
rom[91306] = 12'hfff;
rom[91307] = 12'hfff;
rom[91308] = 12'hfff;
rom[91309] = 12'hfff;
rom[91310] = 12'hfff;
rom[91311] = 12'hfff;
rom[91312] = 12'hfff;
rom[91313] = 12'hfff;
rom[91314] = 12'hfff;
rom[91315] = 12'hfff;
rom[91316] = 12'hfff;
rom[91317] = 12'hfff;
rom[91318] = 12'hfff;
rom[91319] = 12'hfff;
rom[91320] = 12'hfff;
rom[91321] = 12'hfff;
rom[91322] = 12'hfff;
rom[91323] = 12'hfff;
rom[91324] = 12'hfff;
rom[91325] = 12'hfff;
rom[91326] = 12'hfff;
rom[91327] = 12'hfff;
rom[91328] = 12'hfff;
rom[91329] = 12'hfff;
rom[91330] = 12'hfff;
rom[91331] = 12'hfff;
rom[91332] = 12'hfff;
rom[91333] = 12'hfff;
rom[91334] = 12'hfff;
rom[91335] = 12'hfff;
rom[91336] = 12'heee;
rom[91337] = 12'heee;
rom[91338] = 12'heee;
rom[91339] = 12'hddd;
rom[91340] = 12'hddd;
rom[91341] = 12'hccc;
rom[91342] = 12'hccc;
rom[91343] = 12'hbbb;
rom[91344] = 12'hbbb;
rom[91345] = 12'haaa;
rom[91346] = 12'haaa;
rom[91347] = 12'haaa;
rom[91348] = 12'h999;
rom[91349] = 12'h999;
rom[91350] = 12'h999;
rom[91351] = 12'h999;
rom[91352] = 12'h999;
rom[91353] = 12'h999;
rom[91354] = 12'h999;
rom[91355] = 12'h999;
rom[91356] = 12'h888;
rom[91357] = 12'h888;
rom[91358] = 12'h888;
rom[91359] = 12'h888;
rom[91360] = 12'h777;
rom[91361] = 12'h777;
rom[91362] = 12'h777;
rom[91363] = 12'h777;
rom[91364] = 12'h777;
rom[91365] = 12'h777;
rom[91366] = 12'h777;
rom[91367] = 12'h777;
rom[91368] = 12'h777;
rom[91369] = 12'h777;
rom[91370] = 12'h777;
rom[91371] = 12'h777;
rom[91372] = 12'h777;
rom[91373] = 12'h777;
rom[91374] = 12'h777;
rom[91375] = 12'h777;
rom[91376] = 12'h777;
rom[91377] = 12'h777;
rom[91378] = 12'h777;
rom[91379] = 12'h777;
rom[91380] = 12'h777;
rom[91381] = 12'h777;
rom[91382] = 12'h777;
rom[91383] = 12'h777;
rom[91384] = 12'h777;
rom[91385] = 12'h777;
rom[91386] = 12'h777;
rom[91387] = 12'h777;
rom[91388] = 12'h777;
rom[91389] = 12'h777;
rom[91390] = 12'h777;
rom[91391] = 12'h777;
rom[91392] = 12'h777;
rom[91393] = 12'h777;
rom[91394] = 12'h777;
rom[91395] = 12'h777;
rom[91396] = 12'h777;
rom[91397] = 12'h777;
rom[91398] = 12'h666;
rom[91399] = 12'h666;
rom[91400] = 12'h666;
rom[91401] = 12'h666;
rom[91402] = 12'h666;
rom[91403] = 12'h666;
rom[91404] = 12'h666;
rom[91405] = 12'h555;
rom[91406] = 12'h555;
rom[91407] = 12'h555;
rom[91408] = 12'h555;
rom[91409] = 12'h555;
rom[91410] = 12'h555;
rom[91411] = 12'h444;
rom[91412] = 12'h444;
rom[91413] = 12'h444;
rom[91414] = 12'h444;
rom[91415] = 12'h333;
rom[91416] = 12'h333;
rom[91417] = 12'h333;
rom[91418] = 12'h222;
rom[91419] = 12'h222;
rom[91420] = 12'h222;
rom[91421] = 12'h222;
rom[91422] = 12'h222;
rom[91423] = 12'h222;
rom[91424] = 12'h222;
rom[91425] = 12'h333;
rom[91426] = 12'h444;
rom[91427] = 12'h666;
rom[91428] = 12'h777;
rom[91429] = 12'h888;
rom[91430] = 12'h777;
rom[91431] = 12'h777;
rom[91432] = 12'h666;
rom[91433] = 12'h555;
rom[91434] = 12'h555;
rom[91435] = 12'h444;
rom[91436] = 12'h333;
rom[91437] = 12'h222;
rom[91438] = 12'h222;
rom[91439] = 12'h222;
rom[91440] = 12'h222;
rom[91441] = 12'h222;
rom[91442] = 12'h222;
rom[91443] = 12'h111;
rom[91444] = 12'h111;
rom[91445] = 12'h111;
rom[91446] = 12'h111;
rom[91447] = 12'h  0;
rom[91448] = 12'h  0;
rom[91449] = 12'h  0;
rom[91450] = 12'h  0;
rom[91451] = 12'h  0;
rom[91452] = 12'h  0;
rom[91453] = 12'h  0;
rom[91454] = 12'h  0;
rom[91455] = 12'h111;
rom[91456] = 12'h  0;
rom[91457] = 12'h  0;
rom[91458] = 12'h  0;
rom[91459] = 12'h  0;
rom[91460] = 12'h111;
rom[91461] = 12'h111;
rom[91462] = 12'h111;
rom[91463] = 12'h111;
rom[91464] = 12'h111;
rom[91465] = 12'h111;
rom[91466] = 12'h111;
rom[91467] = 12'h111;
rom[91468] = 12'h111;
rom[91469] = 12'h222;
rom[91470] = 12'h222;
rom[91471] = 12'h222;
rom[91472] = 12'h333;
rom[91473] = 12'h333;
rom[91474] = 12'h444;
rom[91475] = 12'h555;
rom[91476] = 12'h666;
rom[91477] = 12'h777;
rom[91478] = 12'h888;
rom[91479] = 12'h999;
rom[91480] = 12'h888;
rom[91481] = 12'h888;
rom[91482] = 12'h888;
rom[91483] = 12'h777;
rom[91484] = 12'h777;
rom[91485] = 12'h777;
rom[91486] = 12'h777;
rom[91487] = 12'h777;
rom[91488] = 12'h777;
rom[91489] = 12'h777;
rom[91490] = 12'h777;
rom[91491] = 12'h888;
rom[91492] = 12'h888;
rom[91493] = 12'h888;
rom[91494] = 12'h999;
rom[91495] = 12'h999;
rom[91496] = 12'h999;
rom[91497] = 12'hbbb;
rom[91498] = 12'hddd;
rom[91499] = 12'hddd;
rom[91500] = 12'hddd;
rom[91501] = 12'hbbb;
rom[91502] = 12'haaa;
rom[91503] = 12'h999;
rom[91504] = 12'h999;
rom[91505] = 12'h999;
rom[91506] = 12'h888;
rom[91507] = 12'h888;
rom[91508] = 12'h888;
rom[91509] = 12'h777;
rom[91510] = 12'h555;
rom[91511] = 12'h555;
rom[91512] = 12'h444;
rom[91513] = 12'h444;
rom[91514] = 12'h444;
rom[91515] = 12'h444;
rom[91516] = 12'h444;
rom[91517] = 12'h444;
rom[91518] = 12'h333;
rom[91519] = 12'h333;
rom[91520] = 12'h333;
rom[91521] = 12'h333;
rom[91522] = 12'h333;
rom[91523] = 12'h333;
rom[91524] = 12'h333;
rom[91525] = 12'h333;
rom[91526] = 12'h333;
rom[91527] = 12'h333;
rom[91528] = 12'h333;
rom[91529] = 12'h333;
rom[91530] = 12'h333;
rom[91531] = 12'h333;
rom[91532] = 12'h333;
rom[91533] = 12'h333;
rom[91534] = 12'h333;
rom[91535] = 12'h333;
rom[91536] = 12'h333;
rom[91537] = 12'h333;
rom[91538] = 12'h333;
rom[91539] = 12'h333;
rom[91540] = 12'h333;
rom[91541] = 12'h333;
rom[91542] = 12'h222;
rom[91543] = 12'h222;
rom[91544] = 12'h222;
rom[91545] = 12'h222;
rom[91546] = 12'h333;
rom[91547] = 12'h333;
rom[91548] = 12'h333;
rom[91549] = 12'h333;
rom[91550] = 12'h333;
rom[91551] = 12'h333;
rom[91552] = 12'h444;
rom[91553] = 12'h444;
rom[91554] = 12'h555;
rom[91555] = 12'h666;
rom[91556] = 12'h888;
rom[91557] = 12'hbbb;
rom[91558] = 12'hddd;
rom[91559] = 12'heee;
rom[91560] = 12'hfff;
rom[91561] = 12'heee;
rom[91562] = 12'hddd;
rom[91563] = 12'hbbb;
rom[91564] = 12'h999;
rom[91565] = 12'h888;
rom[91566] = 12'h666;
rom[91567] = 12'h555;
rom[91568] = 12'h555;
rom[91569] = 12'h555;
rom[91570] = 12'h444;
rom[91571] = 12'h444;
rom[91572] = 12'h444;
rom[91573] = 12'h444;
rom[91574] = 12'h333;
rom[91575] = 12'h333;
rom[91576] = 12'h333;
rom[91577] = 12'h333;
rom[91578] = 12'h333;
rom[91579] = 12'h222;
rom[91580] = 12'h222;
rom[91581] = 12'h222;
rom[91582] = 12'h222;
rom[91583] = 12'h333;
rom[91584] = 12'h222;
rom[91585] = 12'h222;
rom[91586] = 12'h222;
rom[91587] = 12'h222;
rom[91588] = 12'h222;
rom[91589] = 12'h222;
rom[91590] = 12'h222;
rom[91591] = 12'h222;
rom[91592] = 12'h222;
rom[91593] = 12'h222;
rom[91594] = 12'h222;
rom[91595] = 12'h222;
rom[91596] = 12'h333;
rom[91597] = 12'h333;
rom[91598] = 12'h333;
rom[91599] = 12'h333;
rom[91600] = 12'hfff;
rom[91601] = 12'hfff;
rom[91602] = 12'hfff;
rom[91603] = 12'hfff;
rom[91604] = 12'hfff;
rom[91605] = 12'hfff;
rom[91606] = 12'hfff;
rom[91607] = 12'hfff;
rom[91608] = 12'hfff;
rom[91609] = 12'hfff;
rom[91610] = 12'hfff;
rom[91611] = 12'hfff;
rom[91612] = 12'hfff;
rom[91613] = 12'hfff;
rom[91614] = 12'hfff;
rom[91615] = 12'hfff;
rom[91616] = 12'hfff;
rom[91617] = 12'hfff;
rom[91618] = 12'hfff;
rom[91619] = 12'hfff;
rom[91620] = 12'hfff;
rom[91621] = 12'hfff;
rom[91622] = 12'hfff;
rom[91623] = 12'hfff;
rom[91624] = 12'hfff;
rom[91625] = 12'hfff;
rom[91626] = 12'hfff;
rom[91627] = 12'hfff;
rom[91628] = 12'hfff;
rom[91629] = 12'hfff;
rom[91630] = 12'hfff;
rom[91631] = 12'hfff;
rom[91632] = 12'hfff;
rom[91633] = 12'hfff;
rom[91634] = 12'hfff;
rom[91635] = 12'hfff;
rom[91636] = 12'hfff;
rom[91637] = 12'hfff;
rom[91638] = 12'hfff;
rom[91639] = 12'hfff;
rom[91640] = 12'hfff;
rom[91641] = 12'hfff;
rom[91642] = 12'hfff;
rom[91643] = 12'hfff;
rom[91644] = 12'hfff;
rom[91645] = 12'hfff;
rom[91646] = 12'hfff;
rom[91647] = 12'hfff;
rom[91648] = 12'hfff;
rom[91649] = 12'hfff;
rom[91650] = 12'hfff;
rom[91651] = 12'hfff;
rom[91652] = 12'hfff;
rom[91653] = 12'hfff;
rom[91654] = 12'hfff;
rom[91655] = 12'hfff;
rom[91656] = 12'hfff;
rom[91657] = 12'hfff;
rom[91658] = 12'hfff;
rom[91659] = 12'hfff;
rom[91660] = 12'hfff;
rom[91661] = 12'hfff;
rom[91662] = 12'hfff;
rom[91663] = 12'hfff;
rom[91664] = 12'hfff;
rom[91665] = 12'hfff;
rom[91666] = 12'hfff;
rom[91667] = 12'hfff;
rom[91668] = 12'hfff;
rom[91669] = 12'hfff;
rom[91670] = 12'hfff;
rom[91671] = 12'hfff;
rom[91672] = 12'hfff;
rom[91673] = 12'hfff;
rom[91674] = 12'hfff;
rom[91675] = 12'hfff;
rom[91676] = 12'hfff;
rom[91677] = 12'hfff;
rom[91678] = 12'hfff;
rom[91679] = 12'hfff;
rom[91680] = 12'hfff;
rom[91681] = 12'hfff;
rom[91682] = 12'hfff;
rom[91683] = 12'hfff;
rom[91684] = 12'hfff;
rom[91685] = 12'hfff;
rom[91686] = 12'hfff;
rom[91687] = 12'hfff;
rom[91688] = 12'hfff;
rom[91689] = 12'hfff;
rom[91690] = 12'hfff;
rom[91691] = 12'hfff;
rom[91692] = 12'hfff;
rom[91693] = 12'hfff;
rom[91694] = 12'hfff;
rom[91695] = 12'hfff;
rom[91696] = 12'hfff;
rom[91697] = 12'hfff;
rom[91698] = 12'hfff;
rom[91699] = 12'hfff;
rom[91700] = 12'hfff;
rom[91701] = 12'hfff;
rom[91702] = 12'hfff;
rom[91703] = 12'hfff;
rom[91704] = 12'hfff;
rom[91705] = 12'hfff;
rom[91706] = 12'hfff;
rom[91707] = 12'hfff;
rom[91708] = 12'hfff;
rom[91709] = 12'hfff;
rom[91710] = 12'hfff;
rom[91711] = 12'hfff;
rom[91712] = 12'hfff;
rom[91713] = 12'hfff;
rom[91714] = 12'hfff;
rom[91715] = 12'hfff;
rom[91716] = 12'hfff;
rom[91717] = 12'hfff;
rom[91718] = 12'hfff;
rom[91719] = 12'hfff;
rom[91720] = 12'hfff;
rom[91721] = 12'hfff;
rom[91722] = 12'hfff;
rom[91723] = 12'hfff;
rom[91724] = 12'hfff;
rom[91725] = 12'hfff;
rom[91726] = 12'hfff;
rom[91727] = 12'hfff;
rom[91728] = 12'hfff;
rom[91729] = 12'hfff;
rom[91730] = 12'hfff;
rom[91731] = 12'hfff;
rom[91732] = 12'hfff;
rom[91733] = 12'hfff;
rom[91734] = 12'hfff;
rom[91735] = 12'hfff;
rom[91736] = 12'hfff;
rom[91737] = 12'heee;
rom[91738] = 12'heee;
rom[91739] = 12'heee;
rom[91740] = 12'heee;
rom[91741] = 12'hddd;
rom[91742] = 12'hddd;
rom[91743] = 12'hccc;
rom[91744] = 12'hccc;
rom[91745] = 12'hbbb;
rom[91746] = 12'hbbb;
rom[91747] = 12'haaa;
rom[91748] = 12'haaa;
rom[91749] = 12'haaa;
rom[91750] = 12'h999;
rom[91751] = 12'h999;
rom[91752] = 12'h999;
rom[91753] = 12'h999;
rom[91754] = 12'h999;
rom[91755] = 12'h999;
rom[91756] = 12'h999;
rom[91757] = 12'h888;
rom[91758] = 12'h888;
rom[91759] = 12'h888;
rom[91760] = 12'h777;
rom[91761] = 12'h777;
rom[91762] = 12'h777;
rom[91763] = 12'h777;
rom[91764] = 12'h777;
rom[91765] = 12'h777;
rom[91766] = 12'h777;
rom[91767] = 12'h777;
rom[91768] = 12'h777;
rom[91769] = 12'h777;
rom[91770] = 12'h777;
rom[91771] = 12'h777;
rom[91772] = 12'h777;
rom[91773] = 12'h777;
rom[91774] = 12'h777;
rom[91775] = 12'h777;
rom[91776] = 12'h777;
rom[91777] = 12'h777;
rom[91778] = 12'h777;
rom[91779] = 12'h777;
rom[91780] = 12'h777;
rom[91781] = 12'h777;
rom[91782] = 12'h777;
rom[91783] = 12'h777;
rom[91784] = 12'h777;
rom[91785] = 12'h777;
rom[91786] = 12'h777;
rom[91787] = 12'h777;
rom[91788] = 12'h777;
rom[91789] = 12'h777;
rom[91790] = 12'h777;
rom[91791] = 12'h777;
rom[91792] = 12'h777;
rom[91793] = 12'h777;
rom[91794] = 12'h777;
rom[91795] = 12'h777;
rom[91796] = 12'h777;
rom[91797] = 12'h777;
rom[91798] = 12'h777;
rom[91799] = 12'h777;
rom[91800] = 12'h666;
rom[91801] = 12'h666;
rom[91802] = 12'h666;
rom[91803] = 12'h666;
rom[91804] = 12'h666;
rom[91805] = 12'h666;
rom[91806] = 12'h555;
rom[91807] = 12'h555;
rom[91808] = 12'h555;
rom[91809] = 12'h555;
rom[91810] = 12'h555;
rom[91811] = 12'h555;
rom[91812] = 12'h444;
rom[91813] = 12'h444;
rom[91814] = 12'h444;
rom[91815] = 12'h444;
rom[91816] = 12'h333;
rom[91817] = 12'h333;
rom[91818] = 12'h222;
rom[91819] = 12'h222;
rom[91820] = 12'h222;
rom[91821] = 12'h222;
rom[91822] = 12'h222;
rom[91823] = 12'h222;
rom[91824] = 12'h222;
rom[91825] = 12'h222;
rom[91826] = 12'h333;
rom[91827] = 12'h444;
rom[91828] = 12'h666;
rom[91829] = 12'h777;
rom[91830] = 12'h888;
rom[91831] = 12'h777;
rom[91832] = 12'h777;
rom[91833] = 12'h666;
rom[91834] = 12'h666;
rom[91835] = 12'h555;
rom[91836] = 12'h444;
rom[91837] = 12'h333;
rom[91838] = 12'h222;
rom[91839] = 12'h222;
rom[91840] = 12'h222;
rom[91841] = 12'h222;
rom[91842] = 12'h222;
rom[91843] = 12'h111;
rom[91844] = 12'h111;
rom[91845] = 12'h111;
rom[91846] = 12'h111;
rom[91847] = 12'h111;
rom[91848] = 12'h111;
rom[91849] = 12'h  0;
rom[91850] = 12'h  0;
rom[91851] = 12'h  0;
rom[91852] = 12'h  0;
rom[91853] = 12'h111;
rom[91854] = 12'h111;
rom[91855] = 12'h111;
rom[91856] = 12'h111;
rom[91857] = 12'h111;
rom[91858] = 12'h111;
rom[91859] = 12'h111;
rom[91860] = 12'h111;
rom[91861] = 12'h111;
rom[91862] = 12'h111;
rom[91863] = 12'h111;
rom[91864] = 12'h111;
rom[91865] = 12'h111;
rom[91866] = 12'h111;
rom[91867] = 12'h222;
rom[91868] = 12'h222;
rom[91869] = 12'h222;
rom[91870] = 12'h333;
rom[91871] = 12'h333;
rom[91872] = 12'h333;
rom[91873] = 12'h444;
rom[91874] = 12'h555;
rom[91875] = 12'h666;
rom[91876] = 12'h777;
rom[91877] = 12'h888;
rom[91878] = 12'h888;
rom[91879] = 12'h888;
rom[91880] = 12'h888;
rom[91881] = 12'h888;
rom[91882] = 12'h888;
rom[91883] = 12'h777;
rom[91884] = 12'h777;
rom[91885] = 12'h777;
rom[91886] = 12'h777;
rom[91887] = 12'h777;
rom[91888] = 12'h777;
rom[91889] = 12'h888;
rom[91890] = 12'h888;
rom[91891] = 12'h888;
rom[91892] = 12'h888;
rom[91893] = 12'h888;
rom[91894] = 12'h999;
rom[91895] = 12'h999;
rom[91896] = 12'haaa;
rom[91897] = 12'hccc;
rom[91898] = 12'hddd;
rom[91899] = 12'hddd;
rom[91900] = 12'hccc;
rom[91901] = 12'hbbb;
rom[91902] = 12'hbbb;
rom[91903] = 12'haaa;
rom[91904] = 12'haaa;
rom[91905] = 12'h999;
rom[91906] = 12'h999;
rom[91907] = 12'h999;
rom[91908] = 12'h888;
rom[91909] = 12'h777;
rom[91910] = 12'h666;
rom[91911] = 12'h555;
rom[91912] = 12'h444;
rom[91913] = 12'h444;
rom[91914] = 12'h333;
rom[91915] = 12'h333;
rom[91916] = 12'h444;
rom[91917] = 12'h444;
rom[91918] = 12'h333;
rom[91919] = 12'h333;
rom[91920] = 12'h333;
rom[91921] = 12'h333;
rom[91922] = 12'h333;
rom[91923] = 12'h444;
rom[91924] = 12'h444;
rom[91925] = 12'h333;
rom[91926] = 12'h333;
rom[91927] = 12'h333;
rom[91928] = 12'h333;
rom[91929] = 12'h333;
rom[91930] = 12'h333;
rom[91931] = 12'h333;
rom[91932] = 12'h333;
rom[91933] = 12'h333;
rom[91934] = 12'h333;
rom[91935] = 12'h333;
rom[91936] = 12'h333;
rom[91937] = 12'h333;
rom[91938] = 12'h222;
rom[91939] = 12'h222;
rom[91940] = 12'h222;
rom[91941] = 12'h222;
rom[91942] = 12'h222;
rom[91943] = 12'h222;
rom[91944] = 12'h111;
rom[91945] = 12'h222;
rom[91946] = 12'h222;
rom[91947] = 12'h222;
rom[91948] = 12'h222;
rom[91949] = 12'h222;
rom[91950] = 12'h222;
rom[91951] = 12'h333;
rom[91952] = 12'h333;
rom[91953] = 12'h333;
rom[91954] = 12'h444;
rom[91955] = 12'h444;
rom[91956] = 12'h555;
rom[91957] = 12'h666;
rom[91958] = 12'h999;
rom[91959] = 12'haaa;
rom[91960] = 12'hddd;
rom[91961] = 12'heee;
rom[91962] = 12'hfff;
rom[91963] = 12'heee;
rom[91964] = 12'hddd;
rom[91965] = 12'hbbb;
rom[91966] = 12'h888;
rom[91967] = 12'h666;
rom[91968] = 12'h555;
rom[91969] = 12'h555;
rom[91970] = 12'h444;
rom[91971] = 12'h444;
rom[91972] = 12'h444;
rom[91973] = 12'h444;
rom[91974] = 12'h444;
rom[91975] = 12'h444;
rom[91976] = 12'h333;
rom[91977] = 12'h333;
rom[91978] = 12'h333;
rom[91979] = 12'h333;
rom[91980] = 12'h222;
rom[91981] = 12'h222;
rom[91982] = 12'h222;
rom[91983] = 12'h333;
rom[91984] = 12'h222;
rom[91985] = 12'h222;
rom[91986] = 12'h222;
rom[91987] = 12'h222;
rom[91988] = 12'h222;
rom[91989] = 12'h222;
rom[91990] = 12'h222;
rom[91991] = 12'h222;
rom[91992] = 12'h222;
rom[91993] = 12'h222;
rom[91994] = 12'h222;
rom[91995] = 12'h222;
rom[91996] = 12'h222;
rom[91997] = 12'h222;
rom[91998] = 12'h222;
rom[91999] = 12'h333;
rom[92000] = 12'hfff;
rom[92001] = 12'hfff;
rom[92002] = 12'hfff;
rom[92003] = 12'hfff;
rom[92004] = 12'hfff;
rom[92005] = 12'hfff;
rom[92006] = 12'hfff;
rom[92007] = 12'hfff;
rom[92008] = 12'hfff;
rom[92009] = 12'hfff;
rom[92010] = 12'hfff;
rom[92011] = 12'hfff;
rom[92012] = 12'hfff;
rom[92013] = 12'hfff;
rom[92014] = 12'hfff;
rom[92015] = 12'hfff;
rom[92016] = 12'hfff;
rom[92017] = 12'hfff;
rom[92018] = 12'hfff;
rom[92019] = 12'hfff;
rom[92020] = 12'hfff;
rom[92021] = 12'hfff;
rom[92022] = 12'hfff;
rom[92023] = 12'hfff;
rom[92024] = 12'hfff;
rom[92025] = 12'hfff;
rom[92026] = 12'hfff;
rom[92027] = 12'hfff;
rom[92028] = 12'hfff;
rom[92029] = 12'hfff;
rom[92030] = 12'hfff;
rom[92031] = 12'hfff;
rom[92032] = 12'hfff;
rom[92033] = 12'hfff;
rom[92034] = 12'hfff;
rom[92035] = 12'hfff;
rom[92036] = 12'hfff;
rom[92037] = 12'hfff;
rom[92038] = 12'hfff;
rom[92039] = 12'hfff;
rom[92040] = 12'hfff;
rom[92041] = 12'hfff;
rom[92042] = 12'hfff;
rom[92043] = 12'hfff;
rom[92044] = 12'hfff;
rom[92045] = 12'hfff;
rom[92046] = 12'hfff;
rom[92047] = 12'hfff;
rom[92048] = 12'hfff;
rom[92049] = 12'hfff;
rom[92050] = 12'hfff;
rom[92051] = 12'hfff;
rom[92052] = 12'hfff;
rom[92053] = 12'hfff;
rom[92054] = 12'hfff;
rom[92055] = 12'hfff;
rom[92056] = 12'hfff;
rom[92057] = 12'hfff;
rom[92058] = 12'hfff;
rom[92059] = 12'hfff;
rom[92060] = 12'hfff;
rom[92061] = 12'hfff;
rom[92062] = 12'hfff;
rom[92063] = 12'hfff;
rom[92064] = 12'hfff;
rom[92065] = 12'hfff;
rom[92066] = 12'hfff;
rom[92067] = 12'hfff;
rom[92068] = 12'hfff;
rom[92069] = 12'hfff;
rom[92070] = 12'hfff;
rom[92071] = 12'hfff;
rom[92072] = 12'hfff;
rom[92073] = 12'hfff;
rom[92074] = 12'hfff;
rom[92075] = 12'hfff;
rom[92076] = 12'hfff;
rom[92077] = 12'hfff;
rom[92078] = 12'hfff;
rom[92079] = 12'hfff;
rom[92080] = 12'hfff;
rom[92081] = 12'hfff;
rom[92082] = 12'hfff;
rom[92083] = 12'hfff;
rom[92084] = 12'hfff;
rom[92085] = 12'hfff;
rom[92086] = 12'hfff;
rom[92087] = 12'hfff;
rom[92088] = 12'hfff;
rom[92089] = 12'hfff;
rom[92090] = 12'hfff;
rom[92091] = 12'hfff;
rom[92092] = 12'hfff;
rom[92093] = 12'hfff;
rom[92094] = 12'hfff;
rom[92095] = 12'hfff;
rom[92096] = 12'hfff;
rom[92097] = 12'hfff;
rom[92098] = 12'hfff;
rom[92099] = 12'hfff;
rom[92100] = 12'hfff;
rom[92101] = 12'hfff;
rom[92102] = 12'hfff;
rom[92103] = 12'hfff;
rom[92104] = 12'hfff;
rom[92105] = 12'hfff;
rom[92106] = 12'hfff;
rom[92107] = 12'hfff;
rom[92108] = 12'hfff;
rom[92109] = 12'hfff;
rom[92110] = 12'hfff;
rom[92111] = 12'hfff;
rom[92112] = 12'hfff;
rom[92113] = 12'hfff;
rom[92114] = 12'hfff;
rom[92115] = 12'hfff;
rom[92116] = 12'hfff;
rom[92117] = 12'hfff;
rom[92118] = 12'hfff;
rom[92119] = 12'hfff;
rom[92120] = 12'hfff;
rom[92121] = 12'hfff;
rom[92122] = 12'hfff;
rom[92123] = 12'hfff;
rom[92124] = 12'hfff;
rom[92125] = 12'hfff;
rom[92126] = 12'hfff;
rom[92127] = 12'hfff;
rom[92128] = 12'hfff;
rom[92129] = 12'hfff;
rom[92130] = 12'hfff;
rom[92131] = 12'hfff;
rom[92132] = 12'hfff;
rom[92133] = 12'hfff;
rom[92134] = 12'heee;
rom[92135] = 12'heee;
rom[92136] = 12'heee;
rom[92137] = 12'heee;
rom[92138] = 12'heee;
rom[92139] = 12'heee;
rom[92140] = 12'heee;
rom[92141] = 12'heee;
rom[92142] = 12'hddd;
rom[92143] = 12'hddd;
rom[92144] = 12'hddd;
rom[92145] = 12'hccc;
rom[92146] = 12'hccc;
rom[92147] = 12'hbbb;
rom[92148] = 12'hbbb;
rom[92149] = 12'haaa;
rom[92150] = 12'haaa;
rom[92151] = 12'haaa;
rom[92152] = 12'h999;
rom[92153] = 12'h999;
rom[92154] = 12'h999;
rom[92155] = 12'h999;
rom[92156] = 12'h999;
rom[92157] = 12'h999;
rom[92158] = 12'h888;
rom[92159] = 12'h888;
rom[92160] = 12'h888;
rom[92161] = 12'h888;
rom[92162] = 12'h777;
rom[92163] = 12'h777;
rom[92164] = 12'h777;
rom[92165] = 12'h777;
rom[92166] = 12'h777;
rom[92167] = 12'h777;
rom[92168] = 12'h888;
rom[92169] = 12'h888;
rom[92170] = 12'h777;
rom[92171] = 12'h777;
rom[92172] = 12'h777;
rom[92173] = 12'h777;
rom[92174] = 12'h888;
rom[92175] = 12'h888;
rom[92176] = 12'h888;
rom[92177] = 12'h888;
rom[92178] = 12'h777;
rom[92179] = 12'h777;
rom[92180] = 12'h777;
rom[92181] = 12'h777;
rom[92182] = 12'h777;
rom[92183] = 12'h777;
rom[92184] = 12'h888;
rom[92185] = 12'h888;
rom[92186] = 12'h888;
rom[92187] = 12'h888;
rom[92188] = 12'h888;
rom[92189] = 12'h888;
rom[92190] = 12'h888;
rom[92191] = 12'h888;
rom[92192] = 12'h777;
rom[92193] = 12'h777;
rom[92194] = 12'h777;
rom[92195] = 12'h777;
rom[92196] = 12'h777;
rom[92197] = 12'h777;
rom[92198] = 12'h777;
rom[92199] = 12'h777;
rom[92200] = 12'h777;
rom[92201] = 12'h777;
rom[92202] = 12'h666;
rom[92203] = 12'h666;
rom[92204] = 12'h666;
rom[92205] = 12'h666;
rom[92206] = 12'h666;
rom[92207] = 12'h666;
rom[92208] = 12'h666;
rom[92209] = 12'h555;
rom[92210] = 12'h555;
rom[92211] = 12'h555;
rom[92212] = 12'h555;
rom[92213] = 12'h444;
rom[92214] = 12'h444;
rom[92215] = 12'h444;
rom[92216] = 12'h333;
rom[92217] = 12'h333;
rom[92218] = 12'h333;
rom[92219] = 12'h333;
rom[92220] = 12'h333;
rom[92221] = 12'h222;
rom[92222] = 12'h222;
rom[92223] = 12'h222;
rom[92224] = 12'h222;
rom[92225] = 12'h222;
rom[92226] = 12'h333;
rom[92227] = 12'h444;
rom[92228] = 12'h555;
rom[92229] = 12'h666;
rom[92230] = 12'h777;
rom[92231] = 12'h777;
rom[92232] = 12'h888;
rom[92233] = 12'h777;
rom[92234] = 12'h777;
rom[92235] = 12'h666;
rom[92236] = 12'h555;
rom[92237] = 12'h444;
rom[92238] = 12'h333;
rom[92239] = 12'h333;
rom[92240] = 12'h222;
rom[92241] = 12'h222;
rom[92242] = 12'h222;
rom[92243] = 12'h222;
rom[92244] = 12'h111;
rom[92245] = 12'h111;
rom[92246] = 12'h111;
rom[92247] = 12'h111;
rom[92248] = 12'h111;
rom[92249] = 12'h111;
rom[92250] = 12'h111;
rom[92251] = 12'h111;
rom[92252] = 12'h111;
rom[92253] = 12'h111;
rom[92254] = 12'h111;
rom[92255] = 12'h111;
rom[92256] = 12'h111;
rom[92257] = 12'h111;
rom[92258] = 12'h111;
rom[92259] = 12'h111;
rom[92260] = 12'h111;
rom[92261] = 12'h111;
rom[92262] = 12'h111;
rom[92263] = 12'h111;
rom[92264] = 12'h222;
rom[92265] = 12'h222;
rom[92266] = 12'h222;
rom[92267] = 12'h222;
rom[92268] = 12'h222;
rom[92269] = 12'h222;
rom[92270] = 12'h333;
rom[92271] = 12'h333;
rom[92272] = 12'h444;
rom[92273] = 12'h444;
rom[92274] = 12'h666;
rom[92275] = 12'h777;
rom[92276] = 12'h888;
rom[92277] = 12'h888;
rom[92278] = 12'h888;
rom[92279] = 12'h888;
rom[92280] = 12'h888;
rom[92281] = 12'h888;
rom[92282] = 12'h777;
rom[92283] = 12'h777;
rom[92284] = 12'h777;
rom[92285] = 12'h777;
rom[92286] = 12'h777;
rom[92287] = 12'h777;
rom[92288] = 12'h777;
rom[92289] = 12'h888;
rom[92290] = 12'h888;
rom[92291] = 12'h888;
rom[92292] = 12'h999;
rom[92293] = 12'h999;
rom[92294] = 12'haaa;
rom[92295] = 12'haaa;
rom[92296] = 12'hbbb;
rom[92297] = 12'hddd;
rom[92298] = 12'heee;
rom[92299] = 12'hddd;
rom[92300] = 12'hccc;
rom[92301] = 12'hccc;
rom[92302] = 12'hccc;
rom[92303] = 12'hccc;
rom[92304] = 12'hccc;
rom[92305] = 12'haaa;
rom[92306] = 12'h999;
rom[92307] = 12'h999;
rom[92308] = 12'h999;
rom[92309] = 12'h888;
rom[92310] = 12'h777;
rom[92311] = 12'h666;
rom[92312] = 12'h444;
rom[92313] = 12'h444;
rom[92314] = 12'h333;
rom[92315] = 12'h333;
rom[92316] = 12'h444;
rom[92317] = 12'h444;
rom[92318] = 12'h444;
rom[92319] = 12'h333;
rom[92320] = 12'h333;
rom[92321] = 12'h333;
rom[92322] = 12'h333;
rom[92323] = 12'h444;
rom[92324] = 12'h444;
rom[92325] = 12'h444;
rom[92326] = 12'h333;
rom[92327] = 12'h333;
rom[92328] = 12'h333;
rom[92329] = 12'h333;
rom[92330] = 12'h333;
rom[92331] = 12'h333;
rom[92332] = 12'h333;
rom[92333] = 12'h333;
rom[92334] = 12'h333;
rom[92335] = 12'h333;
rom[92336] = 12'h333;
rom[92337] = 12'h222;
rom[92338] = 12'h222;
rom[92339] = 12'h222;
rom[92340] = 12'h222;
rom[92341] = 12'h222;
rom[92342] = 12'h222;
rom[92343] = 12'h222;
rom[92344] = 12'h111;
rom[92345] = 12'h222;
rom[92346] = 12'h222;
rom[92347] = 12'h222;
rom[92348] = 12'h222;
rom[92349] = 12'h222;
rom[92350] = 12'h222;
rom[92351] = 12'h222;
rom[92352] = 12'h333;
rom[92353] = 12'h333;
rom[92354] = 12'h333;
rom[92355] = 12'h333;
rom[92356] = 12'h333;
rom[92357] = 12'h444;
rom[92358] = 12'h555;
rom[92359] = 12'h666;
rom[92360] = 12'h999;
rom[92361] = 12'hbbb;
rom[92362] = 12'hddd;
rom[92363] = 12'heee;
rom[92364] = 12'heee;
rom[92365] = 12'heee;
rom[92366] = 12'hccc;
rom[92367] = 12'haaa;
rom[92368] = 12'h888;
rom[92369] = 12'h666;
rom[92370] = 12'h555;
rom[92371] = 12'h444;
rom[92372] = 12'h444;
rom[92373] = 12'h444;
rom[92374] = 12'h444;
rom[92375] = 12'h444;
rom[92376] = 12'h333;
rom[92377] = 12'h333;
rom[92378] = 12'h333;
rom[92379] = 12'h333;
rom[92380] = 12'h333;
rom[92381] = 12'h222;
rom[92382] = 12'h333;
rom[92383] = 12'h333;
rom[92384] = 12'h222;
rom[92385] = 12'h222;
rom[92386] = 12'h222;
rom[92387] = 12'h222;
rom[92388] = 12'h222;
rom[92389] = 12'h222;
rom[92390] = 12'h222;
rom[92391] = 12'h222;
rom[92392] = 12'h222;
rom[92393] = 12'h111;
rom[92394] = 12'h111;
rom[92395] = 12'h111;
rom[92396] = 12'h222;
rom[92397] = 12'h222;
rom[92398] = 12'h222;
rom[92399] = 12'h222;
rom[92400] = 12'hfff;
rom[92401] = 12'hfff;
rom[92402] = 12'hfff;
rom[92403] = 12'hfff;
rom[92404] = 12'hfff;
rom[92405] = 12'hfff;
rom[92406] = 12'hfff;
rom[92407] = 12'hfff;
rom[92408] = 12'hfff;
rom[92409] = 12'hfff;
rom[92410] = 12'hfff;
rom[92411] = 12'hfff;
rom[92412] = 12'hfff;
rom[92413] = 12'hfff;
rom[92414] = 12'hfff;
rom[92415] = 12'hfff;
rom[92416] = 12'hfff;
rom[92417] = 12'hfff;
rom[92418] = 12'hfff;
rom[92419] = 12'hfff;
rom[92420] = 12'hfff;
rom[92421] = 12'hfff;
rom[92422] = 12'hfff;
rom[92423] = 12'hfff;
rom[92424] = 12'hfff;
rom[92425] = 12'hfff;
rom[92426] = 12'hfff;
rom[92427] = 12'hfff;
rom[92428] = 12'hfff;
rom[92429] = 12'hfff;
rom[92430] = 12'hfff;
rom[92431] = 12'hfff;
rom[92432] = 12'hfff;
rom[92433] = 12'hfff;
rom[92434] = 12'hfff;
rom[92435] = 12'hfff;
rom[92436] = 12'hfff;
rom[92437] = 12'hfff;
rom[92438] = 12'hfff;
rom[92439] = 12'hfff;
rom[92440] = 12'hfff;
rom[92441] = 12'hfff;
rom[92442] = 12'hfff;
rom[92443] = 12'hfff;
rom[92444] = 12'hfff;
rom[92445] = 12'hfff;
rom[92446] = 12'hfff;
rom[92447] = 12'hfff;
rom[92448] = 12'hfff;
rom[92449] = 12'hfff;
rom[92450] = 12'hfff;
rom[92451] = 12'hfff;
rom[92452] = 12'hfff;
rom[92453] = 12'hfff;
rom[92454] = 12'hfff;
rom[92455] = 12'hfff;
rom[92456] = 12'hfff;
rom[92457] = 12'hfff;
rom[92458] = 12'hfff;
rom[92459] = 12'hfff;
rom[92460] = 12'hfff;
rom[92461] = 12'hfff;
rom[92462] = 12'hfff;
rom[92463] = 12'hfff;
rom[92464] = 12'hfff;
rom[92465] = 12'hfff;
rom[92466] = 12'hfff;
rom[92467] = 12'hfff;
rom[92468] = 12'hfff;
rom[92469] = 12'hfff;
rom[92470] = 12'hfff;
rom[92471] = 12'hfff;
rom[92472] = 12'hfff;
rom[92473] = 12'hfff;
rom[92474] = 12'hfff;
rom[92475] = 12'hfff;
rom[92476] = 12'hfff;
rom[92477] = 12'hfff;
rom[92478] = 12'hfff;
rom[92479] = 12'hfff;
rom[92480] = 12'hfff;
rom[92481] = 12'hfff;
rom[92482] = 12'hfff;
rom[92483] = 12'hfff;
rom[92484] = 12'hfff;
rom[92485] = 12'hfff;
rom[92486] = 12'hfff;
rom[92487] = 12'hfff;
rom[92488] = 12'hfff;
rom[92489] = 12'hfff;
rom[92490] = 12'hfff;
rom[92491] = 12'hfff;
rom[92492] = 12'hfff;
rom[92493] = 12'hfff;
rom[92494] = 12'hfff;
rom[92495] = 12'hfff;
rom[92496] = 12'hfff;
rom[92497] = 12'hfff;
rom[92498] = 12'hfff;
rom[92499] = 12'hfff;
rom[92500] = 12'hfff;
rom[92501] = 12'hfff;
rom[92502] = 12'hfff;
rom[92503] = 12'hfff;
rom[92504] = 12'hfff;
rom[92505] = 12'hfff;
rom[92506] = 12'hfff;
rom[92507] = 12'hfff;
rom[92508] = 12'hfff;
rom[92509] = 12'hfff;
rom[92510] = 12'hfff;
rom[92511] = 12'hfff;
rom[92512] = 12'hfff;
rom[92513] = 12'hfff;
rom[92514] = 12'hfff;
rom[92515] = 12'hfff;
rom[92516] = 12'hfff;
rom[92517] = 12'hfff;
rom[92518] = 12'hfff;
rom[92519] = 12'hfff;
rom[92520] = 12'hfff;
rom[92521] = 12'hfff;
rom[92522] = 12'hfff;
rom[92523] = 12'hfff;
rom[92524] = 12'hfff;
rom[92525] = 12'hfff;
rom[92526] = 12'hfff;
rom[92527] = 12'hfff;
rom[92528] = 12'hfff;
rom[92529] = 12'hfff;
rom[92530] = 12'hfff;
rom[92531] = 12'hfff;
rom[92532] = 12'hfff;
rom[92533] = 12'heee;
rom[92534] = 12'heee;
rom[92535] = 12'heee;
rom[92536] = 12'heee;
rom[92537] = 12'heee;
rom[92538] = 12'heee;
rom[92539] = 12'heee;
rom[92540] = 12'heee;
rom[92541] = 12'heee;
rom[92542] = 12'heee;
rom[92543] = 12'heee;
rom[92544] = 12'hddd;
rom[92545] = 12'hddd;
rom[92546] = 12'hccc;
rom[92547] = 12'hccc;
rom[92548] = 12'hccc;
rom[92549] = 12'hbbb;
rom[92550] = 12'haaa;
rom[92551] = 12'haaa;
rom[92552] = 12'h999;
rom[92553] = 12'h999;
rom[92554] = 12'h999;
rom[92555] = 12'h999;
rom[92556] = 12'h999;
rom[92557] = 12'h999;
rom[92558] = 12'h888;
rom[92559] = 12'h888;
rom[92560] = 12'h888;
rom[92561] = 12'h888;
rom[92562] = 12'h888;
rom[92563] = 12'h888;
rom[92564] = 12'h888;
rom[92565] = 12'h888;
rom[92566] = 12'h888;
rom[92567] = 12'h888;
rom[92568] = 12'h888;
rom[92569] = 12'h888;
rom[92570] = 12'h777;
rom[92571] = 12'h777;
rom[92572] = 12'h777;
rom[92573] = 12'h777;
rom[92574] = 12'h888;
rom[92575] = 12'h888;
rom[92576] = 12'h888;
rom[92577] = 12'h888;
rom[92578] = 12'h888;
rom[92579] = 12'h777;
rom[92580] = 12'h777;
rom[92581] = 12'h777;
rom[92582] = 12'h777;
rom[92583] = 12'h888;
rom[92584] = 12'h888;
rom[92585] = 12'h888;
rom[92586] = 12'h888;
rom[92587] = 12'h888;
rom[92588] = 12'h888;
rom[92589] = 12'h888;
rom[92590] = 12'h888;
rom[92591] = 12'h888;
rom[92592] = 12'h888;
rom[92593] = 12'h888;
rom[92594] = 12'h777;
rom[92595] = 12'h777;
rom[92596] = 12'h777;
rom[92597] = 12'h777;
rom[92598] = 12'h777;
rom[92599] = 12'h777;
rom[92600] = 12'h777;
rom[92601] = 12'h777;
rom[92602] = 12'h777;
rom[92603] = 12'h777;
rom[92604] = 12'h666;
rom[92605] = 12'h666;
rom[92606] = 12'h666;
rom[92607] = 12'h666;
rom[92608] = 12'h666;
rom[92609] = 12'h666;
rom[92610] = 12'h555;
rom[92611] = 12'h555;
rom[92612] = 12'h555;
rom[92613] = 12'h444;
rom[92614] = 12'h444;
rom[92615] = 12'h444;
rom[92616] = 12'h333;
rom[92617] = 12'h333;
rom[92618] = 12'h333;
rom[92619] = 12'h333;
rom[92620] = 12'h333;
rom[92621] = 12'h333;
rom[92622] = 12'h222;
rom[92623] = 12'h222;
rom[92624] = 12'h222;
rom[92625] = 12'h222;
rom[92626] = 12'h333;
rom[92627] = 12'h444;
rom[92628] = 12'h555;
rom[92629] = 12'h666;
rom[92630] = 12'h777;
rom[92631] = 12'h777;
rom[92632] = 12'h888;
rom[92633] = 12'h888;
rom[92634] = 12'h777;
rom[92635] = 12'h666;
rom[92636] = 12'h555;
rom[92637] = 12'h444;
rom[92638] = 12'h444;
rom[92639] = 12'h333;
rom[92640] = 12'h333;
rom[92641] = 12'h222;
rom[92642] = 12'h222;
rom[92643] = 12'h222;
rom[92644] = 12'h111;
rom[92645] = 12'h111;
rom[92646] = 12'h111;
rom[92647] = 12'h111;
rom[92648] = 12'h111;
rom[92649] = 12'h111;
rom[92650] = 12'h111;
rom[92651] = 12'h111;
rom[92652] = 12'h111;
rom[92653] = 12'h111;
rom[92654] = 12'h111;
rom[92655] = 12'h111;
rom[92656] = 12'h111;
rom[92657] = 12'h111;
rom[92658] = 12'h111;
rom[92659] = 12'h111;
rom[92660] = 12'h111;
rom[92661] = 12'h111;
rom[92662] = 12'h111;
rom[92663] = 12'h111;
rom[92664] = 12'h222;
rom[92665] = 12'h222;
rom[92666] = 12'h222;
rom[92667] = 12'h222;
rom[92668] = 12'h222;
rom[92669] = 12'h333;
rom[92670] = 12'h333;
rom[92671] = 12'h333;
rom[92672] = 12'h444;
rom[92673] = 12'h555;
rom[92674] = 12'h666;
rom[92675] = 12'h888;
rom[92676] = 12'h999;
rom[92677] = 12'h999;
rom[92678] = 12'h888;
rom[92679] = 12'h777;
rom[92680] = 12'h777;
rom[92681] = 12'h777;
rom[92682] = 12'h777;
rom[92683] = 12'h777;
rom[92684] = 12'h777;
rom[92685] = 12'h777;
rom[92686] = 12'h777;
rom[92687] = 12'h777;
rom[92688] = 12'h777;
rom[92689] = 12'h888;
rom[92690] = 12'h999;
rom[92691] = 12'h999;
rom[92692] = 12'h999;
rom[92693] = 12'haaa;
rom[92694] = 12'haaa;
rom[92695] = 12'haaa;
rom[92696] = 12'hddd;
rom[92697] = 12'heee;
rom[92698] = 12'heee;
rom[92699] = 12'hddd;
rom[92700] = 12'hccc;
rom[92701] = 12'hccc;
rom[92702] = 12'hddd;
rom[92703] = 12'hccc;
rom[92704] = 12'hddd;
rom[92705] = 12'hbbb;
rom[92706] = 12'haaa;
rom[92707] = 12'h999;
rom[92708] = 12'h999;
rom[92709] = 12'h999;
rom[92710] = 12'h777;
rom[92711] = 12'h777;
rom[92712] = 12'h555;
rom[92713] = 12'h444;
rom[92714] = 12'h333;
rom[92715] = 12'h333;
rom[92716] = 12'h444;
rom[92717] = 12'h444;
rom[92718] = 12'h444;
rom[92719] = 12'h444;
rom[92720] = 12'h333;
rom[92721] = 12'h333;
rom[92722] = 12'h333;
rom[92723] = 12'h444;
rom[92724] = 12'h444;
rom[92725] = 12'h444;
rom[92726] = 12'h444;
rom[92727] = 12'h333;
rom[92728] = 12'h333;
rom[92729] = 12'h333;
rom[92730] = 12'h333;
rom[92731] = 12'h333;
rom[92732] = 12'h333;
rom[92733] = 12'h222;
rom[92734] = 12'h222;
rom[92735] = 12'h222;
rom[92736] = 12'h222;
rom[92737] = 12'h222;
rom[92738] = 12'h222;
rom[92739] = 12'h222;
rom[92740] = 12'h222;
rom[92741] = 12'h222;
rom[92742] = 12'h222;
rom[92743] = 12'h222;
rom[92744] = 12'h111;
rom[92745] = 12'h111;
rom[92746] = 12'h111;
rom[92747] = 12'h111;
rom[92748] = 12'h222;
rom[92749] = 12'h222;
rom[92750] = 12'h222;
rom[92751] = 12'h222;
rom[92752] = 12'h222;
rom[92753] = 12'h222;
rom[92754] = 12'h333;
rom[92755] = 12'h333;
rom[92756] = 12'h333;
rom[92757] = 12'h333;
rom[92758] = 12'h333;
rom[92759] = 12'h444;
rom[92760] = 12'h555;
rom[92761] = 12'h777;
rom[92762] = 12'h888;
rom[92763] = 12'haaa;
rom[92764] = 12'hddd;
rom[92765] = 12'hfff;
rom[92766] = 12'hfff;
rom[92767] = 12'heee;
rom[92768] = 12'hccc;
rom[92769] = 12'h999;
rom[92770] = 12'h777;
rom[92771] = 12'h555;
rom[92772] = 12'h555;
rom[92773] = 12'h444;
rom[92774] = 12'h333;
rom[92775] = 12'h333;
rom[92776] = 12'h333;
rom[92777] = 12'h333;
rom[92778] = 12'h333;
rom[92779] = 12'h333;
rom[92780] = 12'h333;
rom[92781] = 12'h222;
rom[92782] = 12'h222;
rom[92783] = 12'h222;
rom[92784] = 12'h222;
rom[92785] = 12'h222;
rom[92786] = 12'h222;
rom[92787] = 12'h222;
rom[92788] = 12'h222;
rom[92789] = 12'h222;
rom[92790] = 12'h222;
rom[92791] = 12'h222;
rom[92792] = 12'h111;
rom[92793] = 12'h111;
rom[92794] = 12'h222;
rom[92795] = 12'h222;
rom[92796] = 12'h222;
rom[92797] = 12'h222;
rom[92798] = 12'h222;
rom[92799] = 12'h111;
rom[92800] = 12'hfff;
rom[92801] = 12'hfff;
rom[92802] = 12'hfff;
rom[92803] = 12'hfff;
rom[92804] = 12'hfff;
rom[92805] = 12'hfff;
rom[92806] = 12'hfff;
rom[92807] = 12'hfff;
rom[92808] = 12'hfff;
rom[92809] = 12'hfff;
rom[92810] = 12'hfff;
rom[92811] = 12'hfff;
rom[92812] = 12'hfff;
rom[92813] = 12'hfff;
rom[92814] = 12'hfff;
rom[92815] = 12'hfff;
rom[92816] = 12'hfff;
rom[92817] = 12'hfff;
rom[92818] = 12'hfff;
rom[92819] = 12'hfff;
rom[92820] = 12'hfff;
rom[92821] = 12'hfff;
rom[92822] = 12'hfff;
rom[92823] = 12'hfff;
rom[92824] = 12'hfff;
rom[92825] = 12'hfff;
rom[92826] = 12'hfff;
rom[92827] = 12'hfff;
rom[92828] = 12'hfff;
rom[92829] = 12'hfff;
rom[92830] = 12'hfff;
rom[92831] = 12'hfff;
rom[92832] = 12'hfff;
rom[92833] = 12'hfff;
rom[92834] = 12'hfff;
rom[92835] = 12'hfff;
rom[92836] = 12'hfff;
rom[92837] = 12'hfff;
rom[92838] = 12'hfff;
rom[92839] = 12'hfff;
rom[92840] = 12'hfff;
rom[92841] = 12'hfff;
rom[92842] = 12'hfff;
rom[92843] = 12'hfff;
rom[92844] = 12'hfff;
rom[92845] = 12'hfff;
rom[92846] = 12'hfff;
rom[92847] = 12'hfff;
rom[92848] = 12'hfff;
rom[92849] = 12'hfff;
rom[92850] = 12'hfff;
rom[92851] = 12'hfff;
rom[92852] = 12'hfff;
rom[92853] = 12'hfff;
rom[92854] = 12'hfff;
rom[92855] = 12'hfff;
rom[92856] = 12'hfff;
rom[92857] = 12'hfff;
rom[92858] = 12'hfff;
rom[92859] = 12'hfff;
rom[92860] = 12'hfff;
rom[92861] = 12'hfff;
rom[92862] = 12'hfff;
rom[92863] = 12'hfff;
rom[92864] = 12'hfff;
rom[92865] = 12'hfff;
rom[92866] = 12'hfff;
rom[92867] = 12'hfff;
rom[92868] = 12'hfff;
rom[92869] = 12'hfff;
rom[92870] = 12'hfff;
rom[92871] = 12'hfff;
rom[92872] = 12'hfff;
rom[92873] = 12'hfff;
rom[92874] = 12'hfff;
rom[92875] = 12'hfff;
rom[92876] = 12'hfff;
rom[92877] = 12'hfff;
rom[92878] = 12'hfff;
rom[92879] = 12'hfff;
rom[92880] = 12'hfff;
rom[92881] = 12'hfff;
rom[92882] = 12'hfff;
rom[92883] = 12'hfff;
rom[92884] = 12'hfff;
rom[92885] = 12'hfff;
rom[92886] = 12'hfff;
rom[92887] = 12'hfff;
rom[92888] = 12'hfff;
rom[92889] = 12'hfff;
rom[92890] = 12'hfff;
rom[92891] = 12'hfff;
rom[92892] = 12'hfff;
rom[92893] = 12'hfff;
rom[92894] = 12'hfff;
rom[92895] = 12'hfff;
rom[92896] = 12'hfff;
rom[92897] = 12'hfff;
rom[92898] = 12'hfff;
rom[92899] = 12'hfff;
rom[92900] = 12'hfff;
rom[92901] = 12'hfff;
rom[92902] = 12'hfff;
rom[92903] = 12'hfff;
rom[92904] = 12'hfff;
rom[92905] = 12'hfff;
rom[92906] = 12'hfff;
rom[92907] = 12'hfff;
rom[92908] = 12'hfff;
rom[92909] = 12'hfff;
rom[92910] = 12'hfff;
rom[92911] = 12'hfff;
rom[92912] = 12'hfff;
rom[92913] = 12'hfff;
rom[92914] = 12'hfff;
rom[92915] = 12'hfff;
rom[92916] = 12'hfff;
rom[92917] = 12'hfff;
rom[92918] = 12'hfff;
rom[92919] = 12'hfff;
rom[92920] = 12'hfff;
rom[92921] = 12'hfff;
rom[92922] = 12'hfff;
rom[92923] = 12'hfff;
rom[92924] = 12'hfff;
rom[92925] = 12'hfff;
rom[92926] = 12'hfff;
rom[92927] = 12'hfff;
rom[92928] = 12'hfff;
rom[92929] = 12'hfff;
rom[92930] = 12'hfff;
rom[92931] = 12'hfff;
rom[92932] = 12'hfff;
rom[92933] = 12'hfff;
rom[92934] = 12'heee;
rom[92935] = 12'heee;
rom[92936] = 12'heee;
rom[92937] = 12'heee;
rom[92938] = 12'heee;
rom[92939] = 12'heee;
rom[92940] = 12'heee;
rom[92941] = 12'heee;
rom[92942] = 12'heee;
rom[92943] = 12'heee;
rom[92944] = 12'hddd;
rom[92945] = 12'hddd;
rom[92946] = 12'hddd;
rom[92947] = 12'hddd;
rom[92948] = 12'hddd;
rom[92949] = 12'hccc;
rom[92950] = 12'hbbb;
rom[92951] = 12'hbbb;
rom[92952] = 12'haaa;
rom[92953] = 12'haaa;
rom[92954] = 12'haaa;
rom[92955] = 12'h999;
rom[92956] = 12'h999;
rom[92957] = 12'h999;
rom[92958] = 12'h888;
rom[92959] = 12'h888;
rom[92960] = 12'h888;
rom[92961] = 12'h888;
rom[92962] = 12'h888;
rom[92963] = 12'h888;
rom[92964] = 12'h888;
rom[92965] = 12'h888;
rom[92966] = 12'h888;
rom[92967] = 12'h888;
rom[92968] = 12'h888;
rom[92969] = 12'h888;
rom[92970] = 12'h888;
rom[92971] = 12'h888;
rom[92972] = 12'h888;
rom[92973] = 12'h888;
rom[92974] = 12'h888;
rom[92975] = 12'h888;
rom[92976] = 12'h888;
rom[92977] = 12'h888;
rom[92978] = 12'h888;
rom[92979] = 12'h888;
rom[92980] = 12'h888;
rom[92981] = 12'h888;
rom[92982] = 12'h888;
rom[92983] = 12'h888;
rom[92984] = 12'h888;
rom[92985] = 12'h888;
rom[92986] = 12'h888;
rom[92987] = 12'h888;
rom[92988] = 12'h888;
rom[92989] = 12'h888;
rom[92990] = 12'h888;
rom[92991] = 12'h888;
rom[92992] = 12'h888;
rom[92993] = 12'h888;
rom[92994] = 12'h888;
rom[92995] = 12'h888;
rom[92996] = 12'h888;
rom[92997] = 12'h888;
rom[92998] = 12'h777;
rom[92999] = 12'h777;
rom[93000] = 12'h777;
rom[93001] = 12'h777;
rom[93002] = 12'h777;
rom[93003] = 12'h777;
rom[93004] = 12'h777;
rom[93005] = 12'h777;
rom[93006] = 12'h666;
rom[93007] = 12'h666;
rom[93008] = 12'h666;
rom[93009] = 12'h666;
rom[93010] = 12'h666;
rom[93011] = 12'h555;
rom[93012] = 12'h555;
rom[93013] = 12'h555;
rom[93014] = 12'h555;
rom[93015] = 12'h444;
rom[93016] = 12'h444;
rom[93017] = 12'h333;
rom[93018] = 12'h333;
rom[93019] = 12'h333;
rom[93020] = 12'h333;
rom[93021] = 12'h333;
rom[93022] = 12'h333;
rom[93023] = 12'h333;
rom[93024] = 12'h222;
rom[93025] = 12'h333;
rom[93026] = 12'h333;
rom[93027] = 12'h444;
rom[93028] = 12'h444;
rom[93029] = 12'h555;
rom[93030] = 12'h666;
rom[93031] = 12'h777;
rom[93032] = 12'h888;
rom[93033] = 12'h888;
rom[93034] = 12'h888;
rom[93035] = 12'h888;
rom[93036] = 12'h777;
rom[93037] = 12'h666;
rom[93038] = 12'h555;
rom[93039] = 12'h444;
rom[93040] = 12'h333;
rom[93041] = 12'h333;
rom[93042] = 12'h333;
rom[93043] = 12'h222;
rom[93044] = 12'h222;
rom[93045] = 12'h222;
rom[93046] = 12'h222;
rom[93047] = 12'h111;
rom[93048] = 12'h222;
rom[93049] = 12'h111;
rom[93050] = 12'h111;
rom[93051] = 12'h111;
rom[93052] = 12'h111;
rom[93053] = 12'h111;
rom[93054] = 12'h111;
rom[93055] = 12'h111;
rom[93056] = 12'h111;
rom[93057] = 12'h111;
rom[93058] = 12'h111;
rom[93059] = 12'h111;
rom[93060] = 12'h111;
rom[93061] = 12'h111;
rom[93062] = 12'h222;
rom[93063] = 12'h222;
rom[93064] = 12'h222;
rom[93065] = 12'h222;
rom[93066] = 12'h222;
rom[93067] = 12'h222;
rom[93068] = 12'h333;
rom[93069] = 12'h333;
rom[93070] = 12'h444;
rom[93071] = 12'h555;
rom[93072] = 12'h666;
rom[93073] = 12'h777;
rom[93074] = 12'h888;
rom[93075] = 12'h888;
rom[93076] = 12'h999;
rom[93077] = 12'h999;
rom[93078] = 12'h888;
rom[93079] = 12'h888;
rom[93080] = 12'h777;
rom[93081] = 12'h888;
rom[93082] = 12'h888;
rom[93083] = 12'h777;
rom[93084] = 12'h777;
rom[93085] = 12'h888;
rom[93086] = 12'h888;
rom[93087] = 12'h888;
rom[93088] = 12'h888;
rom[93089] = 12'h888;
rom[93090] = 12'h999;
rom[93091] = 12'h999;
rom[93092] = 12'h999;
rom[93093] = 12'haaa;
rom[93094] = 12'hbbb;
rom[93095] = 12'hccc;
rom[93096] = 12'hddd;
rom[93097] = 12'heee;
rom[93098] = 12'heee;
rom[93099] = 12'hddd;
rom[93100] = 12'hccc;
rom[93101] = 12'hddd;
rom[93102] = 12'hddd;
rom[93103] = 12'hddd;
rom[93104] = 12'hddd;
rom[93105] = 12'hddd;
rom[93106] = 12'hccc;
rom[93107] = 12'hbbb;
rom[93108] = 12'haaa;
rom[93109] = 12'haaa;
rom[93110] = 12'h999;
rom[93111] = 12'h888;
rom[93112] = 12'h666;
rom[93113] = 12'h555;
rom[93114] = 12'h444;
rom[93115] = 12'h444;
rom[93116] = 12'h444;
rom[93117] = 12'h444;
rom[93118] = 12'h444;
rom[93119] = 12'h444;
rom[93120] = 12'h333;
rom[93121] = 12'h333;
rom[93122] = 12'h333;
rom[93123] = 12'h333;
rom[93124] = 12'h333;
rom[93125] = 12'h444;
rom[93126] = 12'h333;
rom[93127] = 12'h333;
rom[93128] = 12'h333;
rom[93129] = 12'h444;
rom[93130] = 12'h333;
rom[93131] = 12'h333;
rom[93132] = 12'h222;
rom[93133] = 12'h222;
rom[93134] = 12'h222;
rom[93135] = 12'h222;
rom[93136] = 12'h222;
rom[93137] = 12'h222;
rom[93138] = 12'h222;
rom[93139] = 12'h222;
rom[93140] = 12'h111;
rom[93141] = 12'h111;
rom[93142] = 12'h111;
rom[93143] = 12'h111;
rom[93144] = 12'h111;
rom[93145] = 12'h111;
rom[93146] = 12'h111;
rom[93147] = 12'h111;
rom[93148] = 12'h111;
rom[93149] = 12'h111;
rom[93150] = 12'h111;
rom[93151] = 12'h111;
rom[93152] = 12'h222;
rom[93153] = 12'h222;
rom[93154] = 12'h222;
rom[93155] = 12'h222;
rom[93156] = 12'h333;
rom[93157] = 12'h333;
rom[93158] = 12'h333;
rom[93159] = 12'h333;
rom[93160] = 12'h444;
rom[93161] = 12'h444;
rom[93162] = 12'h555;
rom[93163] = 12'h666;
rom[93164] = 12'h888;
rom[93165] = 12'hbbb;
rom[93166] = 12'hddd;
rom[93167] = 12'heee;
rom[93168] = 12'heee;
rom[93169] = 12'heee;
rom[93170] = 12'hbbb;
rom[93171] = 12'h888;
rom[93172] = 12'h666;
rom[93173] = 12'h555;
rom[93174] = 12'h444;
rom[93175] = 12'h333;
rom[93176] = 12'h333;
rom[93177] = 12'h333;
rom[93178] = 12'h333;
rom[93179] = 12'h333;
rom[93180] = 12'h333;
rom[93181] = 12'h222;
rom[93182] = 12'h222;
rom[93183] = 12'h222;
rom[93184] = 12'h222;
rom[93185] = 12'h222;
rom[93186] = 12'h222;
rom[93187] = 12'h222;
rom[93188] = 12'h222;
rom[93189] = 12'h222;
rom[93190] = 12'h111;
rom[93191] = 12'h111;
rom[93192] = 12'h111;
rom[93193] = 12'h111;
rom[93194] = 12'h111;
rom[93195] = 12'h111;
rom[93196] = 12'h111;
rom[93197] = 12'h111;
rom[93198] = 12'h111;
rom[93199] = 12'h111;
rom[93200] = 12'hfff;
rom[93201] = 12'hfff;
rom[93202] = 12'hfff;
rom[93203] = 12'hfff;
rom[93204] = 12'hfff;
rom[93205] = 12'hfff;
rom[93206] = 12'hfff;
rom[93207] = 12'hfff;
rom[93208] = 12'hfff;
rom[93209] = 12'hfff;
rom[93210] = 12'hfff;
rom[93211] = 12'hfff;
rom[93212] = 12'hfff;
rom[93213] = 12'hfff;
rom[93214] = 12'hfff;
rom[93215] = 12'hfff;
rom[93216] = 12'hfff;
rom[93217] = 12'hfff;
rom[93218] = 12'hfff;
rom[93219] = 12'hfff;
rom[93220] = 12'hfff;
rom[93221] = 12'hfff;
rom[93222] = 12'hfff;
rom[93223] = 12'hfff;
rom[93224] = 12'hfff;
rom[93225] = 12'hfff;
rom[93226] = 12'hfff;
rom[93227] = 12'hfff;
rom[93228] = 12'hfff;
rom[93229] = 12'hfff;
rom[93230] = 12'hfff;
rom[93231] = 12'hfff;
rom[93232] = 12'hfff;
rom[93233] = 12'hfff;
rom[93234] = 12'hfff;
rom[93235] = 12'hfff;
rom[93236] = 12'hfff;
rom[93237] = 12'hfff;
rom[93238] = 12'hfff;
rom[93239] = 12'hfff;
rom[93240] = 12'hfff;
rom[93241] = 12'hfff;
rom[93242] = 12'hfff;
rom[93243] = 12'hfff;
rom[93244] = 12'hfff;
rom[93245] = 12'hfff;
rom[93246] = 12'hfff;
rom[93247] = 12'hfff;
rom[93248] = 12'hfff;
rom[93249] = 12'hfff;
rom[93250] = 12'hfff;
rom[93251] = 12'hfff;
rom[93252] = 12'hfff;
rom[93253] = 12'hfff;
rom[93254] = 12'hfff;
rom[93255] = 12'hfff;
rom[93256] = 12'hfff;
rom[93257] = 12'hfff;
rom[93258] = 12'hfff;
rom[93259] = 12'hfff;
rom[93260] = 12'hfff;
rom[93261] = 12'hfff;
rom[93262] = 12'hfff;
rom[93263] = 12'hfff;
rom[93264] = 12'hfff;
rom[93265] = 12'hfff;
rom[93266] = 12'hfff;
rom[93267] = 12'hfff;
rom[93268] = 12'hfff;
rom[93269] = 12'hfff;
rom[93270] = 12'hfff;
rom[93271] = 12'hfff;
rom[93272] = 12'hfff;
rom[93273] = 12'hfff;
rom[93274] = 12'hfff;
rom[93275] = 12'hfff;
rom[93276] = 12'hfff;
rom[93277] = 12'hfff;
rom[93278] = 12'hfff;
rom[93279] = 12'hfff;
rom[93280] = 12'hfff;
rom[93281] = 12'hfff;
rom[93282] = 12'hfff;
rom[93283] = 12'hfff;
rom[93284] = 12'hfff;
rom[93285] = 12'hfff;
rom[93286] = 12'hfff;
rom[93287] = 12'hfff;
rom[93288] = 12'hfff;
rom[93289] = 12'hfff;
rom[93290] = 12'hfff;
rom[93291] = 12'hfff;
rom[93292] = 12'hfff;
rom[93293] = 12'hfff;
rom[93294] = 12'hfff;
rom[93295] = 12'hfff;
rom[93296] = 12'hfff;
rom[93297] = 12'hfff;
rom[93298] = 12'hfff;
rom[93299] = 12'hfff;
rom[93300] = 12'hfff;
rom[93301] = 12'hfff;
rom[93302] = 12'hfff;
rom[93303] = 12'hfff;
rom[93304] = 12'hfff;
rom[93305] = 12'hfff;
rom[93306] = 12'hfff;
rom[93307] = 12'hfff;
rom[93308] = 12'hfff;
rom[93309] = 12'hfff;
rom[93310] = 12'hfff;
rom[93311] = 12'hfff;
rom[93312] = 12'hfff;
rom[93313] = 12'hfff;
rom[93314] = 12'hfff;
rom[93315] = 12'hfff;
rom[93316] = 12'hfff;
rom[93317] = 12'hfff;
rom[93318] = 12'hfff;
rom[93319] = 12'hfff;
rom[93320] = 12'hfff;
rom[93321] = 12'hfff;
rom[93322] = 12'hfff;
rom[93323] = 12'hfff;
rom[93324] = 12'hfff;
rom[93325] = 12'hfff;
rom[93326] = 12'hfff;
rom[93327] = 12'hfff;
rom[93328] = 12'hfff;
rom[93329] = 12'hfff;
rom[93330] = 12'hfff;
rom[93331] = 12'hfff;
rom[93332] = 12'hfff;
rom[93333] = 12'hfff;
rom[93334] = 12'heee;
rom[93335] = 12'heee;
rom[93336] = 12'heee;
rom[93337] = 12'heee;
rom[93338] = 12'hddd;
rom[93339] = 12'hddd;
rom[93340] = 12'hddd;
rom[93341] = 12'hddd;
rom[93342] = 12'hddd;
rom[93343] = 12'hddd;
rom[93344] = 12'heee;
rom[93345] = 12'heee;
rom[93346] = 12'heee;
rom[93347] = 12'heee;
rom[93348] = 12'heee;
rom[93349] = 12'hddd;
rom[93350] = 12'hddd;
rom[93351] = 12'hddd;
rom[93352] = 12'hbbb;
rom[93353] = 12'hbbb;
rom[93354] = 12'hbbb;
rom[93355] = 12'haaa;
rom[93356] = 12'haaa;
rom[93357] = 12'haaa;
rom[93358] = 12'h999;
rom[93359] = 12'h999;
rom[93360] = 12'h888;
rom[93361] = 12'h888;
rom[93362] = 12'h888;
rom[93363] = 12'h888;
rom[93364] = 12'h888;
rom[93365] = 12'h888;
rom[93366] = 12'h888;
rom[93367] = 12'h888;
rom[93368] = 12'h888;
rom[93369] = 12'h888;
rom[93370] = 12'h888;
rom[93371] = 12'h888;
rom[93372] = 12'h888;
rom[93373] = 12'h888;
rom[93374] = 12'h888;
rom[93375] = 12'h888;
rom[93376] = 12'h888;
rom[93377] = 12'h888;
rom[93378] = 12'h888;
rom[93379] = 12'h999;
rom[93380] = 12'h888;
rom[93381] = 12'h888;
rom[93382] = 12'h888;
rom[93383] = 12'h888;
rom[93384] = 12'h888;
rom[93385] = 12'h888;
rom[93386] = 12'h888;
rom[93387] = 12'h888;
rom[93388] = 12'h888;
rom[93389] = 12'h888;
rom[93390] = 12'h888;
rom[93391] = 12'h888;
rom[93392] = 12'h888;
rom[93393] = 12'h888;
rom[93394] = 12'h888;
rom[93395] = 12'h888;
rom[93396] = 12'h888;
rom[93397] = 12'h888;
rom[93398] = 12'h888;
rom[93399] = 12'h888;
rom[93400] = 12'h777;
rom[93401] = 12'h777;
rom[93402] = 12'h777;
rom[93403] = 12'h777;
rom[93404] = 12'h777;
rom[93405] = 12'h777;
rom[93406] = 12'h777;
rom[93407] = 12'h777;
rom[93408] = 12'h666;
rom[93409] = 12'h666;
rom[93410] = 12'h666;
rom[93411] = 12'h666;
rom[93412] = 12'h555;
rom[93413] = 12'h555;
rom[93414] = 12'h555;
rom[93415] = 12'h444;
rom[93416] = 12'h444;
rom[93417] = 12'h444;
rom[93418] = 12'h333;
rom[93419] = 12'h333;
rom[93420] = 12'h333;
rom[93421] = 12'h333;
rom[93422] = 12'h333;
rom[93423] = 12'h333;
rom[93424] = 12'h222;
rom[93425] = 12'h333;
rom[93426] = 12'h444;
rom[93427] = 12'h444;
rom[93428] = 12'h444;
rom[93429] = 12'h555;
rom[93430] = 12'h666;
rom[93431] = 12'h777;
rom[93432] = 12'h777;
rom[93433] = 12'h777;
rom[93434] = 12'h888;
rom[93435] = 12'h888;
rom[93436] = 12'h777;
rom[93437] = 12'h777;
rom[93438] = 12'h666;
rom[93439] = 12'h555;
rom[93440] = 12'h444;
rom[93441] = 12'h444;
rom[93442] = 12'h333;
rom[93443] = 12'h222;
rom[93444] = 12'h222;
rom[93445] = 12'h222;
rom[93446] = 12'h222;
rom[93447] = 12'h222;
rom[93448] = 12'h222;
rom[93449] = 12'h111;
rom[93450] = 12'h111;
rom[93451] = 12'h111;
rom[93452] = 12'h111;
rom[93453] = 12'h111;
rom[93454] = 12'h111;
rom[93455] = 12'h111;
rom[93456] = 12'h111;
rom[93457] = 12'h111;
rom[93458] = 12'h111;
rom[93459] = 12'h111;
rom[93460] = 12'h111;
rom[93461] = 12'h111;
rom[93462] = 12'h222;
rom[93463] = 12'h222;
rom[93464] = 12'h222;
rom[93465] = 12'h222;
rom[93466] = 12'h222;
rom[93467] = 12'h333;
rom[93468] = 12'h333;
rom[93469] = 12'h444;
rom[93470] = 12'h555;
rom[93471] = 12'h666;
rom[93472] = 12'h777;
rom[93473] = 12'h888;
rom[93474] = 12'h888;
rom[93475] = 12'h888;
rom[93476] = 12'h888;
rom[93477] = 12'h888;
rom[93478] = 12'h777;
rom[93479] = 12'h777;
rom[93480] = 12'h777;
rom[93481] = 12'h777;
rom[93482] = 12'h888;
rom[93483] = 12'h888;
rom[93484] = 12'h888;
rom[93485] = 12'h888;
rom[93486] = 12'h888;
rom[93487] = 12'h999;
rom[93488] = 12'h999;
rom[93489] = 12'h999;
rom[93490] = 12'h999;
rom[93491] = 12'h999;
rom[93492] = 12'h999;
rom[93493] = 12'haaa;
rom[93494] = 12'hbbb;
rom[93495] = 12'hddd;
rom[93496] = 12'heee;
rom[93497] = 12'heee;
rom[93498] = 12'hddd;
rom[93499] = 12'hccc;
rom[93500] = 12'hccc;
rom[93501] = 12'hddd;
rom[93502] = 12'hddd;
rom[93503] = 12'hddd;
rom[93504] = 12'heee;
rom[93505] = 12'heee;
rom[93506] = 12'heee;
rom[93507] = 12'hddd;
rom[93508] = 12'hccc;
rom[93509] = 12'hbbb;
rom[93510] = 12'haaa;
rom[93511] = 12'h999;
rom[93512] = 12'h777;
rom[93513] = 12'h666;
rom[93514] = 12'h555;
rom[93515] = 12'h444;
rom[93516] = 12'h444;
rom[93517] = 12'h444;
rom[93518] = 12'h444;
rom[93519] = 12'h333;
rom[93520] = 12'h444;
rom[93521] = 12'h444;
rom[93522] = 12'h333;
rom[93523] = 12'h333;
rom[93524] = 12'h444;
rom[93525] = 12'h444;
rom[93526] = 12'h444;
rom[93527] = 12'h444;
rom[93528] = 12'h333;
rom[93529] = 12'h333;
rom[93530] = 12'h444;
rom[93531] = 12'h333;
rom[93532] = 12'h333;
rom[93533] = 12'h333;
rom[93534] = 12'h222;
rom[93535] = 12'h222;
rom[93536] = 12'h222;
rom[93537] = 12'h222;
rom[93538] = 12'h222;
rom[93539] = 12'h222;
rom[93540] = 12'h111;
rom[93541] = 12'h111;
rom[93542] = 12'h111;
rom[93543] = 12'h111;
rom[93544] = 12'h111;
rom[93545] = 12'h111;
rom[93546] = 12'h111;
rom[93547] = 12'h111;
rom[93548] = 12'h111;
rom[93549] = 12'h111;
rom[93550] = 12'h111;
rom[93551] = 12'h222;
rom[93552] = 12'h111;
rom[93553] = 12'h222;
rom[93554] = 12'h222;
rom[93555] = 12'h222;
rom[93556] = 12'h222;
rom[93557] = 12'h222;
rom[93558] = 12'h333;
rom[93559] = 12'h333;
rom[93560] = 12'h333;
rom[93561] = 12'h333;
rom[93562] = 12'h444;
rom[93563] = 12'h555;
rom[93564] = 12'h666;
rom[93565] = 12'h777;
rom[93566] = 12'h999;
rom[93567] = 12'haaa;
rom[93568] = 12'heee;
rom[93569] = 12'heee;
rom[93570] = 12'heee;
rom[93571] = 12'hccc;
rom[93572] = 12'haaa;
rom[93573] = 12'h888;
rom[93574] = 12'h666;
rom[93575] = 12'h444;
rom[93576] = 12'h333;
rom[93577] = 12'h333;
rom[93578] = 12'h333;
rom[93579] = 12'h333;
rom[93580] = 12'h333;
rom[93581] = 12'h333;
rom[93582] = 12'h222;
rom[93583] = 12'h222;
rom[93584] = 12'h222;
rom[93585] = 12'h222;
rom[93586] = 12'h222;
rom[93587] = 12'h222;
rom[93588] = 12'h222;
rom[93589] = 12'h222;
rom[93590] = 12'h222;
rom[93591] = 12'h111;
rom[93592] = 12'h111;
rom[93593] = 12'h111;
rom[93594] = 12'h111;
rom[93595] = 12'h111;
rom[93596] = 12'h111;
rom[93597] = 12'h111;
rom[93598] = 12'h111;
rom[93599] = 12'h111;
rom[93600] = 12'hfff;
rom[93601] = 12'hfff;
rom[93602] = 12'hfff;
rom[93603] = 12'hfff;
rom[93604] = 12'hfff;
rom[93605] = 12'hfff;
rom[93606] = 12'hfff;
rom[93607] = 12'hfff;
rom[93608] = 12'hfff;
rom[93609] = 12'hfff;
rom[93610] = 12'hfff;
rom[93611] = 12'hfff;
rom[93612] = 12'hfff;
rom[93613] = 12'hfff;
rom[93614] = 12'hfff;
rom[93615] = 12'hfff;
rom[93616] = 12'hfff;
rom[93617] = 12'hfff;
rom[93618] = 12'hfff;
rom[93619] = 12'hfff;
rom[93620] = 12'hfff;
rom[93621] = 12'hfff;
rom[93622] = 12'hfff;
rom[93623] = 12'hfff;
rom[93624] = 12'hfff;
rom[93625] = 12'hfff;
rom[93626] = 12'hfff;
rom[93627] = 12'hfff;
rom[93628] = 12'hfff;
rom[93629] = 12'hfff;
rom[93630] = 12'hfff;
rom[93631] = 12'hfff;
rom[93632] = 12'hfff;
rom[93633] = 12'hfff;
rom[93634] = 12'hfff;
rom[93635] = 12'hfff;
rom[93636] = 12'hfff;
rom[93637] = 12'hfff;
rom[93638] = 12'hfff;
rom[93639] = 12'hfff;
rom[93640] = 12'hfff;
rom[93641] = 12'hfff;
rom[93642] = 12'hfff;
rom[93643] = 12'hfff;
rom[93644] = 12'hfff;
rom[93645] = 12'hfff;
rom[93646] = 12'hfff;
rom[93647] = 12'hfff;
rom[93648] = 12'hfff;
rom[93649] = 12'hfff;
rom[93650] = 12'hfff;
rom[93651] = 12'hfff;
rom[93652] = 12'hfff;
rom[93653] = 12'hfff;
rom[93654] = 12'hfff;
rom[93655] = 12'hfff;
rom[93656] = 12'hfff;
rom[93657] = 12'hfff;
rom[93658] = 12'hfff;
rom[93659] = 12'hfff;
rom[93660] = 12'hfff;
rom[93661] = 12'hfff;
rom[93662] = 12'hfff;
rom[93663] = 12'hfff;
rom[93664] = 12'hfff;
rom[93665] = 12'hfff;
rom[93666] = 12'hfff;
rom[93667] = 12'hfff;
rom[93668] = 12'hfff;
rom[93669] = 12'hfff;
rom[93670] = 12'hfff;
rom[93671] = 12'hfff;
rom[93672] = 12'hfff;
rom[93673] = 12'hfff;
rom[93674] = 12'hfff;
rom[93675] = 12'hfff;
rom[93676] = 12'hfff;
rom[93677] = 12'hfff;
rom[93678] = 12'hfff;
rom[93679] = 12'hfff;
rom[93680] = 12'hfff;
rom[93681] = 12'hfff;
rom[93682] = 12'hfff;
rom[93683] = 12'hfff;
rom[93684] = 12'hfff;
rom[93685] = 12'hfff;
rom[93686] = 12'hfff;
rom[93687] = 12'hfff;
rom[93688] = 12'hfff;
rom[93689] = 12'hfff;
rom[93690] = 12'hfff;
rom[93691] = 12'hfff;
rom[93692] = 12'hfff;
rom[93693] = 12'hfff;
rom[93694] = 12'hfff;
rom[93695] = 12'hfff;
rom[93696] = 12'hfff;
rom[93697] = 12'hfff;
rom[93698] = 12'hfff;
rom[93699] = 12'hfff;
rom[93700] = 12'hfff;
rom[93701] = 12'hfff;
rom[93702] = 12'hfff;
rom[93703] = 12'hfff;
rom[93704] = 12'hfff;
rom[93705] = 12'hfff;
rom[93706] = 12'hfff;
rom[93707] = 12'hfff;
rom[93708] = 12'hfff;
rom[93709] = 12'hfff;
rom[93710] = 12'hfff;
rom[93711] = 12'hfff;
rom[93712] = 12'hfff;
rom[93713] = 12'hfff;
rom[93714] = 12'hfff;
rom[93715] = 12'hfff;
rom[93716] = 12'hfff;
rom[93717] = 12'hfff;
rom[93718] = 12'hfff;
rom[93719] = 12'hfff;
rom[93720] = 12'hfff;
rom[93721] = 12'hfff;
rom[93722] = 12'hfff;
rom[93723] = 12'hfff;
rom[93724] = 12'hfff;
rom[93725] = 12'hfff;
rom[93726] = 12'hfff;
rom[93727] = 12'hfff;
rom[93728] = 12'hfff;
rom[93729] = 12'hfff;
rom[93730] = 12'hfff;
rom[93731] = 12'hfff;
rom[93732] = 12'hfff;
rom[93733] = 12'hfff;
rom[93734] = 12'hfff;
rom[93735] = 12'heee;
rom[93736] = 12'heee;
rom[93737] = 12'heee;
rom[93738] = 12'hddd;
rom[93739] = 12'hddd;
rom[93740] = 12'hddd;
rom[93741] = 12'hddd;
rom[93742] = 12'hddd;
rom[93743] = 12'hddd;
rom[93744] = 12'hddd;
rom[93745] = 12'hddd;
rom[93746] = 12'hddd;
rom[93747] = 12'hddd;
rom[93748] = 12'hddd;
rom[93749] = 12'heee;
rom[93750] = 12'hddd;
rom[93751] = 12'hddd;
rom[93752] = 12'hccc;
rom[93753] = 12'hccc;
rom[93754] = 12'hccc;
rom[93755] = 12'hbbb;
rom[93756] = 12'hbbb;
rom[93757] = 12'hbbb;
rom[93758] = 12'haaa;
rom[93759] = 12'haaa;
rom[93760] = 12'h999;
rom[93761] = 12'h999;
rom[93762] = 12'h999;
rom[93763] = 12'h999;
rom[93764] = 12'h999;
rom[93765] = 12'h999;
rom[93766] = 12'h888;
rom[93767] = 12'h888;
rom[93768] = 12'h888;
rom[93769] = 12'h888;
rom[93770] = 12'h888;
rom[93771] = 12'h888;
rom[93772] = 12'h888;
rom[93773] = 12'h888;
rom[93774] = 12'h888;
rom[93775] = 12'h888;
rom[93776] = 12'h888;
rom[93777] = 12'h999;
rom[93778] = 12'h999;
rom[93779] = 12'h999;
rom[93780] = 12'h999;
rom[93781] = 12'h999;
rom[93782] = 12'h888;
rom[93783] = 12'h888;
rom[93784] = 12'h888;
rom[93785] = 12'h888;
rom[93786] = 12'h888;
rom[93787] = 12'h888;
rom[93788] = 12'h888;
rom[93789] = 12'h888;
rom[93790] = 12'h888;
rom[93791] = 12'h888;
rom[93792] = 12'h888;
rom[93793] = 12'h888;
rom[93794] = 12'h888;
rom[93795] = 12'h888;
rom[93796] = 12'h888;
rom[93797] = 12'h888;
rom[93798] = 12'h888;
rom[93799] = 12'h888;
rom[93800] = 12'h888;
rom[93801] = 12'h888;
rom[93802] = 12'h888;
rom[93803] = 12'h888;
rom[93804] = 12'h777;
rom[93805] = 12'h777;
rom[93806] = 12'h777;
rom[93807] = 12'h777;
rom[93808] = 12'h777;
rom[93809] = 12'h777;
rom[93810] = 12'h666;
rom[93811] = 12'h666;
rom[93812] = 12'h666;
rom[93813] = 12'h555;
rom[93814] = 12'h555;
rom[93815] = 12'h555;
rom[93816] = 12'h444;
rom[93817] = 12'h444;
rom[93818] = 12'h444;
rom[93819] = 12'h444;
rom[93820] = 12'h444;
rom[93821] = 12'h333;
rom[93822] = 12'h333;
rom[93823] = 12'h333;
rom[93824] = 12'h333;
rom[93825] = 12'h333;
rom[93826] = 12'h444;
rom[93827] = 12'h444;
rom[93828] = 12'h555;
rom[93829] = 12'h555;
rom[93830] = 12'h666;
rom[93831] = 12'h777;
rom[93832] = 12'h777;
rom[93833] = 12'h777;
rom[93834] = 12'h888;
rom[93835] = 12'h888;
rom[93836] = 12'h888;
rom[93837] = 12'h777;
rom[93838] = 12'h777;
rom[93839] = 12'h666;
rom[93840] = 12'h555;
rom[93841] = 12'h555;
rom[93842] = 12'h444;
rom[93843] = 12'h333;
rom[93844] = 12'h222;
rom[93845] = 12'h222;
rom[93846] = 12'h222;
rom[93847] = 12'h222;
rom[93848] = 12'h222;
rom[93849] = 12'h222;
rom[93850] = 12'h222;
rom[93851] = 12'h222;
rom[93852] = 12'h222;
rom[93853] = 12'h222;
rom[93854] = 12'h222;
rom[93855] = 12'h222;
rom[93856] = 12'h222;
rom[93857] = 12'h222;
rom[93858] = 12'h222;
rom[93859] = 12'h222;
rom[93860] = 12'h222;
rom[93861] = 12'h222;
rom[93862] = 12'h222;
rom[93863] = 12'h222;
rom[93864] = 12'h333;
rom[93865] = 12'h333;
rom[93866] = 12'h333;
rom[93867] = 12'h444;
rom[93868] = 12'h555;
rom[93869] = 12'h666;
rom[93870] = 12'h777;
rom[93871] = 12'h888;
rom[93872] = 12'h999;
rom[93873] = 12'h999;
rom[93874] = 12'h888;
rom[93875] = 12'h888;
rom[93876] = 12'h888;
rom[93877] = 12'h888;
rom[93878] = 12'h777;
rom[93879] = 12'h777;
rom[93880] = 12'h777;
rom[93881] = 12'h888;
rom[93882] = 12'h888;
rom[93883] = 12'h888;
rom[93884] = 12'h888;
rom[93885] = 12'h999;
rom[93886] = 12'h999;
rom[93887] = 12'h999;
rom[93888] = 12'h999;
rom[93889] = 12'h999;
rom[93890] = 12'haaa;
rom[93891] = 12'haaa;
rom[93892] = 12'haaa;
rom[93893] = 12'haaa;
rom[93894] = 12'hccc;
rom[93895] = 12'heee;
rom[93896] = 12'hfff;
rom[93897] = 12'hddd;
rom[93898] = 12'hccc;
rom[93899] = 12'hccc;
rom[93900] = 12'hddd;
rom[93901] = 12'hddd;
rom[93902] = 12'hddd;
rom[93903] = 12'heee;
rom[93904] = 12'heee;
rom[93905] = 12'hfff;
rom[93906] = 12'hfff;
rom[93907] = 12'hfff;
rom[93908] = 12'heee;
rom[93909] = 12'hddd;
rom[93910] = 12'hccc;
rom[93911] = 12'hbbb;
rom[93912] = 12'h999;
rom[93913] = 12'h888;
rom[93914] = 12'h666;
rom[93915] = 12'h555;
rom[93916] = 12'h444;
rom[93917] = 12'h444;
rom[93918] = 12'h444;
rom[93919] = 12'h444;
rom[93920] = 12'h444;
rom[93921] = 12'h444;
rom[93922] = 12'h444;
rom[93923] = 12'h333;
rom[93924] = 12'h333;
rom[93925] = 12'h333;
rom[93926] = 12'h333;
rom[93927] = 12'h333;
rom[93928] = 12'h333;
rom[93929] = 12'h333;
rom[93930] = 12'h444;
rom[93931] = 12'h444;
rom[93932] = 12'h444;
rom[93933] = 12'h333;
rom[93934] = 12'h222;
rom[93935] = 12'h222;
rom[93936] = 12'h222;
rom[93937] = 12'h222;
rom[93938] = 12'h111;
rom[93939] = 12'h111;
rom[93940] = 12'h111;
rom[93941] = 12'h111;
rom[93942] = 12'h111;
rom[93943] = 12'h111;
rom[93944] = 12'h111;
rom[93945] = 12'h111;
rom[93946] = 12'h111;
rom[93947] = 12'h111;
rom[93948] = 12'h111;
rom[93949] = 12'h111;
rom[93950] = 12'h111;
rom[93951] = 12'h111;
rom[93952] = 12'h111;
rom[93953] = 12'h111;
rom[93954] = 12'h222;
rom[93955] = 12'h222;
rom[93956] = 12'h222;
rom[93957] = 12'h222;
rom[93958] = 12'h222;
rom[93959] = 12'h222;
rom[93960] = 12'h222;
rom[93961] = 12'h333;
rom[93962] = 12'h333;
rom[93963] = 12'h333;
rom[93964] = 12'h444;
rom[93965] = 12'h444;
rom[93966] = 12'h666;
rom[93967] = 12'h777;
rom[93968] = 12'haaa;
rom[93969] = 12'hbbb;
rom[93970] = 12'hddd;
rom[93971] = 12'heee;
rom[93972] = 12'hddd;
rom[93973] = 12'hccc;
rom[93974] = 12'haaa;
rom[93975] = 12'h888;
rom[93976] = 12'h555;
rom[93977] = 12'h444;
rom[93978] = 12'h333;
rom[93979] = 12'h333;
rom[93980] = 12'h333;
rom[93981] = 12'h333;
rom[93982] = 12'h222;
rom[93983] = 12'h222;
rom[93984] = 12'h222;
rom[93985] = 12'h222;
rom[93986] = 12'h222;
rom[93987] = 12'h222;
rom[93988] = 12'h222;
rom[93989] = 12'h222;
rom[93990] = 12'h111;
rom[93991] = 12'h111;
rom[93992] = 12'h111;
rom[93993] = 12'h111;
rom[93994] = 12'h111;
rom[93995] = 12'h111;
rom[93996] = 12'h111;
rom[93997] = 12'h111;
rom[93998] = 12'h111;
rom[93999] = 12'h111;
rom[94000] = 12'hfff;
rom[94001] = 12'hfff;
rom[94002] = 12'hfff;
rom[94003] = 12'hfff;
rom[94004] = 12'hfff;
rom[94005] = 12'hfff;
rom[94006] = 12'hfff;
rom[94007] = 12'hfff;
rom[94008] = 12'hfff;
rom[94009] = 12'hfff;
rom[94010] = 12'hfff;
rom[94011] = 12'hfff;
rom[94012] = 12'hfff;
rom[94013] = 12'hfff;
rom[94014] = 12'hfff;
rom[94015] = 12'hfff;
rom[94016] = 12'hfff;
rom[94017] = 12'hfff;
rom[94018] = 12'hfff;
rom[94019] = 12'hfff;
rom[94020] = 12'hfff;
rom[94021] = 12'hfff;
rom[94022] = 12'hfff;
rom[94023] = 12'hfff;
rom[94024] = 12'hfff;
rom[94025] = 12'hfff;
rom[94026] = 12'hfff;
rom[94027] = 12'hfff;
rom[94028] = 12'hfff;
rom[94029] = 12'hfff;
rom[94030] = 12'hfff;
rom[94031] = 12'hfff;
rom[94032] = 12'hfff;
rom[94033] = 12'hfff;
rom[94034] = 12'hfff;
rom[94035] = 12'hfff;
rom[94036] = 12'hfff;
rom[94037] = 12'hfff;
rom[94038] = 12'hfff;
rom[94039] = 12'hfff;
rom[94040] = 12'hfff;
rom[94041] = 12'hfff;
rom[94042] = 12'hfff;
rom[94043] = 12'hfff;
rom[94044] = 12'hfff;
rom[94045] = 12'hfff;
rom[94046] = 12'hfff;
rom[94047] = 12'hfff;
rom[94048] = 12'hfff;
rom[94049] = 12'hfff;
rom[94050] = 12'hfff;
rom[94051] = 12'hfff;
rom[94052] = 12'hfff;
rom[94053] = 12'hfff;
rom[94054] = 12'hfff;
rom[94055] = 12'hfff;
rom[94056] = 12'hfff;
rom[94057] = 12'hfff;
rom[94058] = 12'hfff;
rom[94059] = 12'hfff;
rom[94060] = 12'hfff;
rom[94061] = 12'hfff;
rom[94062] = 12'hfff;
rom[94063] = 12'hfff;
rom[94064] = 12'hfff;
rom[94065] = 12'hfff;
rom[94066] = 12'hfff;
rom[94067] = 12'hfff;
rom[94068] = 12'hfff;
rom[94069] = 12'hfff;
rom[94070] = 12'hfff;
rom[94071] = 12'hfff;
rom[94072] = 12'hfff;
rom[94073] = 12'hfff;
rom[94074] = 12'hfff;
rom[94075] = 12'hfff;
rom[94076] = 12'hfff;
rom[94077] = 12'hfff;
rom[94078] = 12'hfff;
rom[94079] = 12'hfff;
rom[94080] = 12'hfff;
rom[94081] = 12'hfff;
rom[94082] = 12'hfff;
rom[94083] = 12'hfff;
rom[94084] = 12'hfff;
rom[94085] = 12'hfff;
rom[94086] = 12'hfff;
rom[94087] = 12'hfff;
rom[94088] = 12'hfff;
rom[94089] = 12'hfff;
rom[94090] = 12'hfff;
rom[94091] = 12'hfff;
rom[94092] = 12'hfff;
rom[94093] = 12'hfff;
rom[94094] = 12'hfff;
rom[94095] = 12'hfff;
rom[94096] = 12'hfff;
rom[94097] = 12'hfff;
rom[94098] = 12'hfff;
rom[94099] = 12'hfff;
rom[94100] = 12'hfff;
rom[94101] = 12'hfff;
rom[94102] = 12'hfff;
rom[94103] = 12'hfff;
rom[94104] = 12'hfff;
rom[94105] = 12'hfff;
rom[94106] = 12'hfff;
rom[94107] = 12'hfff;
rom[94108] = 12'hfff;
rom[94109] = 12'hfff;
rom[94110] = 12'hfff;
rom[94111] = 12'hfff;
rom[94112] = 12'hfff;
rom[94113] = 12'hfff;
rom[94114] = 12'hfff;
rom[94115] = 12'hfff;
rom[94116] = 12'hfff;
rom[94117] = 12'hfff;
rom[94118] = 12'hfff;
rom[94119] = 12'hfff;
rom[94120] = 12'hfff;
rom[94121] = 12'hfff;
rom[94122] = 12'hfff;
rom[94123] = 12'hfff;
rom[94124] = 12'hfff;
rom[94125] = 12'hfff;
rom[94126] = 12'hfff;
rom[94127] = 12'hfff;
rom[94128] = 12'hfff;
rom[94129] = 12'hfff;
rom[94130] = 12'hfff;
rom[94131] = 12'hfff;
rom[94132] = 12'hfff;
rom[94133] = 12'hfff;
rom[94134] = 12'hfff;
rom[94135] = 12'hfff;
rom[94136] = 12'heee;
rom[94137] = 12'heee;
rom[94138] = 12'heee;
rom[94139] = 12'hddd;
rom[94140] = 12'hddd;
rom[94141] = 12'hddd;
rom[94142] = 12'hddd;
rom[94143] = 12'hddd;
rom[94144] = 12'hccc;
rom[94145] = 12'hccc;
rom[94146] = 12'hccc;
rom[94147] = 12'hccc;
rom[94148] = 12'hddd;
rom[94149] = 12'hddd;
rom[94150] = 12'hddd;
rom[94151] = 12'hddd;
rom[94152] = 12'hddd;
rom[94153] = 12'hddd;
rom[94154] = 12'hddd;
rom[94155] = 12'hccc;
rom[94156] = 12'hccc;
rom[94157] = 12'hccc;
rom[94158] = 12'hbbb;
rom[94159] = 12'hbbb;
rom[94160] = 12'hbbb;
rom[94161] = 12'haaa;
rom[94162] = 12'haaa;
rom[94163] = 12'haaa;
rom[94164] = 12'h999;
rom[94165] = 12'h999;
rom[94166] = 12'h999;
rom[94167] = 12'h999;
rom[94168] = 12'h999;
rom[94169] = 12'h999;
rom[94170] = 12'h999;
rom[94171] = 12'h999;
rom[94172] = 12'h999;
rom[94173] = 12'h999;
rom[94174] = 12'h999;
rom[94175] = 12'h999;
rom[94176] = 12'h999;
rom[94177] = 12'h999;
rom[94178] = 12'h999;
rom[94179] = 12'h999;
rom[94180] = 12'h999;
rom[94181] = 12'h999;
rom[94182] = 12'h888;
rom[94183] = 12'h888;
rom[94184] = 12'h888;
rom[94185] = 12'h888;
rom[94186] = 12'h888;
rom[94187] = 12'h888;
rom[94188] = 12'h888;
rom[94189] = 12'h888;
rom[94190] = 12'h888;
rom[94191] = 12'h888;
rom[94192] = 12'h888;
rom[94193] = 12'h888;
rom[94194] = 12'h888;
rom[94195] = 12'h888;
rom[94196] = 12'h888;
rom[94197] = 12'h888;
rom[94198] = 12'h888;
rom[94199] = 12'h888;
rom[94200] = 12'h888;
rom[94201] = 12'h888;
rom[94202] = 12'h888;
rom[94203] = 12'h888;
rom[94204] = 12'h888;
rom[94205] = 12'h888;
rom[94206] = 12'h888;
rom[94207] = 12'h888;
rom[94208] = 12'h777;
rom[94209] = 12'h777;
rom[94210] = 12'h777;
rom[94211] = 12'h777;
rom[94212] = 12'h777;
rom[94213] = 12'h666;
rom[94214] = 12'h666;
rom[94215] = 12'h555;
rom[94216] = 12'h555;
rom[94217] = 12'h555;
rom[94218] = 12'h444;
rom[94219] = 12'h444;
rom[94220] = 12'h444;
rom[94221] = 12'h444;
rom[94222] = 12'h444;
rom[94223] = 12'h333;
rom[94224] = 12'h444;
rom[94225] = 12'h444;
rom[94226] = 12'h444;
rom[94227] = 12'h555;
rom[94228] = 12'h555;
rom[94229] = 12'h555;
rom[94230] = 12'h666;
rom[94231] = 12'h777;
rom[94232] = 12'h777;
rom[94233] = 12'h777;
rom[94234] = 12'h888;
rom[94235] = 12'h888;
rom[94236] = 12'h888;
rom[94237] = 12'h888;
rom[94238] = 12'h777;
rom[94239] = 12'h777;
rom[94240] = 12'h666;
rom[94241] = 12'h666;
rom[94242] = 12'h555;
rom[94243] = 12'h444;
rom[94244] = 12'h333;
rom[94245] = 12'h333;
rom[94246] = 12'h333;
rom[94247] = 12'h333;
rom[94248] = 12'h333;
rom[94249] = 12'h222;
rom[94250] = 12'h222;
rom[94251] = 12'h222;
rom[94252] = 12'h222;
rom[94253] = 12'h222;
rom[94254] = 12'h222;
rom[94255] = 12'h222;
rom[94256] = 12'h222;
rom[94257] = 12'h222;
rom[94258] = 12'h222;
rom[94259] = 12'h222;
rom[94260] = 12'h333;
rom[94261] = 12'h333;
rom[94262] = 12'h333;
rom[94263] = 12'h333;
rom[94264] = 12'h444;
rom[94265] = 12'h444;
rom[94266] = 12'h444;
rom[94267] = 12'h555;
rom[94268] = 12'h666;
rom[94269] = 12'h777;
rom[94270] = 12'h888;
rom[94271] = 12'h999;
rom[94272] = 12'h999;
rom[94273] = 12'h999;
rom[94274] = 12'h888;
rom[94275] = 12'h888;
rom[94276] = 12'h888;
rom[94277] = 12'h888;
rom[94278] = 12'h888;
rom[94279] = 12'h888;
rom[94280] = 12'h888;
rom[94281] = 12'h888;
rom[94282] = 12'h888;
rom[94283] = 12'h888;
rom[94284] = 12'h888;
rom[94285] = 12'h999;
rom[94286] = 12'h999;
rom[94287] = 12'h999;
rom[94288] = 12'h999;
rom[94289] = 12'h999;
rom[94290] = 12'haaa;
rom[94291] = 12'haaa;
rom[94292] = 12'hbbb;
rom[94293] = 12'hccc;
rom[94294] = 12'hddd;
rom[94295] = 12'heee;
rom[94296] = 12'heee;
rom[94297] = 12'hddd;
rom[94298] = 12'hbbb;
rom[94299] = 12'hccc;
rom[94300] = 12'hccc;
rom[94301] = 12'hccc;
rom[94302] = 12'hddd;
rom[94303] = 12'heee;
rom[94304] = 12'heee;
rom[94305] = 12'hfff;
rom[94306] = 12'hfff;
rom[94307] = 12'hfff;
rom[94308] = 12'hfff;
rom[94309] = 12'hfff;
rom[94310] = 12'heee;
rom[94311] = 12'hddd;
rom[94312] = 12'hccc;
rom[94313] = 12'hbbb;
rom[94314] = 12'h999;
rom[94315] = 12'h777;
rom[94316] = 12'h555;
rom[94317] = 12'h444;
rom[94318] = 12'h444;
rom[94319] = 12'h444;
rom[94320] = 12'h444;
rom[94321] = 12'h444;
rom[94322] = 12'h444;
rom[94323] = 12'h444;
rom[94324] = 12'h333;
rom[94325] = 12'h333;
rom[94326] = 12'h333;
rom[94327] = 12'h333;
rom[94328] = 12'h333;
rom[94329] = 12'h333;
rom[94330] = 12'h333;
rom[94331] = 12'h333;
rom[94332] = 12'h333;
rom[94333] = 12'h333;
rom[94334] = 12'h333;
rom[94335] = 12'h222;
rom[94336] = 12'h222;
rom[94337] = 12'h222;
rom[94338] = 12'h111;
rom[94339] = 12'h111;
rom[94340] = 12'h111;
rom[94341] = 12'h111;
rom[94342] = 12'h111;
rom[94343] = 12'h111;
rom[94344] = 12'h111;
rom[94345] = 12'h111;
rom[94346] = 12'h111;
rom[94347] = 12'h111;
rom[94348] = 12'h111;
rom[94349] = 12'h111;
rom[94350] = 12'h111;
rom[94351] = 12'h111;
rom[94352] = 12'h111;
rom[94353] = 12'h111;
rom[94354] = 12'h222;
rom[94355] = 12'h222;
rom[94356] = 12'h222;
rom[94357] = 12'h222;
rom[94358] = 12'h222;
rom[94359] = 12'h222;
rom[94360] = 12'h222;
rom[94361] = 12'h333;
rom[94362] = 12'h333;
rom[94363] = 12'h333;
rom[94364] = 12'h333;
rom[94365] = 12'h333;
rom[94366] = 12'h444;
rom[94367] = 12'h555;
rom[94368] = 12'h555;
rom[94369] = 12'h777;
rom[94370] = 12'h999;
rom[94371] = 12'hbbb;
rom[94372] = 12'hddd;
rom[94373] = 12'hddd;
rom[94374] = 12'hccc;
rom[94375] = 12'hbbb;
rom[94376] = 12'h999;
rom[94377] = 12'h777;
rom[94378] = 12'h555;
rom[94379] = 12'h333;
rom[94380] = 12'h333;
rom[94381] = 12'h222;
rom[94382] = 12'h222;
rom[94383] = 12'h222;
rom[94384] = 12'h222;
rom[94385] = 12'h222;
rom[94386] = 12'h222;
rom[94387] = 12'h222;
rom[94388] = 12'h222;
rom[94389] = 12'h222;
rom[94390] = 12'h111;
rom[94391] = 12'h111;
rom[94392] = 12'h111;
rom[94393] = 12'h111;
rom[94394] = 12'h111;
rom[94395] = 12'h111;
rom[94396] = 12'h111;
rom[94397] = 12'h111;
rom[94398] = 12'h111;
rom[94399] = 12'h111;
rom[94400] = 12'hfff;
rom[94401] = 12'hfff;
rom[94402] = 12'hfff;
rom[94403] = 12'hfff;
rom[94404] = 12'hfff;
rom[94405] = 12'hfff;
rom[94406] = 12'hfff;
rom[94407] = 12'hfff;
rom[94408] = 12'hfff;
rom[94409] = 12'hfff;
rom[94410] = 12'hfff;
rom[94411] = 12'hfff;
rom[94412] = 12'hfff;
rom[94413] = 12'hfff;
rom[94414] = 12'hfff;
rom[94415] = 12'hfff;
rom[94416] = 12'hfff;
rom[94417] = 12'hfff;
rom[94418] = 12'hfff;
rom[94419] = 12'hfff;
rom[94420] = 12'hfff;
rom[94421] = 12'hfff;
rom[94422] = 12'hfff;
rom[94423] = 12'hfff;
rom[94424] = 12'hfff;
rom[94425] = 12'hfff;
rom[94426] = 12'hfff;
rom[94427] = 12'hfff;
rom[94428] = 12'hfff;
rom[94429] = 12'hfff;
rom[94430] = 12'hfff;
rom[94431] = 12'hfff;
rom[94432] = 12'hfff;
rom[94433] = 12'hfff;
rom[94434] = 12'hfff;
rom[94435] = 12'hfff;
rom[94436] = 12'hfff;
rom[94437] = 12'hfff;
rom[94438] = 12'hfff;
rom[94439] = 12'hfff;
rom[94440] = 12'hfff;
rom[94441] = 12'hfff;
rom[94442] = 12'hfff;
rom[94443] = 12'hfff;
rom[94444] = 12'hfff;
rom[94445] = 12'hfff;
rom[94446] = 12'hfff;
rom[94447] = 12'hfff;
rom[94448] = 12'hfff;
rom[94449] = 12'hfff;
rom[94450] = 12'hfff;
rom[94451] = 12'hfff;
rom[94452] = 12'hfff;
rom[94453] = 12'hfff;
rom[94454] = 12'hfff;
rom[94455] = 12'hfff;
rom[94456] = 12'hfff;
rom[94457] = 12'hfff;
rom[94458] = 12'hfff;
rom[94459] = 12'hfff;
rom[94460] = 12'hfff;
rom[94461] = 12'hfff;
rom[94462] = 12'hfff;
rom[94463] = 12'hfff;
rom[94464] = 12'hfff;
rom[94465] = 12'hfff;
rom[94466] = 12'hfff;
rom[94467] = 12'hfff;
rom[94468] = 12'hfff;
rom[94469] = 12'hfff;
rom[94470] = 12'hfff;
rom[94471] = 12'hfff;
rom[94472] = 12'hfff;
rom[94473] = 12'hfff;
rom[94474] = 12'hfff;
rom[94475] = 12'hfff;
rom[94476] = 12'hfff;
rom[94477] = 12'hfff;
rom[94478] = 12'hfff;
rom[94479] = 12'hfff;
rom[94480] = 12'hfff;
rom[94481] = 12'hfff;
rom[94482] = 12'hfff;
rom[94483] = 12'hfff;
rom[94484] = 12'hfff;
rom[94485] = 12'hfff;
rom[94486] = 12'hfff;
rom[94487] = 12'hfff;
rom[94488] = 12'hfff;
rom[94489] = 12'hfff;
rom[94490] = 12'hfff;
rom[94491] = 12'hfff;
rom[94492] = 12'hfff;
rom[94493] = 12'hfff;
rom[94494] = 12'hfff;
rom[94495] = 12'hfff;
rom[94496] = 12'hfff;
rom[94497] = 12'hfff;
rom[94498] = 12'hfff;
rom[94499] = 12'hfff;
rom[94500] = 12'hfff;
rom[94501] = 12'hfff;
rom[94502] = 12'hfff;
rom[94503] = 12'hfff;
rom[94504] = 12'hfff;
rom[94505] = 12'hfff;
rom[94506] = 12'hfff;
rom[94507] = 12'hfff;
rom[94508] = 12'hfff;
rom[94509] = 12'hfff;
rom[94510] = 12'hfff;
rom[94511] = 12'hfff;
rom[94512] = 12'hfff;
rom[94513] = 12'hfff;
rom[94514] = 12'hfff;
rom[94515] = 12'hfff;
rom[94516] = 12'hfff;
rom[94517] = 12'hfff;
rom[94518] = 12'hfff;
rom[94519] = 12'hfff;
rom[94520] = 12'hfff;
rom[94521] = 12'hfff;
rom[94522] = 12'hfff;
rom[94523] = 12'hfff;
rom[94524] = 12'hfff;
rom[94525] = 12'hfff;
rom[94526] = 12'hfff;
rom[94527] = 12'hfff;
rom[94528] = 12'hfff;
rom[94529] = 12'hfff;
rom[94530] = 12'hfff;
rom[94531] = 12'hfff;
rom[94532] = 12'hfff;
rom[94533] = 12'hfff;
rom[94534] = 12'hfff;
rom[94535] = 12'hfff;
rom[94536] = 12'hfff;
rom[94537] = 12'heee;
rom[94538] = 12'heee;
rom[94539] = 12'heee;
rom[94540] = 12'heee;
rom[94541] = 12'hddd;
rom[94542] = 12'hddd;
rom[94543] = 12'hddd;
rom[94544] = 12'hddd;
rom[94545] = 12'hccc;
rom[94546] = 12'hccc;
rom[94547] = 12'hccc;
rom[94548] = 12'hccc;
rom[94549] = 12'hddd;
rom[94550] = 12'hddd;
rom[94551] = 12'hddd;
rom[94552] = 12'hddd;
rom[94553] = 12'hddd;
rom[94554] = 12'hddd;
rom[94555] = 12'hddd;
rom[94556] = 12'hccc;
rom[94557] = 12'hccc;
rom[94558] = 12'hccc;
rom[94559] = 12'hccc;
rom[94560] = 12'hccc;
rom[94561] = 12'hbbb;
rom[94562] = 12'hbbb;
rom[94563] = 12'hbbb;
rom[94564] = 12'haaa;
rom[94565] = 12'haaa;
rom[94566] = 12'haaa;
rom[94567] = 12'haaa;
rom[94568] = 12'haaa;
rom[94569] = 12'haaa;
rom[94570] = 12'haaa;
rom[94571] = 12'haaa;
rom[94572] = 12'haaa;
rom[94573] = 12'haaa;
rom[94574] = 12'haaa;
rom[94575] = 12'haaa;
rom[94576] = 12'h999;
rom[94577] = 12'h999;
rom[94578] = 12'h999;
rom[94579] = 12'h999;
rom[94580] = 12'h999;
rom[94581] = 12'h999;
rom[94582] = 12'h888;
rom[94583] = 12'h888;
rom[94584] = 12'h888;
rom[94585] = 12'h888;
rom[94586] = 12'h888;
rom[94587] = 12'h888;
rom[94588] = 12'h888;
rom[94589] = 12'h888;
rom[94590] = 12'h888;
rom[94591] = 12'h888;
rom[94592] = 12'h888;
rom[94593] = 12'h888;
rom[94594] = 12'h888;
rom[94595] = 12'h888;
rom[94596] = 12'h888;
rom[94597] = 12'h888;
rom[94598] = 12'h888;
rom[94599] = 12'h888;
rom[94600] = 12'h888;
rom[94601] = 12'h888;
rom[94602] = 12'h888;
rom[94603] = 12'h888;
rom[94604] = 12'h888;
rom[94605] = 12'h888;
rom[94606] = 12'h888;
rom[94607] = 12'h888;
rom[94608] = 12'h888;
rom[94609] = 12'h888;
rom[94610] = 12'h888;
rom[94611] = 12'h777;
rom[94612] = 12'h777;
rom[94613] = 12'h777;
rom[94614] = 12'h666;
rom[94615] = 12'h666;
rom[94616] = 12'h555;
rom[94617] = 12'h555;
rom[94618] = 12'h555;
rom[94619] = 12'h555;
rom[94620] = 12'h555;
rom[94621] = 12'h555;
rom[94622] = 12'h555;
rom[94623] = 12'h444;
rom[94624] = 12'h555;
rom[94625] = 12'h555;
rom[94626] = 12'h555;
rom[94627] = 12'h555;
rom[94628] = 12'h555;
rom[94629] = 12'h666;
rom[94630] = 12'h666;
rom[94631] = 12'h777;
rom[94632] = 12'h777;
rom[94633] = 12'h888;
rom[94634] = 12'h888;
rom[94635] = 12'h888;
rom[94636] = 12'h888;
rom[94637] = 12'h888;
rom[94638] = 12'h888;
rom[94639] = 12'h777;
rom[94640] = 12'h777;
rom[94641] = 12'h666;
rom[94642] = 12'h666;
rom[94643] = 12'h555;
rom[94644] = 12'h555;
rom[94645] = 12'h444;
rom[94646] = 12'h444;
rom[94647] = 12'h333;
rom[94648] = 12'h333;
rom[94649] = 12'h333;
rom[94650] = 12'h333;
rom[94651] = 12'h333;
rom[94652] = 12'h333;
rom[94653] = 12'h333;
rom[94654] = 12'h333;
rom[94655] = 12'h222;
rom[94656] = 12'h333;
rom[94657] = 12'h333;
rom[94658] = 12'h333;
rom[94659] = 12'h333;
rom[94660] = 12'h444;
rom[94661] = 12'h444;
rom[94662] = 12'h444;
rom[94663] = 12'h444;
rom[94664] = 12'h555;
rom[94665] = 12'h555;
rom[94666] = 12'h666;
rom[94667] = 12'h777;
rom[94668] = 12'h777;
rom[94669] = 12'h888;
rom[94670] = 12'h888;
rom[94671] = 12'h999;
rom[94672] = 12'h999;
rom[94673] = 12'h888;
rom[94674] = 12'h888;
rom[94675] = 12'h888;
rom[94676] = 12'h888;
rom[94677] = 12'h888;
rom[94678] = 12'h888;
rom[94679] = 12'h888;
rom[94680] = 12'h888;
rom[94681] = 12'h888;
rom[94682] = 12'h888;
rom[94683] = 12'h888;
rom[94684] = 12'h888;
rom[94685] = 12'h888;
rom[94686] = 12'h999;
rom[94687] = 12'h999;
rom[94688] = 12'h999;
rom[94689] = 12'h999;
rom[94690] = 12'haaa;
rom[94691] = 12'haaa;
rom[94692] = 12'hccc;
rom[94693] = 12'hddd;
rom[94694] = 12'heee;
rom[94695] = 12'hfff;
rom[94696] = 12'heee;
rom[94697] = 12'hccc;
rom[94698] = 12'hbbb;
rom[94699] = 12'hbbb;
rom[94700] = 12'hbbb;
rom[94701] = 12'haaa;
rom[94702] = 12'hbbb;
rom[94703] = 12'hccc;
rom[94704] = 12'hddd;
rom[94705] = 12'heee;
rom[94706] = 12'hfff;
rom[94707] = 12'hfff;
rom[94708] = 12'hfff;
rom[94709] = 12'hfff;
rom[94710] = 12'hfff;
rom[94711] = 12'hfff;
rom[94712] = 12'heee;
rom[94713] = 12'hddd;
rom[94714] = 12'hccc;
rom[94715] = 12'haaa;
rom[94716] = 12'h777;
rom[94717] = 12'h555;
rom[94718] = 12'h444;
rom[94719] = 12'h444;
rom[94720] = 12'h444;
rom[94721] = 12'h444;
rom[94722] = 12'h444;
rom[94723] = 12'h444;
rom[94724] = 12'h444;
rom[94725] = 12'h333;
rom[94726] = 12'h333;
rom[94727] = 12'h333;
rom[94728] = 12'h333;
rom[94729] = 12'h333;
rom[94730] = 12'h222;
rom[94731] = 12'h222;
rom[94732] = 12'h333;
rom[94733] = 12'h333;
rom[94734] = 12'h333;
rom[94735] = 12'h333;
rom[94736] = 12'h222;
rom[94737] = 12'h222;
rom[94738] = 12'h222;
rom[94739] = 12'h111;
rom[94740] = 12'h111;
rom[94741] = 12'h111;
rom[94742] = 12'h111;
rom[94743] = 12'h111;
rom[94744] = 12'h  0;
rom[94745] = 12'h111;
rom[94746] = 12'h111;
rom[94747] = 12'h111;
rom[94748] = 12'h111;
rom[94749] = 12'h111;
rom[94750] = 12'h111;
rom[94751] = 12'h  0;
rom[94752] = 12'h111;
rom[94753] = 12'h111;
rom[94754] = 12'h111;
rom[94755] = 12'h222;
rom[94756] = 12'h222;
rom[94757] = 12'h222;
rom[94758] = 12'h222;
rom[94759] = 12'h222;
rom[94760] = 12'h222;
rom[94761] = 12'h222;
rom[94762] = 12'h222;
rom[94763] = 12'h222;
rom[94764] = 12'h333;
rom[94765] = 12'h333;
rom[94766] = 12'h333;
rom[94767] = 12'h444;
rom[94768] = 12'h444;
rom[94769] = 12'h555;
rom[94770] = 12'h666;
rom[94771] = 12'h888;
rom[94772] = 12'haaa;
rom[94773] = 12'hbbb;
rom[94774] = 12'hccc;
rom[94775] = 12'hccc;
rom[94776] = 12'hbbb;
rom[94777] = 12'haaa;
rom[94778] = 12'h888;
rom[94779] = 12'h666;
rom[94780] = 12'h555;
rom[94781] = 12'h444;
rom[94782] = 12'h333;
rom[94783] = 12'h222;
rom[94784] = 12'h222;
rom[94785] = 12'h222;
rom[94786] = 12'h222;
rom[94787] = 12'h222;
rom[94788] = 12'h222;
rom[94789] = 12'h222;
rom[94790] = 12'h222;
rom[94791] = 12'h111;
rom[94792] = 12'h111;
rom[94793] = 12'h111;
rom[94794] = 12'h111;
rom[94795] = 12'h111;
rom[94796] = 12'h111;
rom[94797] = 12'h111;
rom[94798] = 12'h111;
rom[94799] = 12'h111;
rom[94800] = 12'hfff;
rom[94801] = 12'hfff;
rom[94802] = 12'hfff;
rom[94803] = 12'hfff;
rom[94804] = 12'hfff;
rom[94805] = 12'hfff;
rom[94806] = 12'hfff;
rom[94807] = 12'hfff;
rom[94808] = 12'hfff;
rom[94809] = 12'hfff;
rom[94810] = 12'hfff;
rom[94811] = 12'hfff;
rom[94812] = 12'hfff;
rom[94813] = 12'hfff;
rom[94814] = 12'hfff;
rom[94815] = 12'hfff;
rom[94816] = 12'hfff;
rom[94817] = 12'hfff;
rom[94818] = 12'hfff;
rom[94819] = 12'hfff;
rom[94820] = 12'hfff;
rom[94821] = 12'hfff;
rom[94822] = 12'hfff;
rom[94823] = 12'hfff;
rom[94824] = 12'hfff;
rom[94825] = 12'hfff;
rom[94826] = 12'hfff;
rom[94827] = 12'hfff;
rom[94828] = 12'hfff;
rom[94829] = 12'hfff;
rom[94830] = 12'hfff;
rom[94831] = 12'hfff;
rom[94832] = 12'hfff;
rom[94833] = 12'hfff;
rom[94834] = 12'hfff;
rom[94835] = 12'hfff;
rom[94836] = 12'hfff;
rom[94837] = 12'hfff;
rom[94838] = 12'hfff;
rom[94839] = 12'hfff;
rom[94840] = 12'hfff;
rom[94841] = 12'hfff;
rom[94842] = 12'hfff;
rom[94843] = 12'hfff;
rom[94844] = 12'hfff;
rom[94845] = 12'hfff;
rom[94846] = 12'hfff;
rom[94847] = 12'hfff;
rom[94848] = 12'hfff;
rom[94849] = 12'hfff;
rom[94850] = 12'hfff;
rom[94851] = 12'hfff;
rom[94852] = 12'hfff;
rom[94853] = 12'hfff;
rom[94854] = 12'hfff;
rom[94855] = 12'hfff;
rom[94856] = 12'hfff;
rom[94857] = 12'hfff;
rom[94858] = 12'hfff;
rom[94859] = 12'hfff;
rom[94860] = 12'hfff;
rom[94861] = 12'hfff;
rom[94862] = 12'hfff;
rom[94863] = 12'hfff;
rom[94864] = 12'hfff;
rom[94865] = 12'hfff;
rom[94866] = 12'hfff;
rom[94867] = 12'hfff;
rom[94868] = 12'hfff;
rom[94869] = 12'hfff;
rom[94870] = 12'hfff;
rom[94871] = 12'hfff;
rom[94872] = 12'hfff;
rom[94873] = 12'hfff;
rom[94874] = 12'hfff;
rom[94875] = 12'hfff;
rom[94876] = 12'hfff;
rom[94877] = 12'hfff;
rom[94878] = 12'hfff;
rom[94879] = 12'hfff;
rom[94880] = 12'hfff;
rom[94881] = 12'hfff;
rom[94882] = 12'hfff;
rom[94883] = 12'hfff;
rom[94884] = 12'hfff;
rom[94885] = 12'hfff;
rom[94886] = 12'hfff;
rom[94887] = 12'hfff;
rom[94888] = 12'hfff;
rom[94889] = 12'hfff;
rom[94890] = 12'hfff;
rom[94891] = 12'hfff;
rom[94892] = 12'hfff;
rom[94893] = 12'hfff;
rom[94894] = 12'hfff;
rom[94895] = 12'hfff;
rom[94896] = 12'hfff;
rom[94897] = 12'hfff;
rom[94898] = 12'hfff;
rom[94899] = 12'hfff;
rom[94900] = 12'hfff;
rom[94901] = 12'hfff;
rom[94902] = 12'hfff;
rom[94903] = 12'hfff;
rom[94904] = 12'hfff;
rom[94905] = 12'hfff;
rom[94906] = 12'hfff;
rom[94907] = 12'hfff;
rom[94908] = 12'hfff;
rom[94909] = 12'hfff;
rom[94910] = 12'hfff;
rom[94911] = 12'hfff;
rom[94912] = 12'hfff;
rom[94913] = 12'hfff;
rom[94914] = 12'hfff;
rom[94915] = 12'hfff;
rom[94916] = 12'hfff;
rom[94917] = 12'hfff;
rom[94918] = 12'hfff;
rom[94919] = 12'hfff;
rom[94920] = 12'hfff;
rom[94921] = 12'hfff;
rom[94922] = 12'hfff;
rom[94923] = 12'hfff;
rom[94924] = 12'hfff;
rom[94925] = 12'hfff;
rom[94926] = 12'hfff;
rom[94927] = 12'hfff;
rom[94928] = 12'hfff;
rom[94929] = 12'hfff;
rom[94930] = 12'hfff;
rom[94931] = 12'hfff;
rom[94932] = 12'hfff;
rom[94933] = 12'hfff;
rom[94934] = 12'hfff;
rom[94935] = 12'hfff;
rom[94936] = 12'hfff;
rom[94937] = 12'hfff;
rom[94938] = 12'heee;
rom[94939] = 12'heee;
rom[94940] = 12'heee;
rom[94941] = 12'heee;
rom[94942] = 12'hddd;
rom[94943] = 12'hddd;
rom[94944] = 12'hddd;
rom[94945] = 12'hddd;
rom[94946] = 12'hccc;
rom[94947] = 12'hccc;
rom[94948] = 12'hccc;
rom[94949] = 12'hccc;
rom[94950] = 12'hccc;
rom[94951] = 12'hccc;
rom[94952] = 12'hccc;
rom[94953] = 12'hddd;
rom[94954] = 12'hddd;
rom[94955] = 12'hddd;
rom[94956] = 12'hccc;
rom[94957] = 12'hccc;
rom[94958] = 12'hccc;
rom[94959] = 12'hccc;
rom[94960] = 12'hccc;
rom[94961] = 12'hccc;
rom[94962] = 12'hccc;
rom[94963] = 12'hbbb;
rom[94964] = 12'hbbb;
rom[94965] = 12'hbbb;
rom[94966] = 12'hbbb;
rom[94967] = 12'hbbb;
rom[94968] = 12'hbbb;
rom[94969] = 12'hbbb;
rom[94970] = 12'haaa;
rom[94971] = 12'haaa;
rom[94972] = 12'haaa;
rom[94973] = 12'haaa;
rom[94974] = 12'haaa;
rom[94975] = 12'haaa;
rom[94976] = 12'haaa;
rom[94977] = 12'h999;
rom[94978] = 12'h999;
rom[94979] = 12'h999;
rom[94980] = 12'h999;
rom[94981] = 12'h999;
rom[94982] = 12'h999;
rom[94983] = 12'h999;
rom[94984] = 12'h888;
rom[94985] = 12'h888;
rom[94986] = 12'h888;
rom[94987] = 12'h888;
rom[94988] = 12'h888;
rom[94989] = 12'h888;
rom[94990] = 12'h888;
rom[94991] = 12'h888;
rom[94992] = 12'h888;
rom[94993] = 12'h888;
rom[94994] = 12'h888;
rom[94995] = 12'h888;
rom[94996] = 12'h888;
rom[94997] = 12'h888;
rom[94998] = 12'h888;
rom[94999] = 12'h999;
rom[95000] = 12'h888;
rom[95001] = 12'h888;
rom[95002] = 12'h999;
rom[95003] = 12'h999;
rom[95004] = 12'h999;
rom[95005] = 12'h888;
rom[95006] = 12'h888;
rom[95007] = 12'h888;
rom[95008] = 12'h888;
rom[95009] = 12'h888;
rom[95010] = 12'h888;
rom[95011] = 12'h888;
rom[95012] = 12'h888;
rom[95013] = 12'h777;
rom[95014] = 12'h777;
rom[95015] = 12'h666;
rom[95016] = 12'h666;
rom[95017] = 12'h666;
rom[95018] = 12'h555;
rom[95019] = 12'h666;
rom[95020] = 12'h666;
rom[95021] = 12'h666;
rom[95022] = 12'h555;
rom[95023] = 12'h555;
rom[95024] = 12'h666;
rom[95025] = 12'h666;
rom[95026] = 12'h666;
rom[95027] = 12'h666;
rom[95028] = 12'h666;
rom[95029] = 12'h666;
rom[95030] = 12'h777;
rom[95031] = 12'h777;
rom[95032] = 12'h777;
rom[95033] = 12'h888;
rom[95034] = 12'h888;
rom[95035] = 12'h777;
rom[95036] = 12'h888;
rom[95037] = 12'h888;
rom[95038] = 12'h888;
rom[95039] = 12'h888;
rom[95040] = 12'h777;
rom[95041] = 12'h777;
rom[95042] = 12'h666;
rom[95043] = 12'h666;
rom[95044] = 12'h555;
rom[95045] = 12'h555;
rom[95046] = 12'h444;
rom[95047] = 12'h444;
rom[95048] = 12'h444;
rom[95049] = 12'h333;
rom[95050] = 12'h333;
rom[95051] = 12'h333;
rom[95052] = 12'h333;
rom[95053] = 12'h333;
rom[95054] = 12'h333;
rom[95055] = 12'h333;
rom[95056] = 12'h333;
rom[95057] = 12'h444;
rom[95058] = 12'h444;
rom[95059] = 12'h444;
rom[95060] = 12'h444;
rom[95061] = 12'h555;
rom[95062] = 12'h555;
rom[95063] = 12'h666;
rom[95064] = 12'h666;
rom[95065] = 12'h777;
rom[95066] = 12'h888;
rom[95067] = 12'h888;
rom[95068] = 12'h888;
rom[95069] = 12'h888;
rom[95070] = 12'h888;
rom[95071] = 12'h888;
rom[95072] = 12'h888;
rom[95073] = 12'h888;
rom[95074] = 12'h888;
rom[95075] = 12'h888;
rom[95076] = 12'h888;
rom[95077] = 12'h888;
rom[95078] = 12'h777;
rom[95079] = 12'h777;
rom[95080] = 12'h777;
rom[95081] = 12'h777;
rom[95082] = 12'h888;
rom[95083] = 12'h888;
rom[95084] = 12'h888;
rom[95085] = 12'h888;
rom[95086] = 12'h999;
rom[95087] = 12'h999;
rom[95088] = 12'h999;
rom[95089] = 12'h999;
rom[95090] = 12'haaa;
rom[95091] = 12'hbbb;
rom[95092] = 12'hddd;
rom[95093] = 12'heee;
rom[95094] = 12'hfff;
rom[95095] = 12'heee;
rom[95096] = 12'hddd;
rom[95097] = 12'hccc;
rom[95098] = 12'haaa;
rom[95099] = 12'haaa;
rom[95100] = 12'h999;
rom[95101] = 12'h888;
rom[95102] = 12'h888;
rom[95103] = 12'h999;
rom[95104] = 12'haaa;
rom[95105] = 12'hbbb;
rom[95106] = 12'hddd;
rom[95107] = 12'heee;
rom[95108] = 12'hfff;
rom[95109] = 12'hfff;
rom[95110] = 12'hfff;
rom[95111] = 12'hfff;
rom[95112] = 12'hfff;
rom[95113] = 12'hfff;
rom[95114] = 12'hfff;
rom[95115] = 12'hddd;
rom[95116] = 12'hbbb;
rom[95117] = 12'h888;
rom[95118] = 12'h666;
rom[95119] = 12'h555;
rom[95120] = 12'h444;
rom[95121] = 12'h444;
rom[95122] = 12'h444;
rom[95123] = 12'h444;
rom[95124] = 12'h444;
rom[95125] = 12'h333;
rom[95126] = 12'h333;
rom[95127] = 12'h333;
rom[95128] = 12'h333;
rom[95129] = 12'h333;
rom[95130] = 12'h222;
rom[95131] = 12'h222;
rom[95132] = 12'h222;
rom[95133] = 12'h222;
rom[95134] = 12'h333;
rom[95135] = 12'h333;
rom[95136] = 12'h333;
rom[95137] = 12'h333;
rom[95138] = 12'h222;
rom[95139] = 12'h111;
rom[95140] = 12'h111;
rom[95141] = 12'h111;
rom[95142] = 12'h  0;
rom[95143] = 12'h  0;
rom[95144] = 12'h  0;
rom[95145] = 12'h  0;
rom[95146] = 12'h111;
rom[95147] = 12'h111;
rom[95148] = 12'h111;
rom[95149] = 12'h111;
rom[95150] = 12'h  0;
rom[95151] = 12'h  0;
rom[95152] = 12'h111;
rom[95153] = 12'h111;
rom[95154] = 12'h111;
rom[95155] = 12'h111;
rom[95156] = 12'h111;
rom[95157] = 12'h222;
rom[95158] = 12'h222;
rom[95159] = 12'h222;
rom[95160] = 12'h222;
rom[95161] = 12'h222;
rom[95162] = 12'h111;
rom[95163] = 12'h222;
rom[95164] = 12'h222;
rom[95165] = 12'h333;
rom[95166] = 12'h333;
rom[95167] = 12'h222;
rom[95168] = 12'h333;
rom[95169] = 12'h444;
rom[95170] = 12'h555;
rom[95171] = 12'h666;
rom[95172] = 12'h777;
rom[95173] = 12'h888;
rom[95174] = 12'haaa;
rom[95175] = 12'hbbb;
rom[95176] = 12'hbbb;
rom[95177] = 12'hbbb;
rom[95178] = 12'hbbb;
rom[95179] = 12'haaa;
rom[95180] = 12'h888;
rom[95181] = 12'h666;
rom[95182] = 12'h444;
rom[95183] = 12'h333;
rom[95184] = 12'h222;
rom[95185] = 12'h222;
rom[95186] = 12'h111;
rom[95187] = 12'h111;
rom[95188] = 12'h111;
rom[95189] = 12'h111;
rom[95190] = 12'h111;
rom[95191] = 12'h111;
rom[95192] = 12'h111;
rom[95193] = 12'h111;
rom[95194] = 12'h111;
rom[95195] = 12'h111;
rom[95196] = 12'h111;
rom[95197] = 12'h111;
rom[95198] = 12'h111;
rom[95199] = 12'h111;
rom[95200] = 12'hfff;
rom[95201] = 12'hfff;
rom[95202] = 12'hfff;
rom[95203] = 12'hfff;
rom[95204] = 12'hfff;
rom[95205] = 12'hfff;
rom[95206] = 12'hfff;
rom[95207] = 12'hfff;
rom[95208] = 12'hfff;
rom[95209] = 12'hfff;
rom[95210] = 12'hfff;
rom[95211] = 12'hfff;
rom[95212] = 12'hfff;
rom[95213] = 12'hfff;
rom[95214] = 12'hfff;
rom[95215] = 12'hfff;
rom[95216] = 12'hfff;
rom[95217] = 12'hfff;
rom[95218] = 12'hfff;
rom[95219] = 12'hfff;
rom[95220] = 12'hfff;
rom[95221] = 12'hfff;
rom[95222] = 12'hfff;
rom[95223] = 12'hfff;
rom[95224] = 12'hfff;
rom[95225] = 12'hfff;
rom[95226] = 12'hfff;
rom[95227] = 12'hfff;
rom[95228] = 12'hfff;
rom[95229] = 12'hfff;
rom[95230] = 12'hfff;
rom[95231] = 12'hfff;
rom[95232] = 12'hfff;
rom[95233] = 12'hfff;
rom[95234] = 12'hfff;
rom[95235] = 12'hfff;
rom[95236] = 12'hfff;
rom[95237] = 12'hfff;
rom[95238] = 12'hfff;
rom[95239] = 12'hfff;
rom[95240] = 12'hfff;
rom[95241] = 12'hfff;
rom[95242] = 12'hfff;
rom[95243] = 12'hfff;
rom[95244] = 12'hfff;
rom[95245] = 12'hfff;
rom[95246] = 12'hfff;
rom[95247] = 12'hfff;
rom[95248] = 12'hfff;
rom[95249] = 12'hfff;
rom[95250] = 12'hfff;
rom[95251] = 12'hfff;
rom[95252] = 12'hfff;
rom[95253] = 12'hfff;
rom[95254] = 12'hfff;
rom[95255] = 12'hfff;
rom[95256] = 12'hfff;
rom[95257] = 12'hfff;
rom[95258] = 12'hfff;
rom[95259] = 12'hfff;
rom[95260] = 12'hfff;
rom[95261] = 12'hfff;
rom[95262] = 12'hfff;
rom[95263] = 12'hfff;
rom[95264] = 12'hfff;
rom[95265] = 12'hfff;
rom[95266] = 12'hfff;
rom[95267] = 12'hfff;
rom[95268] = 12'hfff;
rom[95269] = 12'hfff;
rom[95270] = 12'hfff;
rom[95271] = 12'hfff;
rom[95272] = 12'hfff;
rom[95273] = 12'hfff;
rom[95274] = 12'hfff;
rom[95275] = 12'hfff;
rom[95276] = 12'hfff;
rom[95277] = 12'hfff;
rom[95278] = 12'hfff;
rom[95279] = 12'hfff;
rom[95280] = 12'hfff;
rom[95281] = 12'hfff;
rom[95282] = 12'hfff;
rom[95283] = 12'hfff;
rom[95284] = 12'hfff;
rom[95285] = 12'hfff;
rom[95286] = 12'hfff;
rom[95287] = 12'hfff;
rom[95288] = 12'hfff;
rom[95289] = 12'hfff;
rom[95290] = 12'hfff;
rom[95291] = 12'hfff;
rom[95292] = 12'hfff;
rom[95293] = 12'hfff;
rom[95294] = 12'hfff;
rom[95295] = 12'hfff;
rom[95296] = 12'hfff;
rom[95297] = 12'hfff;
rom[95298] = 12'hfff;
rom[95299] = 12'hfff;
rom[95300] = 12'hfff;
rom[95301] = 12'hfff;
rom[95302] = 12'hfff;
rom[95303] = 12'hfff;
rom[95304] = 12'hfff;
rom[95305] = 12'hfff;
rom[95306] = 12'hfff;
rom[95307] = 12'hfff;
rom[95308] = 12'hfff;
rom[95309] = 12'hfff;
rom[95310] = 12'hfff;
rom[95311] = 12'hfff;
rom[95312] = 12'hfff;
rom[95313] = 12'hfff;
rom[95314] = 12'hfff;
rom[95315] = 12'hfff;
rom[95316] = 12'hfff;
rom[95317] = 12'hfff;
rom[95318] = 12'hfff;
rom[95319] = 12'hfff;
rom[95320] = 12'hfff;
rom[95321] = 12'hfff;
rom[95322] = 12'hfff;
rom[95323] = 12'hfff;
rom[95324] = 12'hfff;
rom[95325] = 12'hfff;
rom[95326] = 12'hfff;
rom[95327] = 12'hfff;
rom[95328] = 12'hfff;
rom[95329] = 12'hfff;
rom[95330] = 12'hfff;
rom[95331] = 12'hfff;
rom[95332] = 12'hfff;
rom[95333] = 12'hfff;
rom[95334] = 12'hfff;
rom[95335] = 12'hfff;
rom[95336] = 12'hfff;
rom[95337] = 12'hfff;
rom[95338] = 12'hfff;
rom[95339] = 12'heee;
rom[95340] = 12'heee;
rom[95341] = 12'heee;
rom[95342] = 12'heee;
rom[95343] = 12'hddd;
rom[95344] = 12'hddd;
rom[95345] = 12'hddd;
rom[95346] = 12'hddd;
rom[95347] = 12'hccc;
rom[95348] = 12'hccc;
rom[95349] = 12'hccc;
rom[95350] = 12'hccc;
rom[95351] = 12'hccc;
rom[95352] = 12'hccc;
rom[95353] = 12'hccc;
rom[95354] = 12'hccc;
rom[95355] = 12'hccc;
rom[95356] = 12'hccc;
rom[95357] = 12'hccc;
rom[95358] = 12'hccc;
rom[95359] = 12'hccc;
rom[95360] = 12'hccc;
rom[95361] = 12'hccc;
rom[95362] = 12'hccc;
rom[95363] = 12'hccc;
rom[95364] = 12'hbbb;
rom[95365] = 12'hbbb;
rom[95366] = 12'hbbb;
rom[95367] = 12'hbbb;
rom[95368] = 12'hbbb;
rom[95369] = 12'hbbb;
rom[95370] = 12'hbbb;
rom[95371] = 12'haaa;
rom[95372] = 12'haaa;
rom[95373] = 12'haaa;
rom[95374] = 12'haaa;
rom[95375] = 12'haaa;
rom[95376] = 12'haaa;
rom[95377] = 12'h999;
rom[95378] = 12'h999;
rom[95379] = 12'h999;
rom[95380] = 12'h999;
rom[95381] = 12'h999;
rom[95382] = 12'h999;
rom[95383] = 12'h999;
rom[95384] = 12'h999;
rom[95385] = 12'h999;
rom[95386] = 12'h888;
rom[95387] = 12'h888;
rom[95388] = 12'h888;
rom[95389] = 12'h888;
rom[95390] = 12'h888;
rom[95391] = 12'h888;
rom[95392] = 12'h888;
rom[95393] = 12'h888;
rom[95394] = 12'h888;
rom[95395] = 12'h888;
rom[95396] = 12'h888;
rom[95397] = 12'h888;
rom[95398] = 12'h999;
rom[95399] = 12'h999;
rom[95400] = 12'h999;
rom[95401] = 12'h999;
rom[95402] = 12'h999;
rom[95403] = 12'h999;
rom[95404] = 12'h999;
rom[95405] = 12'h999;
rom[95406] = 12'h999;
rom[95407] = 12'h999;
rom[95408] = 12'h888;
rom[95409] = 12'h888;
rom[95410] = 12'h888;
rom[95411] = 12'h888;
rom[95412] = 12'h888;
rom[95413] = 12'h888;
rom[95414] = 12'h777;
rom[95415] = 12'h777;
rom[95416] = 12'h777;
rom[95417] = 12'h666;
rom[95418] = 12'h666;
rom[95419] = 12'h666;
rom[95420] = 12'h666;
rom[95421] = 12'h666;
rom[95422] = 12'h666;
rom[95423] = 12'h666;
rom[95424] = 12'h666;
rom[95425] = 12'h666;
rom[95426] = 12'h666;
rom[95427] = 12'h666;
rom[95428] = 12'h666;
rom[95429] = 12'h666;
rom[95430] = 12'h777;
rom[95431] = 12'h777;
rom[95432] = 12'h777;
rom[95433] = 12'h888;
rom[95434] = 12'h888;
rom[95435] = 12'h888;
rom[95436] = 12'h888;
rom[95437] = 12'h999;
rom[95438] = 12'h999;
rom[95439] = 12'h888;
rom[95440] = 12'h888;
rom[95441] = 12'h777;
rom[95442] = 12'h777;
rom[95443] = 12'h666;
rom[95444] = 12'h666;
rom[95445] = 12'h666;
rom[95446] = 12'h555;
rom[95447] = 12'h555;
rom[95448] = 12'h444;
rom[95449] = 12'h444;
rom[95450] = 12'h444;
rom[95451] = 12'h444;
rom[95452] = 12'h444;
rom[95453] = 12'h444;
rom[95454] = 12'h444;
rom[95455] = 12'h444;
rom[95456] = 12'h444;
rom[95457] = 12'h555;
rom[95458] = 12'h555;
rom[95459] = 12'h555;
rom[95460] = 12'h555;
rom[95461] = 12'h666;
rom[95462] = 12'h666;
rom[95463] = 12'h777;
rom[95464] = 12'h777;
rom[95465] = 12'h888;
rom[95466] = 12'h888;
rom[95467] = 12'h999;
rom[95468] = 12'h999;
rom[95469] = 12'h888;
rom[95470] = 12'h888;
rom[95471] = 12'h888;
rom[95472] = 12'h888;
rom[95473] = 12'h888;
rom[95474] = 12'h888;
rom[95475] = 12'h888;
rom[95476] = 12'h777;
rom[95477] = 12'h777;
rom[95478] = 12'h777;
rom[95479] = 12'h777;
rom[95480] = 12'h777;
rom[95481] = 12'h777;
rom[95482] = 12'h888;
rom[95483] = 12'h888;
rom[95484] = 12'h888;
rom[95485] = 12'h888;
rom[95486] = 12'h888;
rom[95487] = 12'h999;
rom[95488] = 12'h999;
rom[95489] = 12'haaa;
rom[95490] = 12'hbbb;
rom[95491] = 12'hccc;
rom[95492] = 12'heee;
rom[95493] = 12'hfff;
rom[95494] = 12'heee;
rom[95495] = 12'heee;
rom[95496] = 12'hccc;
rom[95497] = 12'hbbb;
rom[95498] = 12'haaa;
rom[95499] = 12'h999;
rom[95500] = 12'h888;
rom[95501] = 12'h777;
rom[95502] = 12'h777;
rom[95503] = 12'h777;
rom[95504] = 12'h777;
rom[95505] = 12'h888;
rom[95506] = 12'h999;
rom[95507] = 12'haaa;
rom[95508] = 12'hccc;
rom[95509] = 12'hddd;
rom[95510] = 12'heee;
rom[95511] = 12'hfff;
rom[95512] = 12'hfff;
rom[95513] = 12'hfff;
rom[95514] = 12'hfff;
rom[95515] = 12'hfff;
rom[95516] = 12'heee;
rom[95517] = 12'hccc;
rom[95518] = 12'haaa;
rom[95519] = 12'h888;
rom[95520] = 12'h666;
rom[95521] = 12'h555;
rom[95522] = 12'h444;
rom[95523] = 12'h333;
rom[95524] = 12'h333;
rom[95525] = 12'h333;
rom[95526] = 12'h333;
rom[95527] = 12'h333;
rom[95528] = 12'h333;
rom[95529] = 12'h333;
rom[95530] = 12'h222;
rom[95531] = 12'h222;
rom[95532] = 12'h222;
rom[95533] = 12'h222;
rom[95534] = 12'h222;
rom[95535] = 12'h222;
rom[95536] = 12'h333;
rom[95537] = 12'h333;
rom[95538] = 12'h222;
rom[95539] = 12'h222;
rom[95540] = 12'h111;
rom[95541] = 12'h111;
rom[95542] = 12'h111;
rom[95543] = 12'h  0;
rom[95544] = 12'h  0;
rom[95545] = 12'h  0;
rom[95546] = 12'h  0;
rom[95547] = 12'h111;
rom[95548] = 12'h111;
rom[95549] = 12'h111;
rom[95550] = 12'h  0;
rom[95551] = 12'h  0;
rom[95552] = 12'h111;
rom[95553] = 12'h111;
rom[95554] = 12'h111;
rom[95555] = 12'h111;
rom[95556] = 12'h111;
rom[95557] = 12'h111;
rom[95558] = 12'h222;
rom[95559] = 12'h222;
rom[95560] = 12'h222;
rom[95561] = 12'h222;
rom[95562] = 12'h222;
rom[95563] = 12'h222;
rom[95564] = 12'h222;
rom[95565] = 12'h222;
rom[95566] = 12'h222;
rom[95567] = 12'h222;
rom[95568] = 12'h222;
rom[95569] = 12'h333;
rom[95570] = 12'h333;
rom[95571] = 12'h444;
rom[95572] = 12'h444;
rom[95573] = 12'h666;
rom[95574] = 12'h777;
rom[95575] = 12'h888;
rom[95576] = 12'h999;
rom[95577] = 12'haaa;
rom[95578] = 12'haaa;
rom[95579] = 12'haaa;
rom[95580] = 12'haaa;
rom[95581] = 12'h999;
rom[95582] = 12'h777;
rom[95583] = 12'h666;
rom[95584] = 12'h444;
rom[95585] = 12'h333;
rom[95586] = 12'h333;
rom[95587] = 12'h222;
rom[95588] = 12'h111;
rom[95589] = 12'h111;
rom[95590] = 12'h111;
rom[95591] = 12'h111;
rom[95592] = 12'h111;
rom[95593] = 12'h111;
rom[95594] = 12'h111;
rom[95595] = 12'h111;
rom[95596] = 12'h111;
rom[95597] = 12'h111;
rom[95598] = 12'h111;
rom[95599] = 12'h111;
rom[95600] = 12'hfff;
rom[95601] = 12'hfff;
rom[95602] = 12'hfff;
rom[95603] = 12'hfff;
rom[95604] = 12'hfff;
rom[95605] = 12'hfff;
rom[95606] = 12'hfff;
rom[95607] = 12'hfff;
rom[95608] = 12'hfff;
rom[95609] = 12'hfff;
rom[95610] = 12'hfff;
rom[95611] = 12'hfff;
rom[95612] = 12'hfff;
rom[95613] = 12'hfff;
rom[95614] = 12'hfff;
rom[95615] = 12'hfff;
rom[95616] = 12'hfff;
rom[95617] = 12'hfff;
rom[95618] = 12'hfff;
rom[95619] = 12'hfff;
rom[95620] = 12'hfff;
rom[95621] = 12'hfff;
rom[95622] = 12'hfff;
rom[95623] = 12'hfff;
rom[95624] = 12'hfff;
rom[95625] = 12'hfff;
rom[95626] = 12'hfff;
rom[95627] = 12'hfff;
rom[95628] = 12'hfff;
rom[95629] = 12'hfff;
rom[95630] = 12'hfff;
rom[95631] = 12'hfff;
rom[95632] = 12'hfff;
rom[95633] = 12'hfff;
rom[95634] = 12'hfff;
rom[95635] = 12'hfff;
rom[95636] = 12'hfff;
rom[95637] = 12'hfff;
rom[95638] = 12'hfff;
rom[95639] = 12'hfff;
rom[95640] = 12'hfff;
rom[95641] = 12'hfff;
rom[95642] = 12'hfff;
rom[95643] = 12'hfff;
rom[95644] = 12'hfff;
rom[95645] = 12'hfff;
rom[95646] = 12'hfff;
rom[95647] = 12'hfff;
rom[95648] = 12'hfff;
rom[95649] = 12'hfff;
rom[95650] = 12'hfff;
rom[95651] = 12'hfff;
rom[95652] = 12'hfff;
rom[95653] = 12'hfff;
rom[95654] = 12'hfff;
rom[95655] = 12'hfff;
rom[95656] = 12'hfff;
rom[95657] = 12'hfff;
rom[95658] = 12'hfff;
rom[95659] = 12'hfff;
rom[95660] = 12'hfff;
rom[95661] = 12'hfff;
rom[95662] = 12'hfff;
rom[95663] = 12'hfff;
rom[95664] = 12'hfff;
rom[95665] = 12'hfff;
rom[95666] = 12'hfff;
rom[95667] = 12'hfff;
rom[95668] = 12'hfff;
rom[95669] = 12'hfff;
rom[95670] = 12'hfff;
rom[95671] = 12'hfff;
rom[95672] = 12'hfff;
rom[95673] = 12'hfff;
rom[95674] = 12'hfff;
rom[95675] = 12'hfff;
rom[95676] = 12'hfff;
rom[95677] = 12'hfff;
rom[95678] = 12'hfff;
rom[95679] = 12'hfff;
rom[95680] = 12'hfff;
rom[95681] = 12'hfff;
rom[95682] = 12'hfff;
rom[95683] = 12'hfff;
rom[95684] = 12'hfff;
rom[95685] = 12'hfff;
rom[95686] = 12'hfff;
rom[95687] = 12'hfff;
rom[95688] = 12'hfff;
rom[95689] = 12'hfff;
rom[95690] = 12'hfff;
rom[95691] = 12'hfff;
rom[95692] = 12'hfff;
rom[95693] = 12'hfff;
rom[95694] = 12'hfff;
rom[95695] = 12'hfff;
rom[95696] = 12'hfff;
rom[95697] = 12'hfff;
rom[95698] = 12'hfff;
rom[95699] = 12'hfff;
rom[95700] = 12'hfff;
rom[95701] = 12'hfff;
rom[95702] = 12'hfff;
rom[95703] = 12'hfff;
rom[95704] = 12'hfff;
rom[95705] = 12'hfff;
rom[95706] = 12'hfff;
rom[95707] = 12'hfff;
rom[95708] = 12'hfff;
rom[95709] = 12'hfff;
rom[95710] = 12'hfff;
rom[95711] = 12'hfff;
rom[95712] = 12'hfff;
rom[95713] = 12'hfff;
rom[95714] = 12'hfff;
rom[95715] = 12'hfff;
rom[95716] = 12'hfff;
rom[95717] = 12'hfff;
rom[95718] = 12'hfff;
rom[95719] = 12'hfff;
rom[95720] = 12'hfff;
rom[95721] = 12'hfff;
rom[95722] = 12'hfff;
rom[95723] = 12'hfff;
rom[95724] = 12'hfff;
rom[95725] = 12'hfff;
rom[95726] = 12'hfff;
rom[95727] = 12'hfff;
rom[95728] = 12'hfff;
rom[95729] = 12'hfff;
rom[95730] = 12'hfff;
rom[95731] = 12'hfff;
rom[95732] = 12'hfff;
rom[95733] = 12'hfff;
rom[95734] = 12'hfff;
rom[95735] = 12'hfff;
rom[95736] = 12'hfff;
rom[95737] = 12'hfff;
rom[95738] = 12'hfff;
rom[95739] = 12'hfff;
rom[95740] = 12'heee;
rom[95741] = 12'heee;
rom[95742] = 12'heee;
rom[95743] = 12'heee;
rom[95744] = 12'hddd;
rom[95745] = 12'hddd;
rom[95746] = 12'hddd;
rom[95747] = 12'hccc;
rom[95748] = 12'hccc;
rom[95749] = 12'hccc;
rom[95750] = 12'hccc;
rom[95751] = 12'hccc;
rom[95752] = 12'hccc;
rom[95753] = 12'hccc;
rom[95754] = 12'hccc;
rom[95755] = 12'hccc;
rom[95756] = 12'hccc;
rom[95757] = 12'hccc;
rom[95758] = 12'hccc;
rom[95759] = 12'hccc;
rom[95760] = 12'hccc;
rom[95761] = 12'hccc;
rom[95762] = 12'hccc;
rom[95763] = 12'hccc;
rom[95764] = 12'hbbb;
rom[95765] = 12'hbbb;
rom[95766] = 12'hbbb;
rom[95767] = 12'hbbb;
rom[95768] = 12'haaa;
rom[95769] = 12'haaa;
rom[95770] = 12'haaa;
rom[95771] = 12'haaa;
rom[95772] = 12'haaa;
rom[95773] = 12'haaa;
rom[95774] = 12'haaa;
rom[95775] = 12'haaa;
rom[95776] = 12'h999;
rom[95777] = 12'h999;
rom[95778] = 12'h999;
rom[95779] = 12'h999;
rom[95780] = 12'h999;
rom[95781] = 12'h999;
rom[95782] = 12'h999;
rom[95783] = 12'h999;
rom[95784] = 12'h999;
rom[95785] = 12'h999;
rom[95786] = 12'h999;
rom[95787] = 12'h888;
rom[95788] = 12'h888;
rom[95789] = 12'h888;
rom[95790] = 12'h888;
rom[95791] = 12'h888;
rom[95792] = 12'h888;
rom[95793] = 12'h888;
rom[95794] = 12'h888;
rom[95795] = 12'h888;
rom[95796] = 12'h888;
rom[95797] = 12'h999;
rom[95798] = 12'h999;
rom[95799] = 12'h999;
rom[95800] = 12'h999;
rom[95801] = 12'h999;
rom[95802] = 12'h999;
rom[95803] = 12'h999;
rom[95804] = 12'h999;
rom[95805] = 12'h999;
rom[95806] = 12'h999;
rom[95807] = 12'h999;
rom[95808] = 12'h999;
rom[95809] = 12'h999;
rom[95810] = 12'h999;
rom[95811] = 12'h999;
rom[95812] = 12'h999;
rom[95813] = 12'h888;
rom[95814] = 12'h888;
rom[95815] = 12'h888;
rom[95816] = 12'h777;
rom[95817] = 12'h777;
rom[95818] = 12'h666;
rom[95819] = 12'h666;
rom[95820] = 12'h777;
rom[95821] = 12'h777;
rom[95822] = 12'h777;
rom[95823] = 12'h666;
rom[95824] = 12'h666;
rom[95825] = 12'h666;
rom[95826] = 12'h666;
rom[95827] = 12'h666;
rom[95828] = 12'h777;
rom[95829] = 12'h777;
rom[95830] = 12'h777;
rom[95831] = 12'h777;
rom[95832] = 12'h777;
rom[95833] = 12'h888;
rom[95834] = 12'h888;
rom[95835] = 12'h888;
rom[95836] = 12'h888;
rom[95837] = 12'h999;
rom[95838] = 12'h999;
rom[95839] = 12'h888;
rom[95840] = 12'h888;
rom[95841] = 12'h888;
rom[95842] = 12'h777;
rom[95843] = 12'h777;
rom[95844] = 12'h666;
rom[95845] = 12'h666;
rom[95846] = 12'h666;
rom[95847] = 12'h666;
rom[95848] = 12'h555;
rom[95849] = 12'h555;
rom[95850] = 12'h555;
rom[95851] = 12'h555;
rom[95852] = 12'h555;
rom[95853] = 12'h555;
rom[95854] = 12'h555;
rom[95855] = 12'h555;
rom[95856] = 12'h555;
rom[95857] = 12'h555;
rom[95858] = 12'h666;
rom[95859] = 12'h666;
rom[95860] = 12'h666;
rom[95861] = 12'h666;
rom[95862] = 12'h777;
rom[95863] = 12'h777;
rom[95864] = 12'h888;
rom[95865] = 12'h888;
rom[95866] = 12'h999;
rom[95867] = 12'h999;
rom[95868] = 12'h999;
rom[95869] = 12'h888;
rom[95870] = 12'h888;
rom[95871] = 12'h888;
rom[95872] = 12'h888;
rom[95873] = 12'h888;
rom[95874] = 12'h777;
rom[95875] = 12'h777;
rom[95876] = 12'h777;
rom[95877] = 12'h777;
rom[95878] = 12'h777;
rom[95879] = 12'h777;
rom[95880] = 12'h888;
rom[95881] = 12'h888;
rom[95882] = 12'h888;
rom[95883] = 12'h888;
rom[95884] = 12'h888;
rom[95885] = 12'h888;
rom[95886] = 12'h888;
rom[95887] = 12'h888;
rom[95888] = 12'h999;
rom[95889] = 12'hbbb;
rom[95890] = 12'hccc;
rom[95891] = 12'hddd;
rom[95892] = 12'heee;
rom[95893] = 12'hfff;
rom[95894] = 12'heee;
rom[95895] = 12'hddd;
rom[95896] = 12'hccc;
rom[95897] = 12'hbbb;
rom[95898] = 12'haaa;
rom[95899] = 12'h999;
rom[95900] = 12'h888;
rom[95901] = 12'h777;
rom[95902] = 12'h666;
rom[95903] = 12'h666;
rom[95904] = 12'h666;
rom[95905] = 12'h666;
rom[95906] = 12'h666;
rom[95907] = 12'h777;
rom[95908] = 12'h888;
rom[95909] = 12'haaa;
rom[95910] = 12'hccc;
rom[95911] = 12'hddd;
rom[95912] = 12'hfff;
rom[95913] = 12'hfff;
rom[95914] = 12'hfff;
rom[95915] = 12'hfff;
rom[95916] = 12'hfff;
rom[95917] = 12'hfff;
rom[95918] = 12'hddd;
rom[95919] = 12'hbbb;
rom[95920] = 12'h888;
rom[95921] = 12'h777;
rom[95922] = 12'h555;
rom[95923] = 12'h444;
rom[95924] = 12'h444;
rom[95925] = 12'h444;
rom[95926] = 12'h333;
rom[95927] = 12'h333;
rom[95928] = 12'h333;
rom[95929] = 12'h333;
rom[95930] = 12'h333;
rom[95931] = 12'h333;
rom[95932] = 12'h222;
rom[95933] = 12'h222;
rom[95934] = 12'h222;
rom[95935] = 12'h222;
rom[95936] = 12'h222;
rom[95937] = 12'h222;
rom[95938] = 12'h222;
rom[95939] = 12'h222;
rom[95940] = 12'h222;
rom[95941] = 12'h222;
rom[95942] = 12'h111;
rom[95943] = 12'h111;
rom[95944] = 12'h111;
rom[95945] = 12'h111;
rom[95946] = 12'h  0;
rom[95947] = 12'h  0;
rom[95948] = 12'h  0;
rom[95949] = 12'h  0;
rom[95950] = 12'h111;
rom[95951] = 12'h111;
rom[95952] = 12'h111;
rom[95953] = 12'h111;
rom[95954] = 12'h111;
rom[95955] = 12'h111;
rom[95956] = 12'h111;
rom[95957] = 12'h111;
rom[95958] = 12'h111;
rom[95959] = 12'h222;
rom[95960] = 12'h111;
rom[95961] = 12'h222;
rom[95962] = 12'h222;
rom[95963] = 12'h222;
rom[95964] = 12'h222;
rom[95965] = 12'h222;
rom[95966] = 12'h222;
rom[95967] = 12'h222;
rom[95968] = 12'h222;
rom[95969] = 12'h222;
rom[95970] = 12'h333;
rom[95971] = 12'h333;
rom[95972] = 12'h333;
rom[95973] = 12'h444;
rom[95974] = 12'h555;
rom[95975] = 12'h666;
rom[95976] = 12'h999;
rom[95977] = 12'h999;
rom[95978] = 12'h888;
rom[95979] = 12'h888;
rom[95980] = 12'h999;
rom[95981] = 12'haaa;
rom[95982] = 12'h999;
rom[95983] = 12'h888;
rom[95984] = 12'h777;
rom[95985] = 12'h666;
rom[95986] = 12'h555;
rom[95987] = 12'h333;
rom[95988] = 12'h222;
rom[95989] = 12'h222;
rom[95990] = 12'h111;
rom[95991] = 12'h111;
rom[95992] = 12'h111;
rom[95993] = 12'h111;
rom[95994] = 12'h111;
rom[95995] = 12'h111;
rom[95996] = 12'h111;
rom[95997] = 12'h111;
rom[95998] = 12'h111;
rom[95999] = 12'h111;
rom[96000] = 12'hfff;
rom[96001] = 12'hfff;
rom[96002] = 12'hfff;
rom[96003] = 12'hfff;
rom[96004] = 12'hfff;
rom[96005] = 12'hfff;
rom[96006] = 12'hfff;
rom[96007] = 12'hfff;
rom[96008] = 12'hfff;
rom[96009] = 12'hfff;
rom[96010] = 12'hfff;
rom[96011] = 12'hfff;
rom[96012] = 12'hfff;
rom[96013] = 12'hfff;
rom[96014] = 12'hfff;
rom[96015] = 12'hfff;
rom[96016] = 12'hfff;
rom[96017] = 12'hfff;
rom[96018] = 12'hfff;
rom[96019] = 12'hfff;
rom[96020] = 12'hfff;
rom[96021] = 12'hfff;
rom[96022] = 12'hfff;
rom[96023] = 12'hfff;
rom[96024] = 12'hfff;
rom[96025] = 12'hfff;
rom[96026] = 12'hfff;
rom[96027] = 12'hfff;
rom[96028] = 12'hfff;
rom[96029] = 12'hfff;
rom[96030] = 12'hfff;
rom[96031] = 12'hfff;
rom[96032] = 12'hfff;
rom[96033] = 12'hfff;
rom[96034] = 12'hfff;
rom[96035] = 12'hfff;
rom[96036] = 12'hfff;
rom[96037] = 12'hfff;
rom[96038] = 12'hfff;
rom[96039] = 12'hfff;
rom[96040] = 12'hfff;
rom[96041] = 12'hfff;
rom[96042] = 12'hfff;
rom[96043] = 12'hfff;
rom[96044] = 12'hfff;
rom[96045] = 12'hfff;
rom[96046] = 12'hfff;
rom[96047] = 12'hfff;
rom[96048] = 12'hfff;
rom[96049] = 12'hfff;
rom[96050] = 12'hfff;
rom[96051] = 12'hfff;
rom[96052] = 12'hfff;
rom[96053] = 12'hfff;
rom[96054] = 12'hfff;
rom[96055] = 12'hfff;
rom[96056] = 12'hfff;
rom[96057] = 12'hfff;
rom[96058] = 12'hfff;
rom[96059] = 12'hfff;
rom[96060] = 12'hfff;
rom[96061] = 12'hfff;
rom[96062] = 12'hfff;
rom[96063] = 12'hfff;
rom[96064] = 12'hfff;
rom[96065] = 12'hfff;
rom[96066] = 12'hfff;
rom[96067] = 12'hfff;
rom[96068] = 12'hfff;
rom[96069] = 12'hfff;
rom[96070] = 12'hfff;
rom[96071] = 12'hfff;
rom[96072] = 12'hfff;
rom[96073] = 12'hfff;
rom[96074] = 12'hfff;
rom[96075] = 12'hfff;
rom[96076] = 12'hfff;
rom[96077] = 12'hfff;
rom[96078] = 12'hfff;
rom[96079] = 12'hfff;
rom[96080] = 12'hfff;
rom[96081] = 12'hfff;
rom[96082] = 12'hfff;
rom[96083] = 12'hfff;
rom[96084] = 12'hfff;
rom[96085] = 12'hfff;
rom[96086] = 12'hfff;
rom[96087] = 12'hfff;
rom[96088] = 12'hfff;
rom[96089] = 12'hfff;
rom[96090] = 12'hfff;
rom[96091] = 12'hfff;
rom[96092] = 12'hfff;
rom[96093] = 12'hfff;
rom[96094] = 12'hfff;
rom[96095] = 12'hfff;
rom[96096] = 12'hfff;
rom[96097] = 12'hfff;
rom[96098] = 12'hfff;
rom[96099] = 12'hfff;
rom[96100] = 12'hfff;
rom[96101] = 12'hfff;
rom[96102] = 12'hfff;
rom[96103] = 12'hfff;
rom[96104] = 12'hfff;
rom[96105] = 12'hfff;
rom[96106] = 12'hfff;
rom[96107] = 12'hfff;
rom[96108] = 12'hfff;
rom[96109] = 12'hfff;
rom[96110] = 12'hfff;
rom[96111] = 12'hfff;
rom[96112] = 12'hfff;
rom[96113] = 12'hfff;
rom[96114] = 12'hfff;
rom[96115] = 12'hfff;
rom[96116] = 12'hfff;
rom[96117] = 12'hfff;
rom[96118] = 12'hfff;
rom[96119] = 12'hfff;
rom[96120] = 12'hfff;
rom[96121] = 12'hfff;
rom[96122] = 12'hfff;
rom[96123] = 12'hfff;
rom[96124] = 12'hfff;
rom[96125] = 12'hfff;
rom[96126] = 12'hfff;
rom[96127] = 12'hfff;
rom[96128] = 12'hfff;
rom[96129] = 12'hfff;
rom[96130] = 12'hfff;
rom[96131] = 12'hfff;
rom[96132] = 12'hfff;
rom[96133] = 12'hfff;
rom[96134] = 12'hfff;
rom[96135] = 12'hfff;
rom[96136] = 12'hfff;
rom[96137] = 12'hfff;
rom[96138] = 12'hfff;
rom[96139] = 12'hfff;
rom[96140] = 12'hfff;
rom[96141] = 12'heee;
rom[96142] = 12'heee;
rom[96143] = 12'heee;
rom[96144] = 12'hddd;
rom[96145] = 12'hddd;
rom[96146] = 12'hddd;
rom[96147] = 12'hddd;
rom[96148] = 12'hddd;
rom[96149] = 12'hddd;
rom[96150] = 12'hddd;
rom[96151] = 12'hccc;
rom[96152] = 12'hddd;
rom[96153] = 12'hddd;
rom[96154] = 12'hccc;
rom[96155] = 12'hccc;
rom[96156] = 12'hccc;
rom[96157] = 12'hccc;
rom[96158] = 12'hccc;
rom[96159] = 12'hccc;
rom[96160] = 12'hccc;
rom[96161] = 12'hccc;
rom[96162] = 12'hccc;
rom[96163] = 12'hccc;
rom[96164] = 12'hccc;
rom[96165] = 12'hccc;
rom[96166] = 12'hccc;
rom[96167] = 12'hccc;
rom[96168] = 12'hbbb;
rom[96169] = 12'hbbb;
rom[96170] = 12'haaa;
rom[96171] = 12'haaa;
rom[96172] = 12'haaa;
rom[96173] = 12'haaa;
rom[96174] = 12'haaa;
rom[96175] = 12'haaa;
rom[96176] = 12'h999;
rom[96177] = 12'h999;
rom[96178] = 12'h999;
rom[96179] = 12'h999;
rom[96180] = 12'h999;
rom[96181] = 12'h999;
rom[96182] = 12'h999;
rom[96183] = 12'h999;
rom[96184] = 12'h999;
rom[96185] = 12'h999;
rom[96186] = 12'h999;
rom[96187] = 12'h999;
rom[96188] = 12'h999;
rom[96189] = 12'h999;
rom[96190] = 12'h999;
rom[96191] = 12'h999;
rom[96192] = 12'h999;
rom[96193] = 12'h999;
rom[96194] = 12'h999;
rom[96195] = 12'h999;
rom[96196] = 12'h999;
rom[96197] = 12'h999;
rom[96198] = 12'h999;
rom[96199] = 12'h999;
rom[96200] = 12'h999;
rom[96201] = 12'h999;
rom[96202] = 12'h999;
rom[96203] = 12'h999;
rom[96204] = 12'h999;
rom[96205] = 12'h999;
rom[96206] = 12'h999;
rom[96207] = 12'h999;
rom[96208] = 12'h999;
rom[96209] = 12'h999;
rom[96210] = 12'h999;
rom[96211] = 12'h999;
rom[96212] = 12'h999;
rom[96213] = 12'h999;
rom[96214] = 12'h999;
rom[96215] = 12'h999;
rom[96216] = 12'h888;
rom[96217] = 12'h888;
rom[96218] = 12'h888;
rom[96219] = 12'h777;
rom[96220] = 12'h777;
rom[96221] = 12'h777;
rom[96222] = 12'h777;
rom[96223] = 12'h777;
rom[96224] = 12'h777;
rom[96225] = 12'h777;
rom[96226] = 12'h777;
rom[96227] = 12'h777;
rom[96228] = 12'h777;
rom[96229] = 12'h777;
rom[96230] = 12'h777;
rom[96231] = 12'h777;
rom[96232] = 12'h888;
rom[96233] = 12'h888;
rom[96234] = 12'h888;
rom[96235] = 12'h999;
rom[96236] = 12'h999;
rom[96237] = 12'h999;
rom[96238] = 12'h999;
rom[96239] = 12'h999;
rom[96240] = 12'h888;
rom[96241] = 12'h888;
rom[96242] = 12'h888;
rom[96243] = 12'h777;
rom[96244] = 12'h777;
rom[96245] = 12'h666;
rom[96246] = 12'h777;
rom[96247] = 12'h777;
rom[96248] = 12'h666;
rom[96249] = 12'h666;
rom[96250] = 12'h666;
rom[96251] = 12'h666;
rom[96252] = 12'h666;
rom[96253] = 12'h666;
rom[96254] = 12'h666;
rom[96255] = 12'h666;
rom[96256] = 12'h666;
rom[96257] = 12'h666;
rom[96258] = 12'h777;
rom[96259] = 12'h777;
rom[96260] = 12'h777;
rom[96261] = 12'h888;
rom[96262] = 12'h888;
rom[96263] = 12'h888;
rom[96264] = 12'h999;
rom[96265] = 12'h999;
rom[96266] = 12'h999;
rom[96267] = 12'h999;
rom[96268] = 12'h999;
rom[96269] = 12'h888;
rom[96270] = 12'h888;
rom[96271] = 12'h888;
rom[96272] = 12'h888;
rom[96273] = 12'h888;
rom[96274] = 12'h888;
rom[96275] = 12'h777;
rom[96276] = 12'h777;
rom[96277] = 12'h777;
rom[96278] = 12'h777;
rom[96279] = 12'h777;
rom[96280] = 12'h888;
rom[96281] = 12'h888;
rom[96282] = 12'h888;
rom[96283] = 12'h888;
rom[96284] = 12'h888;
rom[96285] = 12'h888;
rom[96286] = 12'h999;
rom[96287] = 12'h999;
rom[96288] = 12'hbbb;
rom[96289] = 12'hccc;
rom[96290] = 12'heee;
rom[96291] = 12'hfff;
rom[96292] = 12'heee;
rom[96293] = 12'heee;
rom[96294] = 12'hddd;
rom[96295] = 12'hddd;
rom[96296] = 12'hccc;
rom[96297] = 12'hccc;
rom[96298] = 12'hbbb;
rom[96299] = 12'haaa;
rom[96300] = 12'h888;
rom[96301] = 12'h777;
rom[96302] = 12'h777;
rom[96303] = 12'h777;
rom[96304] = 12'h666;
rom[96305] = 12'h555;
rom[96306] = 12'h555;
rom[96307] = 12'h666;
rom[96308] = 12'h666;
rom[96309] = 12'h666;
rom[96310] = 12'h888;
rom[96311] = 12'h999;
rom[96312] = 12'hccc;
rom[96313] = 12'hccc;
rom[96314] = 12'heee;
rom[96315] = 12'hfff;
rom[96316] = 12'hfff;
rom[96317] = 12'hfff;
rom[96318] = 12'hfff;
rom[96319] = 12'hfff;
rom[96320] = 12'hccc;
rom[96321] = 12'haaa;
rom[96322] = 12'h888;
rom[96323] = 12'h666;
rom[96324] = 12'h555;
rom[96325] = 12'h444;
rom[96326] = 12'h444;
rom[96327] = 12'h444;
rom[96328] = 12'h333;
rom[96329] = 12'h333;
rom[96330] = 12'h222;
rom[96331] = 12'h333;
rom[96332] = 12'h333;
rom[96333] = 12'h222;
rom[96334] = 12'h111;
rom[96335] = 12'h111;
rom[96336] = 12'h111;
rom[96337] = 12'h222;
rom[96338] = 12'h222;
rom[96339] = 12'h222;
rom[96340] = 12'h222;
rom[96341] = 12'h333;
rom[96342] = 12'h222;
rom[96343] = 12'h111;
rom[96344] = 12'h  0;
rom[96345] = 12'h  0;
rom[96346] = 12'h  0;
rom[96347] = 12'h  0;
rom[96348] = 12'h111;
rom[96349] = 12'h111;
rom[96350] = 12'h111;
rom[96351] = 12'h  0;
rom[96352] = 12'h111;
rom[96353] = 12'h111;
rom[96354] = 12'h111;
rom[96355] = 12'h111;
rom[96356] = 12'h111;
rom[96357] = 12'h111;
rom[96358] = 12'h111;
rom[96359] = 12'h111;
rom[96360] = 12'h222;
rom[96361] = 12'h222;
rom[96362] = 12'h222;
rom[96363] = 12'h222;
rom[96364] = 12'h222;
rom[96365] = 12'h222;
rom[96366] = 12'h222;
rom[96367] = 12'h222;
rom[96368] = 12'h222;
rom[96369] = 12'h222;
rom[96370] = 12'h222;
rom[96371] = 12'h333;
rom[96372] = 12'h333;
rom[96373] = 12'h333;
rom[96374] = 12'h444;
rom[96375] = 12'h444;
rom[96376] = 12'h666;
rom[96377] = 12'h777;
rom[96378] = 12'h888;
rom[96379] = 12'h888;
rom[96380] = 12'h888;
rom[96381] = 12'h777;
rom[96382] = 12'h888;
rom[96383] = 12'h888;
rom[96384] = 12'h888;
rom[96385] = 12'h777;
rom[96386] = 12'h777;
rom[96387] = 12'h666;
rom[96388] = 12'h555;
rom[96389] = 12'h444;
rom[96390] = 12'h333;
rom[96391] = 12'h222;
rom[96392] = 12'h111;
rom[96393] = 12'h111;
rom[96394] = 12'h111;
rom[96395] = 12'h111;
rom[96396] = 12'h111;
rom[96397] = 12'h111;
rom[96398] = 12'h111;
rom[96399] = 12'h111;
rom[96400] = 12'hfff;
rom[96401] = 12'hfff;
rom[96402] = 12'hfff;
rom[96403] = 12'hfff;
rom[96404] = 12'hfff;
rom[96405] = 12'hfff;
rom[96406] = 12'hfff;
rom[96407] = 12'hfff;
rom[96408] = 12'hfff;
rom[96409] = 12'hfff;
rom[96410] = 12'hfff;
rom[96411] = 12'hfff;
rom[96412] = 12'hfff;
rom[96413] = 12'hfff;
rom[96414] = 12'hfff;
rom[96415] = 12'hfff;
rom[96416] = 12'hfff;
rom[96417] = 12'hfff;
rom[96418] = 12'hfff;
rom[96419] = 12'hfff;
rom[96420] = 12'hfff;
rom[96421] = 12'hfff;
rom[96422] = 12'hfff;
rom[96423] = 12'hfff;
rom[96424] = 12'hfff;
rom[96425] = 12'hfff;
rom[96426] = 12'hfff;
rom[96427] = 12'hfff;
rom[96428] = 12'hfff;
rom[96429] = 12'hfff;
rom[96430] = 12'hfff;
rom[96431] = 12'hfff;
rom[96432] = 12'hfff;
rom[96433] = 12'hfff;
rom[96434] = 12'hfff;
rom[96435] = 12'hfff;
rom[96436] = 12'hfff;
rom[96437] = 12'hfff;
rom[96438] = 12'hfff;
rom[96439] = 12'hfff;
rom[96440] = 12'hfff;
rom[96441] = 12'hfff;
rom[96442] = 12'hfff;
rom[96443] = 12'hfff;
rom[96444] = 12'hfff;
rom[96445] = 12'hfff;
rom[96446] = 12'hfff;
rom[96447] = 12'hfff;
rom[96448] = 12'hfff;
rom[96449] = 12'hfff;
rom[96450] = 12'hfff;
rom[96451] = 12'hfff;
rom[96452] = 12'hfff;
rom[96453] = 12'hfff;
rom[96454] = 12'hfff;
rom[96455] = 12'hfff;
rom[96456] = 12'hfff;
rom[96457] = 12'hfff;
rom[96458] = 12'hfff;
rom[96459] = 12'hfff;
rom[96460] = 12'hfff;
rom[96461] = 12'hfff;
rom[96462] = 12'hfff;
rom[96463] = 12'hfff;
rom[96464] = 12'hfff;
rom[96465] = 12'hfff;
rom[96466] = 12'hfff;
rom[96467] = 12'hfff;
rom[96468] = 12'hfff;
rom[96469] = 12'hfff;
rom[96470] = 12'hfff;
rom[96471] = 12'hfff;
rom[96472] = 12'hfff;
rom[96473] = 12'hfff;
rom[96474] = 12'hfff;
rom[96475] = 12'hfff;
rom[96476] = 12'hfff;
rom[96477] = 12'hfff;
rom[96478] = 12'hfff;
rom[96479] = 12'hfff;
rom[96480] = 12'hfff;
rom[96481] = 12'hfff;
rom[96482] = 12'hfff;
rom[96483] = 12'hfff;
rom[96484] = 12'hfff;
rom[96485] = 12'hfff;
rom[96486] = 12'hfff;
rom[96487] = 12'hfff;
rom[96488] = 12'hfff;
rom[96489] = 12'hfff;
rom[96490] = 12'hfff;
rom[96491] = 12'hfff;
rom[96492] = 12'hfff;
rom[96493] = 12'hfff;
rom[96494] = 12'hfff;
rom[96495] = 12'hfff;
rom[96496] = 12'hfff;
rom[96497] = 12'hfff;
rom[96498] = 12'hfff;
rom[96499] = 12'hfff;
rom[96500] = 12'hfff;
rom[96501] = 12'hfff;
rom[96502] = 12'hfff;
rom[96503] = 12'hfff;
rom[96504] = 12'hfff;
rom[96505] = 12'hfff;
rom[96506] = 12'hfff;
rom[96507] = 12'hfff;
rom[96508] = 12'hfff;
rom[96509] = 12'hfff;
rom[96510] = 12'hfff;
rom[96511] = 12'hfff;
rom[96512] = 12'hfff;
rom[96513] = 12'hfff;
rom[96514] = 12'hfff;
rom[96515] = 12'hfff;
rom[96516] = 12'hfff;
rom[96517] = 12'hfff;
rom[96518] = 12'hfff;
rom[96519] = 12'hfff;
rom[96520] = 12'hfff;
rom[96521] = 12'hfff;
rom[96522] = 12'hfff;
rom[96523] = 12'hfff;
rom[96524] = 12'hfff;
rom[96525] = 12'hfff;
rom[96526] = 12'hfff;
rom[96527] = 12'hfff;
rom[96528] = 12'hfff;
rom[96529] = 12'hfff;
rom[96530] = 12'hfff;
rom[96531] = 12'hfff;
rom[96532] = 12'hfff;
rom[96533] = 12'hfff;
rom[96534] = 12'hfff;
rom[96535] = 12'hfff;
rom[96536] = 12'hfff;
rom[96537] = 12'hfff;
rom[96538] = 12'hfff;
rom[96539] = 12'hfff;
rom[96540] = 12'hfff;
rom[96541] = 12'hfff;
rom[96542] = 12'heee;
rom[96543] = 12'heee;
rom[96544] = 12'heee;
rom[96545] = 12'heee;
rom[96546] = 12'hddd;
rom[96547] = 12'hddd;
rom[96548] = 12'hddd;
rom[96549] = 12'hddd;
rom[96550] = 12'hddd;
rom[96551] = 12'hddd;
rom[96552] = 12'hddd;
rom[96553] = 12'hddd;
rom[96554] = 12'hddd;
rom[96555] = 12'hccc;
rom[96556] = 12'hccc;
rom[96557] = 12'hccc;
rom[96558] = 12'hccc;
rom[96559] = 12'hccc;
rom[96560] = 12'hccc;
rom[96561] = 12'hccc;
rom[96562] = 12'hccc;
rom[96563] = 12'hccc;
rom[96564] = 12'hccc;
rom[96565] = 12'hccc;
rom[96566] = 12'hccc;
rom[96567] = 12'hccc;
rom[96568] = 12'hbbb;
rom[96569] = 12'hbbb;
rom[96570] = 12'hbbb;
rom[96571] = 12'haaa;
rom[96572] = 12'haaa;
rom[96573] = 12'haaa;
rom[96574] = 12'haaa;
rom[96575] = 12'haaa;
rom[96576] = 12'h999;
rom[96577] = 12'h999;
rom[96578] = 12'h999;
rom[96579] = 12'h999;
rom[96580] = 12'h999;
rom[96581] = 12'h999;
rom[96582] = 12'h999;
rom[96583] = 12'h999;
rom[96584] = 12'h999;
rom[96585] = 12'h999;
rom[96586] = 12'h999;
rom[96587] = 12'h999;
rom[96588] = 12'h999;
rom[96589] = 12'h999;
rom[96590] = 12'h999;
rom[96591] = 12'h999;
rom[96592] = 12'h999;
rom[96593] = 12'h999;
rom[96594] = 12'h999;
rom[96595] = 12'h999;
rom[96596] = 12'h999;
rom[96597] = 12'h999;
rom[96598] = 12'h999;
rom[96599] = 12'h999;
rom[96600] = 12'h999;
rom[96601] = 12'h999;
rom[96602] = 12'h999;
rom[96603] = 12'h999;
rom[96604] = 12'h999;
rom[96605] = 12'h999;
rom[96606] = 12'haaa;
rom[96607] = 12'haaa;
rom[96608] = 12'h999;
rom[96609] = 12'haaa;
rom[96610] = 12'haaa;
rom[96611] = 12'haaa;
rom[96612] = 12'haaa;
rom[96613] = 12'h999;
rom[96614] = 12'h999;
rom[96615] = 12'h999;
rom[96616] = 12'h999;
rom[96617] = 12'h888;
rom[96618] = 12'h888;
rom[96619] = 12'h888;
rom[96620] = 12'h888;
rom[96621] = 12'h777;
rom[96622] = 12'h777;
rom[96623] = 12'h888;
rom[96624] = 12'h777;
rom[96625] = 12'h777;
rom[96626] = 12'h777;
rom[96627] = 12'h777;
rom[96628] = 12'h777;
rom[96629] = 12'h777;
rom[96630] = 12'h888;
rom[96631] = 12'h888;
rom[96632] = 12'h888;
rom[96633] = 12'h888;
rom[96634] = 12'h888;
rom[96635] = 12'h999;
rom[96636] = 12'h999;
rom[96637] = 12'h999;
rom[96638] = 12'h999;
rom[96639] = 12'h999;
rom[96640] = 12'h999;
rom[96641] = 12'h999;
rom[96642] = 12'h888;
rom[96643] = 12'h888;
rom[96644] = 12'h777;
rom[96645] = 12'h777;
rom[96646] = 12'h777;
rom[96647] = 12'h777;
rom[96648] = 12'h777;
rom[96649] = 12'h777;
rom[96650] = 12'h777;
rom[96651] = 12'h777;
rom[96652] = 12'h777;
rom[96653] = 12'h777;
rom[96654] = 12'h777;
rom[96655] = 12'h666;
rom[96656] = 12'h777;
rom[96657] = 12'h777;
rom[96658] = 12'h777;
rom[96659] = 12'h888;
rom[96660] = 12'h888;
rom[96661] = 12'h888;
rom[96662] = 12'h888;
rom[96663] = 12'h999;
rom[96664] = 12'h999;
rom[96665] = 12'h999;
rom[96666] = 12'h999;
rom[96667] = 12'h999;
rom[96668] = 12'h999;
rom[96669] = 12'h888;
rom[96670] = 12'h888;
rom[96671] = 12'h888;
rom[96672] = 12'h888;
rom[96673] = 12'h888;
rom[96674] = 12'h888;
rom[96675] = 12'h888;
rom[96676] = 12'h777;
rom[96677] = 12'h777;
rom[96678] = 12'h777;
rom[96679] = 12'h777;
rom[96680] = 12'h777;
rom[96681] = 12'h777;
rom[96682] = 12'h777;
rom[96683] = 12'h888;
rom[96684] = 12'h888;
rom[96685] = 12'h999;
rom[96686] = 12'haaa;
rom[96687] = 12'haaa;
rom[96688] = 12'hccc;
rom[96689] = 12'hddd;
rom[96690] = 12'heee;
rom[96691] = 12'hfff;
rom[96692] = 12'heee;
rom[96693] = 12'hddd;
rom[96694] = 12'hddd;
rom[96695] = 12'hccc;
rom[96696] = 12'hddd;
rom[96697] = 12'hddd;
rom[96698] = 12'hddd;
rom[96699] = 12'hccc;
rom[96700] = 12'haaa;
rom[96701] = 12'h888;
rom[96702] = 12'h777;
rom[96703] = 12'h666;
rom[96704] = 12'h666;
rom[96705] = 12'h666;
rom[96706] = 12'h666;
rom[96707] = 12'h555;
rom[96708] = 12'h555;
rom[96709] = 12'h666;
rom[96710] = 12'h777;
rom[96711] = 12'h777;
rom[96712] = 12'h999;
rom[96713] = 12'haaa;
rom[96714] = 12'hbbb;
rom[96715] = 12'hccc;
rom[96716] = 12'hddd;
rom[96717] = 12'heee;
rom[96718] = 12'hfff;
rom[96719] = 12'hfff;
rom[96720] = 12'hfff;
rom[96721] = 12'heee;
rom[96722] = 12'hccc;
rom[96723] = 12'haaa;
rom[96724] = 12'h777;
rom[96725] = 12'h666;
rom[96726] = 12'h555;
rom[96727] = 12'h444;
rom[96728] = 12'h333;
rom[96729] = 12'h333;
rom[96730] = 12'h222;
rom[96731] = 12'h222;
rom[96732] = 12'h222;
rom[96733] = 12'h222;
rom[96734] = 12'h222;
rom[96735] = 12'h222;
rom[96736] = 12'h111;
rom[96737] = 12'h222;
rom[96738] = 12'h111;
rom[96739] = 12'h111;
rom[96740] = 12'h222;
rom[96741] = 12'h222;
rom[96742] = 12'h222;
rom[96743] = 12'h222;
rom[96744] = 12'h111;
rom[96745] = 12'h111;
rom[96746] = 12'h  0;
rom[96747] = 12'h  0;
rom[96748] = 12'h111;
rom[96749] = 12'h111;
rom[96750] = 12'h111;
rom[96751] = 12'h111;
rom[96752] = 12'h111;
rom[96753] = 12'h111;
rom[96754] = 12'h111;
rom[96755] = 12'h111;
rom[96756] = 12'h111;
rom[96757] = 12'h111;
rom[96758] = 12'h111;
rom[96759] = 12'h111;
rom[96760] = 12'h111;
rom[96761] = 12'h111;
rom[96762] = 12'h111;
rom[96763] = 12'h111;
rom[96764] = 12'h111;
rom[96765] = 12'h111;
rom[96766] = 12'h111;
rom[96767] = 12'h111;
rom[96768] = 12'h222;
rom[96769] = 12'h222;
rom[96770] = 12'h222;
rom[96771] = 12'h222;
rom[96772] = 12'h222;
rom[96773] = 12'h222;
rom[96774] = 12'h333;
rom[96775] = 12'h333;
rom[96776] = 12'h444;
rom[96777] = 12'h555;
rom[96778] = 12'h666;
rom[96779] = 12'h777;
rom[96780] = 12'h777;
rom[96781] = 12'h777;
rom[96782] = 12'h666;
rom[96783] = 12'h666;
rom[96784] = 12'h777;
rom[96785] = 12'h777;
rom[96786] = 12'h777;
rom[96787] = 12'h777;
rom[96788] = 12'h777;
rom[96789] = 12'h666;
rom[96790] = 12'h555;
rom[96791] = 12'h444;
rom[96792] = 12'h333;
rom[96793] = 12'h333;
rom[96794] = 12'h222;
rom[96795] = 12'h111;
rom[96796] = 12'h111;
rom[96797] = 12'h111;
rom[96798] = 12'h111;
rom[96799] = 12'h111;
rom[96800] = 12'hfff;
rom[96801] = 12'hfff;
rom[96802] = 12'hfff;
rom[96803] = 12'hfff;
rom[96804] = 12'hfff;
rom[96805] = 12'hfff;
rom[96806] = 12'hfff;
rom[96807] = 12'hfff;
rom[96808] = 12'hfff;
rom[96809] = 12'hfff;
rom[96810] = 12'hfff;
rom[96811] = 12'hfff;
rom[96812] = 12'hfff;
rom[96813] = 12'hfff;
rom[96814] = 12'hfff;
rom[96815] = 12'hfff;
rom[96816] = 12'hfff;
rom[96817] = 12'hfff;
rom[96818] = 12'hfff;
rom[96819] = 12'hfff;
rom[96820] = 12'hfff;
rom[96821] = 12'hfff;
rom[96822] = 12'hfff;
rom[96823] = 12'hfff;
rom[96824] = 12'hfff;
rom[96825] = 12'hfff;
rom[96826] = 12'hfff;
rom[96827] = 12'hfff;
rom[96828] = 12'hfff;
rom[96829] = 12'hfff;
rom[96830] = 12'hfff;
rom[96831] = 12'hfff;
rom[96832] = 12'hfff;
rom[96833] = 12'hfff;
rom[96834] = 12'hfff;
rom[96835] = 12'hfff;
rom[96836] = 12'hfff;
rom[96837] = 12'hfff;
rom[96838] = 12'hfff;
rom[96839] = 12'hfff;
rom[96840] = 12'hfff;
rom[96841] = 12'hfff;
rom[96842] = 12'hfff;
rom[96843] = 12'hfff;
rom[96844] = 12'hfff;
rom[96845] = 12'hfff;
rom[96846] = 12'hfff;
rom[96847] = 12'hfff;
rom[96848] = 12'hfff;
rom[96849] = 12'hfff;
rom[96850] = 12'hfff;
rom[96851] = 12'hfff;
rom[96852] = 12'hfff;
rom[96853] = 12'hfff;
rom[96854] = 12'hfff;
rom[96855] = 12'hfff;
rom[96856] = 12'hfff;
rom[96857] = 12'hfff;
rom[96858] = 12'hfff;
rom[96859] = 12'hfff;
rom[96860] = 12'hfff;
rom[96861] = 12'hfff;
rom[96862] = 12'hfff;
rom[96863] = 12'hfff;
rom[96864] = 12'hfff;
rom[96865] = 12'hfff;
rom[96866] = 12'hfff;
rom[96867] = 12'hfff;
rom[96868] = 12'hfff;
rom[96869] = 12'hfff;
rom[96870] = 12'hfff;
rom[96871] = 12'hfff;
rom[96872] = 12'hfff;
rom[96873] = 12'hfff;
rom[96874] = 12'hfff;
rom[96875] = 12'hfff;
rom[96876] = 12'hfff;
rom[96877] = 12'hfff;
rom[96878] = 12'hfff;
rom[96879] = 12'hfff;
rom[96880] = 12'hfff;
rom[96881] = 12'hfff;
rom[96882] = 12'hfff;
rom[96883] = 12'hfff;
rom[96884] = 12'hfff;
rom[96885] = 12'hfff;
rom[96886] = 12'hfff;
rom[96887] = 12'hfff;
rom[96888] = 12'hfff;
rom[96889] = 12'hfff;
rom[96890] = 12'hfff;
rom[96891] = 12'hfff;
rom[96892] = 12'hfff;
rom[96893] = 12'hfff;
rom[96894] = 12'hfff;
rom[96895] = 12'hfff;
rom[96896] = 12'hfff;
rom[96897] = 12'hfff;
rom[96898] = 12'hfff;
rom[96899] = 12'hfff;
rom[96900] = 12'hfff;
rom[96901] = 12'hfff;
rom[96902] = 12'hfff;
rom[96903] = 12'hfff;
rom[96904] = 12'hfff;
rom[96905] = 12'hfff;
rom[96906] = 12'hfff;
rom[96907] = 12'hfff;
rom[96908] = 12'hfff;
rom[96909] = 12'hfff;
rom[96910] = 12'hfff;
rom[96911] = 12'hfff;
rom[96912] = 12'hfff;
rom[96913] = 12'hfff;
rom[96914] = 12'hfff;
rom[96915] = 12'hfff;
rom[96916] = 12'hfff;
rom[96917] = 12'hfff;
rom[96918] = 12'hfff;
rom[96919] = 12'hfff;
rom[96920] = 12'hfff;
rom[96921] = 12'hfff;
rom[96922] = 12'hfff;
rom[96923] = 12'hfff;
rom[96924] = 12'hfff;
rom[96925] = 12'hfff;
rom[96926] = 12'hfff;
rom[96927] = 12'hfff;
rom[96928] = 12'hfff;
rom[96929] = 12'hfff;
rom[96930] = 12'hfff;
rom[96931] = 12'hfff;
rom[96932] = 12'hfff;
rom[96933] = 12'hfff;
rom[96934] = 12'hfff;
rom[96935] = 12'hfff;
rom[96936] = 12'hfff;
rom[96937] = 12'hfff;
rom[96938] = 12'hfff;
rom[96939] = 12'hfff;
rom[96940] = 12'hfff;
rom[96941] = 12'hfff;
rom[96942] = 12'hfff;
rom[96943] = 12'hfff;
rom[96944] = 12'heee;
rom[96945] = 12'heee;
rom[96946] = 12'heee;
rom[96947] = 12'heee;
rom[96948] = 12'heee;
rom[96949] = 12'hddd;
rom[96950] = 12'hddd;
rom[96951] = 12'hddd;
rom[96952] = 12'hddd;
rom[96953] = 12'hddd;
rom[96954] = 12'hddd;
rom[96955] = 12'hddd;
rom[96956] = 12'hccc;
rom[96957] = 12'hccc;
rom[96958] = 12'hccc;
rom[96959] = 12'hccc;
rom[96960] = 12'hccc;
rom[96961] = 12'hccc;
rom[96962] = 12'hccc;
rom[96963] = 12'hccc;
rom[96964] = 12'hccc;
rom[96965] = 12'hccc;
rom[96966] = 12'hccc;
rom[96967] = 12'hccc;
rom[96968] = 12'hccc;
rom[96969] = 12'hccc;
rom[96970] = 12'hbbb;
rom[96971] = 12'hbbb;
rom[96972] = 12'hbbb;
rom[96973] = 12'hbbb;
rom[96974] = 12'haaa;
rom[96975] = 12'haaa;
rom[96976] = 12'haaa;
rom[96977] = 12'haaa;
rom[96978] = 12'h999;
rom[96979] = 12'h999;
rom[96980] = 12'h999;
rom[96981] = 12'h999;
rom[96982] = 12'h999;
rom[96983] = 12'h999;
rom[96984] = 12'h999;
rom[96985] = 12'h999;
rom[96986] = 12'h999;
rom[96987] = 12'h999;
rom[96988] = 12'h999;
rom[96989] = 12'h999;
rom[96990] = 12'h999;
rom[96991] = 12'h999;
rom[96992] = 12'h999;
rom[96993] = 12'h999;
rom[96994] = 12'h999;
rom[96995] = 12'h999;
rom[96996] = 12'h999;
rom[96997] = 12'h999;
rom[96998] = 12'h999;
rom[96999] = 12'h999;
rom[97000] = 12'h999;
rom[97001] = 12'h999;
rom[97002] = 12'h999;
rom[97003] = 12'h999;
rom[97004] = 12'h999;
rom[97005] = 12'haaa;
rom[97006] = 12'haaa;
rom[97007] = 12'haaa;
rom[97008] = 12'haaa;
rom[97009] = 12'haaa;
rom[97010] = 12'haaa;
rom[97011] = 12'haaa;
rom[97012] = 12'haaa;
rom[97013] = 12'haaa;
rom[97014] = 12'haaa;
rom[97015] = 12'haaa;
rom[97016] = 12'h999;
rom[97017] = 12'h999;
rom[97018] = 12'h999;
rom[97019] = 12'h888;
rom[97020] = 12'h888;
rom[97021] = 12'h888;
rom[97022] = 12'h888;
rom[97023] = 12'h888;
rom[97024] = 12'h888;
rom[97025] = 12'h888;
rom[97026] = 12'h888;
rom[97027] = 12'h888;
rom[97028] = 12'h888;
rom[97029] = 12'h888;
rom[97030] = 12'h888;
rom[97031] = 12'h888;
rom[97032] = 12'h888;
rom[97033] = 12'h999;
rom[97034] = 12'h999;
rom[97035] = 12'h999;
rom[97036] = 12'h999;
rom[97037] = 12'h999;
rom[97038] = 12'h999;
rom[97039] = 12'h999;
rom[97040] = 12'h999;
rom[97041] = 12'h999;
rom[97042] = 12'h999;
rom[97043] = 12'h888;
rom[97044] = 12'h888;
rom[97045] = 12'h777;
rom[97046] = 12'h777;
rom[97047] = 12'h777;
rom[97048] = 12'h777;
rom[97049] = 12'h777;
rom[97050] = 12'h777;
rom[97051] = 12'h777;
rom[97052] = 12'h888;
rom[97053] = 12'h888;
rom[97054] = 12'h777;
rom[97055] = 12'h777;
rom[97056] = 12'h888;
rom[97057] = 12'h888;
rom[97058] = 12'h888;
rom[97059] = 12'h888;
rom[97060] = 12'h999;
rom[97061] = 12'h999;
rom[97062] = 12'h999;
rom[97063] = 12'h999;
rom[97064] = 12'h999;
rom[97065] = 12'h999;
rom[97066] = 12'h999;
rom[97067] = 12'h999;
rom[97068] = 12'h999;
rom[97069] = 12'h888;
rom[97070] = 12'h888;
rom[97071] = 12'h888;
rom[97072] = 12'h888;
rom[97073] = 12'h888;
rom[97074] = 12'h888;
rom[97075] = 12'h888;
rom[97076] = 12'h888;
rom[97077] = 12'h888;
rom[97078] = 12'h888;
rom[97079] = 12'h888;
rom[97080] = 12'h888;
rom[97081] = 12'h777;
rom[97082] = 12'h888;
rom[97083] = 12'h888;
rom[97084] = 12'h999;
rom[97085] = 12'haaa;
rom[97086] = 12'hbbb;
rom[97087] = 12'hccc;
rom[97088] = 12'heee;
rom[97089] = 12'heee;
rom[97090] = 12'hfff;
rom[97091] = 12'heee;
rom[97092] = 12'hddd;
rom[97093] = 12'hccc;
rom[97094] = 12'hbbb;
rom[97095] = 12'hccc;
rom[97096] = 12'hccc;
rom[97097] = 12'hddd;
rom[97098] = 12'heee;
rom[97099] = 12'heee;
rom[97100] = 12'hccc;
rom[97101] = 12'haaa;
rom[97102] = 12'h888;
rom[97103] = 12'h666;
rom[97104] = 12'h555;
rom[97105] = 12'h666;
rom[97106] = 12'h666;
rom[97107] = 12'h555;
rom[97108] = 12'h555;
rom[97109] = 12'h666;
rom[97110] = 12'h666;
rom[97111] = 12'h555;
rom[97112] = 12'h666;
rom[97113] = 12'h777;
rom[97114] = 12'h999;
rom[97115] = 12'h999;
rom[97116] = 12'haaa;
rom[97117] = 12'hbbb;
rom[97118] = 12'hddd;
rom[97119] = 12'heee;
rom[97120] = 12'hfff;
rom[97121] = 12'hfff;
rom[97122] = 12'hfff;
rom[97123] = 12'hddd;
rom[97124] = 12'hbbb;
rom[97125] = 12'h999;
rom[97126] = 12'h777;
rom[97127] = 12'h555;
rom[97128] = 12'h444;
rom[97129] = 12'h444;
rom[97130] = 12'h333;
rom[97131] = 12'h333;
rom[97132] = 12'h333;
rom[97133] = 12'h222;
rom[97134] = 12'h222;
rom[97135] = 12'h222;
rom[97136] = 12'h222;
rom[97137] = 12'h222;
rom[97138] = 12'h111;
rom[97139] = 12'h111;
rom[97140] = 12'h111;
rom[97141] = 12'h111;
rom[97142] = 12'h222;
rom[97143] = 12'h222;
rom[97144] = 12'h222;
rom[97145] = 12'h222;
rom[97146] = 12'h111;
rom[97147] = 12'h111;
rom[97148] = 12'h  0;
rom[97149] = 12'h  0;
rom[97150] = 12'h111;
rom[97151] = 12'h111;
rom[97152] = 12'h111;
rom[97153] = 12'h111;
rom[97154] = 12'h111;
rom[97155] = 12'h111;
rom[97156] = 12'h111;
rom[97157] = 12'h111;
rom[97158] = 12'h111;
rom[97159] = 12'h111;
rom[97160] = 12'h111;
rom[97161] = 12'h111;
rom[97162] = 12'h111;
rom[97163] = 12'h111;
rom[97164] = 12'h111;
rom[97165] = 12'h111;
rom[97166] = 12'h111;
rom[97167] = 12'h111;
rom[97168] = 12'h111;
rom[97169] = 12'h222;
rom[97170] = 12'h222;
rom[97171] = 12'h222;
rom[97172] = 12'h222;
rom[97173] = 12'h222;
rom[97174] = 12'h222;
rom[97175] = 12'h333;
rom[97176] = 12'h222;
rom[97177] = 12'h333;
rom[97178] = 12'h444;
rom[97179] = 12'h555;
rom[97180] = 12'h666;
rom[97181] = 12'h666;
rom[97182] = 12'h666;
rom[97183] = 12'h555;
rom[97184] = 12'h555;
rom[97185] = 12'h555;
rom[97186] = 12'h666;
rom[97187] = 12'h777;
rom[97188] = 12'h777;
rom[97189] = 12'h777;
rom[97190] = 12'h666;
rom[97191] = 12'h666;
rom[97192] = 12'h555;
rom[97193] = 12'h555;
rom[97194] = 12'h444;
rom[97195] = 12'h333;
rom[97196] = 12'h222;
rom[97197] = 12'h222;
rom[97198] = 12'h222;
rom[97199] = 12'h222;
rom[97200] = 12'hfff;
rom[97201] = 12'hfff;
rom[97202] = 12'hfff;
rom[97203] = 12'hfff;
rom[97204] = 12'hfff;
rom[97205] = 12'hfff;
rom[97206] = 12'hfff;
rom[97207] = 12'hfff;
rom[97208] = 12'hfff;
rom[97209] = 12'hfff;
rom[97210] = 12'hfff;
rom[97211] = 12'hfff;
rom[97212] = 12'hfff;
rom[97213] = 12'hfff;
rom[97214] = 12'hfff;
rom[97215] = 12'hfff;
rom[97216] = 12'hfff;
rom[97217] = 12'hfff;
rom[97218] = 12'hfff;
rom[97219] = 12'hfff;
rom[97220] = 12'hfff;
rom[97221] = 12'hfff;
rom[97222] = 12'hfff;
rom[97223] = 12'hfff;
rom[97224] = 12'hfff;
rom[97225] = 12'hfff;
rom[97226] = 12'hfff;
rom[97227] = 12'hfff;
rom[97228] = 12'hfff;
rom[97229] = 12'hfff;
rom[97230] = 12'hfff;
rom[97231] = 12'hfff;
rom[97232] = 12'hfff;
rom[97233] = 12'hfff;
rom[97234] = 12'hfff;
rom[97235] = 12'hfff;
rom[97236] = 12'hfff;
rom[97237] = 12'hfff;
rom[97238] = 12'hfff;
rom[97239] = 12'hfff;
rom[97240] = 12'hfff;
rom[97241] = 12'hfff;
rom[97242] = 12'hfff;
rom[97243] = 12'hfff;
rom[97244] = 12'hfff;
rom[97245] = 12'hfff;
rom[97246] = 12'hfff;
rom[97247] = 12'hfff;
rom[97248] = 12'hfff;
rom[97249] = 12'hfff;
rom[97250] = 12'hfff;
rom[97251] = 12'hfff;
rom[97252] = 12'hfff;
rom[97253] = 12'hfff;
rom[97254] = 12'hfff;
rom[97255] = 12'hfff;
rom[97256] = 12'hfff;
rom[97257] = 12'hfff;
rom[97258] = 12'hfff;
rom[97259] = 12'hfff;
rom[97260] = 12'hfff;
rom[97261] = 12'hfff;
rom[97262] = 12'hfff;
rom[97263] = 12'hfff;
rom[97264] = 12'hfff;
rom[97265] = 12'hfff;
rom[97266] = 12'hfff;
rom[97267] = 12'hfff;
rom[97268] = 12'hfff;
rom[97269] = 12'hfff;
rom[97270] = 12'hfff;
rom[97271] = 12'hfff;
rom[97272] = 12'hfff;
rom[97273] = 12'hfff;
rom[97274] = 12'hfff;
rom[97275] = 12'hfff;
rom[97276] = 12'hfff;
rom[97277] = 12'hfff;
rom[97278] = 12'hfff;
rom[97279] = 12'hfff;
rom[97280] = 12'hfff;
rom[97281] = 12'hfff;
rom[97282] = 12'hfff;
rom[97283] = 12'hfff;
rom[97284] = 12'hfff;
rom[97285] = 12'hfff;
rom[97286] = 12'hfff;
rom[97287] = 12'hfff;
rom[97288] = 12'hfff;
rom[97289] = 12'hfff;
rom[97290] = 12'hfff;
rom[97291] = 12'hfff;
rom[97292] = 12'hfff;
rom[97293] = 12'hfff;
rom[97294] = 12'hfff;
rom[97295] = 12'hfff;
rom[97296] = 12'hfff;
rom[97297] = 12'hfff;
rom[97298] = 12'hfff;
rom[97299] = 12'hfff;
rom[97300] = 12'hfff;
rom[97301] = 12'hfff;
rom[97302] = 12'hfff;
rom[97303] = 12'hfff;
rom[97304] = 12'hfff;
rom[97305] = 12'hfff;
rom[97306] = 12'hfff;
rom[97307] = 12'hfff;
rom[97308] = 12'hfff;
rom[97309] = 12'hfff;
rom[97310] = 12'hfff;
rom[97311] = 12'hfff;
rom[97312] = 12'hfff;
rom[97313] = 12'hfff;
rom[97314] = 12'hfff;
rom[97315] = 12'hfff;
rom[97316] = 12'hfff;
rom[97317] = 12'hfff;
rom[97318] = 12'hfff;
rom[97319] = 12'hfff;
rom[97320] = 12'hfff;
rom[97321] = 12'hfff;
rom[97322] = 12'hfff;
rom[97323] = 12'hfff;
rom[97324] = 12'hfff;
rom[97325] = 12'hfff;
rom[97326] = 12'hfff;
rom[97327] = 12'hfff;
rom[97328] = 12'hfff;
rom[97329] = 12'hfff;
rom[97330] = 12'hfff;
rom[97331] = 12'hfff;
rom[97332] = 12'hfff;
rom[97333] = 12'hfff;
rom[97334] = 12'hfff;
rom[97335] = 12'hfff;
rom[97336] = 12'hfff;
rom[97337] = 12'hfff;
rom[97338] = 12'hfff;
rom[97339] = 12'hfff;
rom[97340] = 12'hfff;
rom[97341] = 12'hfff;
rom[97342] = 12'hfff;
rom[97343] = 12'hfff;
rom[97344] = 12'hfff;
rom[97345] = 12'heee;
rom[97346] = 12'heee;
rom[97347] = 12'heee;
rom[97348] = 12'heee;
rom[97349] = 12'heee;
rom[97350] = 12'hddd;
rom[97351] = 12'hddd;
rom[97352] = 12'hddd;
rom[97353] = 12'hddd;
rom[97354] = 12'hddd;
rom[97355] = 12'hddd;
rom[97356] = 12'hddd;
rom[97357] = 12'hccc;
rom[97358] = 12'hccc;
rom[97359] = 12'hccc;
rom[97360] = 12'hccc;
rom[97361] = 12'hccc;
rom[97362] = 12'hccc;
rom[97363] = 12'hccc;
rom[97364] = 12'hccc;
rom[97365] = 12'hccc;
rom[97366] = 12'hccc;
rom[97367] = 12'hccc;
rom[97368] = 12'hccc;
rom[97369] = 12'hccc;
rom[97370] = 12'hccc;
rom[97371] = 12'hccc;
rom[97372] = 12'hbbb;
rom[97373] = 12'hbbb;
rom[97374] = 12'hbbb;
rom[97375] = 12'hbbb;
rom[97376] = 12'haaa;
rom[97377] = 12'haaa;
rom[97378] = 12'haaa;
rom[97379] = 12'haaa;
rom[97380] = 12'h999;
rom[97381] = 12'haaa;
rom[97382] = 12'haaa;
rom[97383] = 12'haaa;
rom[97384] = 12'haaa;
rom[97385] = 12'haaa;
rom[97386] = 12'h999;
rom[97387] = 12'h999;
rom[97388] = 12'h999;
rom[97389] = 12'h999;
rom[97390] = 12'h999;
rom[97391] = 12'h999;
rom[97392] = 12'h999;
rom[97393] = 12'h999;
rom[97394] = 12'h999;
rom[97395] = 12'h999;
rom[97396] = 12'h999;
rom[97397] = 12'h999;
rom[97398] = 12'h999;
rom[97399] = 12'h999;
rom[97400] = 12'h999;
rom[97401] = 12'h999;
rom[97402] = 12'h999;
rom[97403] = 12'h999;
rom[97404] = 12'haaa;
rom[97405] = 12'haaa;
rom[97406] = 12'haaa;
rom[97407] = 12'haaa;
rom[97408] = 12'haaa;
rom[97409] = 12'haaa;
rom[97410] = 12'haaa;
rom[97411] = 12'haaa;
rom[97412] = 12'haaa;
rom[97413] = 12'haaa;
rom[97414] = 12'haaa;
rom[97415] = 12'haaa;
rom[97416] = 12'haaa;
rom[97417] = 12'haaa;
rom[97418] = 12'h999;
rom[97419] = 12'h999;
rom[97420] = 12'h999;
rom[97421] = 12'h888;
rom[97422] = 12'h888;
rom[97423] = 12'h888;
rom[97424] = 12'h888;
rom[97425] = 12'h888;
rom[97426] = 12'h888;
rom[97427] = 12'h888;
rom[97428] = 12'h888;
rom[97429] = 12'h888;
rom[97430] = 12'h888;
rom[97431] = 12'h888;
rom[97432] = 12'h999;
rom[97433] = 12'h999;
rom[97434] = 12'h999;
rom[97435] = 12'h999;
rom[97436] = 12'h999;
rom[97437] = 12'h999;
rom[97438] = 12'h999;
rom[97439] = 12'h999;
rom[97440] = 12'h999;
rom[97441] = 12'h999;
rom[97442] = 12'h999;
rom[97443] = 12'h999;
rom[97444] = 12'h888;
rom[97445] = 12'h888;
rom[97446] = 12'h888;
rom[97447] = 12'h888;
rom[97448] = 12'h777;
rom[97449] = 12'h777;
rom[97450] = 12'h777;
rom[97451] = 12'h888;
rom[97452] = 12'h888;
rom[97453] = 12'h888;
rom[97454] = 12'h888;
rom[97455] = 12'h888;
rom[97456] = 12'h888;
rom[97457] = 12'h888;
rom[97458] = 12'h999;
rom[97459] = 12'h999;
rom[97460] = 12'h999;
rom[97461] = 12'h999;
rom[97462] = 12'h999;
rom[97463] = 12'h999;
rom[97464] = 12'h999;
rom[97465] = 12'h999;
rom[97466] = 12'h999;
rom[97467] = 12'h999;
rom[97468] = 12'h888;
rom[97469] = 12'h888;
rom[97470] = 12'h888;
rom[97471] = 12'h888;
rom[97472] = 12'h888;
rom[97473] = 12'h888;
rom[97474] = 12'h888;
rom[97475] = 12'h888;
rom[97476] = 12'h888;
rom[97477] = 12'h888;
rom[97478] = 12'h888;
rom[97479] = 12'h888;
rom[97480] = 12'h888;
rom[97481] = 12'h888;
rom[97482] = 12'h888;
rom[97483] = 12'h999;
rom[97484] = 12'haaa;
rom[97485] = 12'hbbb;
rom[97486] = 12'hddd;
rom[97487] = 12'heee;
rom[97488] = 12'hfff;
rom[97489] = 12'hfff;
rom[97490] = 12'heee;
rom[97491] = 12'hddd;
rom[97492] = 12'hccc;
rom[97493] = 12'haaa;
rom[97494] = 12'haaa;
rom[97495] = 12'haaa;
rom[97496] = 12'hbbb;
rom[97497] = 12'hccc;
rom[97498] = 12'hddd;
rom[97499] = 12'heee;
rom[97500] = 12'heee;
rom[97501] = 12'hddd;
rom[97502] = 12'haaa;
rom[97503] = 12'h888;
rom[97504] = 12'h666;
rom[97505] = 12'h666;
rom[97506] = 12'h555;
rom[97507] = 12'h555;
rom[97508] = 12'h666;
rom[97509] = 12'h666;
rom[97510] = 12'h555;
rom[97511] = 12'h555;
rom[97512] = 12'h555;
rom[97513] = 12'h666;
rom[97514] = 12'h777;
rom[97515] = 12'h888;
rom[97516] = 12'h888;
rom[97517] = 12'h999;
rom[97518] = 12'haaa;
rom[97519] = 12'hbbb;
rom[97520] = 12'hccc;
rom[97521] = 12'heee;
rom[97522] = 12'hfff;
rom[97523] = 12'hfff;
rom[97524] = 12'heee;
rom[97525] = 12'hccc;
rom[97526] = 12'haaa;
rom[97527] = 12'h888;
rom[97528] = 12'h666;
rom[97529] = 12'h555;
rom[97530] = 12'h444;
rom[97531] = 12'h333;
rom[97532] = 12'h333;
rom[97533] = 12'h333;
rom[97534] = 12'h222;
rom[97535] = 12'h222;
rom[97536] = 12'h222;
rom[97537] = 12'h222;
rom[97538] = 12'h111;
rom[97539] = 12'h111;
rom[97540] = 12'h  0;
rom[97541] = 12'h111;
rom[97542] = 12'h111;
rom[97543] = 12'h111;
rom[97544] = 12'h222;
rom[97545] = 12'h222;
rom[97546] = 12'h222;
rom[97547] = 12'h111;
rom[97548] = 12'h111;
rom[97549] = 12'h111;
rom[97550] = 12'h111;
rom[97551] = 12'h111;
rom[97552] = 12'h111;
rom[97553] = 12'h111;
rom[97554] = 12'h111;
rom[97555] = 12'h111;
rom[97556] = 12'h111;
rom[97557] = 12'h111;
rom[97558] = 12'h111;
rom[97559] = 12'h111;
rom[97560] = 12'h111;
rom[97561] = 12'h111;
rom[97562] = 12'h111;
rom[97563] = 12'h111;
rom[97564] = 12'h111;
rom[97565] = 12'h111;
rom[97566] = 12'h111;
rom[97567] = 12'h111;
rom[97568] = 12'h111;
rom[97569] = 12'h111;
rom[97570] = 12'h111;
rom[97571] = 12'h111;
rom[97572] = 12'h111;
rom[97573] = 12'h111;
rom[97574] = 12'h222;
rom[97575] = 12'h222;
rom[97576] = 12'h222;
rom[97577] = 12'h222;
rom[97578] = 12'h333;
rom[97579] = 12'h333;
rom[97580] = 12'h555;
rom[97581] = 12'h555;
rom[97582] = 12'h666;
rom[97583] = 12'h666;
rom[97584] = 12'h444;
rom[97585] = 12'h444;
rom[97586] = 12'h555;
rom[97587] = 12'h555;
rom[97588] = 12'h555;
rom[97589] = 12'h666;
rom[97590] = 12'h666;
rom[97591] = 12'h666;
rom[97592] = 12'h666;
rom[97593] = 12'h666;
rom[97594] = 12'h666;
rom[97595] = 12'h555;
rom[97596] = 12'h555;
rom[97597] = 12'h444;
rom[97598] = 12'h333;
rom[97599] = 12'h333;
rom[97600] = 12'hfff;
rom[97601] = 12'hfff;
rom[97602] = 12'hfff;
rom[97603] = 12'hfff;
rom[97604] = 12'hfff;
rom[97605] = 12'hfff;
rom[97606] = 12'hfff;
rom[97607] = 12'hfff;
rom[97608] = 12'hfff;
rom[97609] = 12'hfff;
rom[97610] = 12'hfff;
rom[97611] = 12'hfff;
rom[97612] = 12'hfff;
rom[97613] = 12'hfff;
rom[97614] = 12'hfff;
rom[97615] = 12'hfff;
rom[97616] = 12'hfff;
rom[97617] = 12'hfff;
rom[97618] = 12'hfff;
rom[97619] = 12'hfff;
rom[97620] = 12'hfff;
rom[97621] = 12'hfff;
rom[97622] = 12'hfff;
rom[97623] = 12'hfff;
rom[97624] = 12'hfff;
rom[97625] = 12'hfff;
rom[97626] = 12'hfff;
rom[97627] = 12'hfff;
rom[97628] = 12'hfff;
rom[97629] = 12'hfff;
rom[97630] = 12'hfff;
rom[97631] = 12'hfff;
rom[97632] = 12'hfff;
rom[97633] = 12'hfff;
rom[97634] = 12'hfff;
rom[97635] = 12'hfff;
rom[97636] = 12'hfff;
rom[97637] = 12'hfff;
rom[97638] = 12'hfff;
rom[97639] = 12'hfff;
rom[97640] = 12'hfff;
rom[97641] = 12'hfff;
rom[97642] = 12'hfff;
rom[97643] = 12'hfff;
rom[97644] = 12'hfff;
rom[97645] = 12'hfff;
rom[97646] = 12'hfff;
rom[97647] = 12'hfff;
rom[97648] = 12'hfff;
rom[97649] = 12'hfff;
rom[97650] = 12'hfff;
rom[97651] = 12'hfff;
rom[97652] = 12'hfff;
rom[97653] = 12'hfff;
rom[97654] = 12'hfff;
rom[97655] = 12'hfff;
rom[97656] = 12'hfff;
rom[97657] = 12'hfff;
rom[97658] = 12'hfff;
rom[97659] = 12'hfff;
rom[97660] = 12'hfff;
rom[97661] = 12'hfff;
rom[97662] = 12'hfff;
rom[97663] = 12'hfff;
rom[97664] = 12'hfff;
rom[97665] = 12'hfff;
rom[97666] = 12'hfff;
rom[97667] = 12'hfff;
rom[97668] = 12'hfff;
rom[97669] = 12'hfff;
rom[97670] = 12'hfff;
rom[97671] = 12'hfff;
rom[97672] = 12'hfff;
rom[97673] = 12'hfff;
rom[97674] = 12'hfff;
rom[97675] = 12'hfff;
rom[97676] = 12'hfff;
rom[97677] = 12'hfff;
rom[97678] = 12'hfff;
rom[97679] = 12'hfff;
rom[97680] = 12'hfff;
rom[97681] = 12'hfff;
rom[97682] = 12'hfff;
rom[97683] = 12'hfff;
rom[97684] = 12'hfff;
rom[97685] = 12'hfff;
rom[97686] = 12'hfff;
rom[97687] = 12'hfff;
rom[97688] = 12'hfff;
rom[97689] = 12'hfff;
rom[97690] = 12'hfff;
rom[97691] = 12'hfff;
rom[97692] = 12'hfff;
rom[97693] = 12'hfff;
rom[97694] = 12'hfff;
rom[97695] = 12'hfff;
rom[97696] = 12'hfff;
rom[97697] = 12'hfff;
rom[97698] = 12'hfff;
rom[97699] = 12'hfff;
rom[97700] = 12'hfff;
rom[97701] = 12'hfff;
rom[97702] = 12'hfff;
rom[97703] = 12'hfff;
rom[97704] = 12'hfff;
rom[97705] = 12'hfff;
rom[97706] = 12'hfff;
rom[97707] = 12'hfff;
rom[97708] = 12'hfff;
rom[97709] = 12'hfff;
rom[97710] = 12'hfff;
rom[97711] = 12'hfff;
rom[97712] = 12'hfff;
rom[97713] = 12'hfff;
rom[97714] = 12'hfff;
rom[97715] = 12'hfff;
rom[97716] = 12'hfff;
rom[97717] = 12'hfff;
rom[97718] = 12'hfff;
rom[97719] = 12'hfff;
rom[97720] = 12'hfff;
rom[97721] = 12'hfff;
rom[97722] = 12'hfff;
rom[97723] = 12'hfff;
rom[97724] = 12'hfff;
rom[97725] = 12'hfff;
rom[97726] = 12'hfff;
rom[97727] = 12'hfff;
rom[97728] = 12'hfff;
rom[97729] = 12'hfff;
rom[97730] = 12'hfff;
rom[97731] = 12'hfff;
rom[97732] = 12'hfff;
rom[97733] = 12'hfff;
rom[97734] = 12'hfff;
rom[97735] = 12'hfff;
rom[97736] = 12'hfff;
rom[97737] = 12'hfff;
rom[97738] = 12'hfff;
rom[97739] = 12'hfff;
rom[97740] = 12'hfff;
rom[97741] = 12'hfff;
rom[97742] = 12'hfff;
rom[97743] = 12'hfff;
rom[97744] = 12'hfff;
rom[97745] = 12'hfff;
rom[97746] = 12'heee;
rom[97747] = 12'heee;
rom[97748] = 12'heee;
rom[97749] = 12'heee;
rom[97750] = 12'heee;
rom[97751] = 12'hddd;
rom[97752] = 12'hddd;
rom[97753] = 12'hddd;
rom[97754] = 12'hddd;
rom[97755] = 12'hddd;
rom[97756] = 12'hddd;
rom[97757] = 12'hccc;
rom[97758] = 12'hccc;
rom[97759] = 12'hccc;
rom[97760] = 12'hccc;
rom[97761] = 12'hccc;
rom[97762] = 12'hccc;
rom[97763] = 12'hccc;
rom[97764] = 12'hccc;
rom[97765] = 12'hccc;
rom[97766] = 12'hccc;
rom[97767] = 12'hccc;
rom[97768] = 12'hccc;
rom[97769] = 12'hccc;
rom[97770] = 12'hccc;
rom[97771] = 12'hccc;
rom[97772] = 12'hccc;
rom[97773] = 12'hccc;
rom[97774] = 12'hbbb;
rom[97775] = 12'hbbb;
rom[97776] = 12'hbbb;
rom[97777] = 12'haaa;
rom[97778] = 12'haaa;
rom[97779] = 12'haaa;
rom[97780] = 12'haaa;
rom[97781] = 12'haaa;
rom[97782] = 12'haaa;
rom[97783] = 12'haaa;
rom[97784] = 12'haaa;
rom[97785] = 12'haaa;
rom[97786] = 12'h999;
rom[97787] = 12'h999;
rom[97788] = 12'h999;
rom[97789] = 12'h999;
rom[97790] = 12'h999;
rom[97791] = 12'h999;
rom[97792] = 12'h999;
rom[97793] = 12'h999;
rom[97794] = 12'h999;
rom[97795] = 12'h999;
rom[97796] = 12'h999;
rom[97797] = 12'h999;
rom[97798] = 12'h999;
rom[97799] = 12'h999;
rom[97800] = 12'h999;
rom[97801] = 12'h999;
rom[97802] = 12'h999;
rom[97803] = 12'haaa;
rom[97804] = 12'haaa;
rom[97805] = 12'haaa;
rom[97806] = 12'haaa;
rom[97807] = 12'haaa;
rom[97808] = 12'haaa;
rom[97809] = 12'haaa;
rom[97810] = 12'haaa;
rom[97811] = 12'haaa;
rom[97812] = 12'haaa;
rom[97813] = 12'haaa;
rom[97814] = 12'haaa;
rom[97815] = 12'haaa;
rom[97816] = 12'haaa;
rom[97817] = 12'haaa;
rom[97818] = 12'haaa;
rom[97819] = 12'haaa;
rom[97820] = 12'h999;
rom[97821] = 12'h999;
rom[97822] = 12'h888;
rom[97823] = 12'h888;
rom[97824] = 12'h888;
rom[97825] = 12'h888;
rom[97826] = 12'h888;
rom[97827] = 12'h888;
rom[97828] = 12'h888;
rom[97829] = 12'h888;
rom[97830] = 12'h888;
rom[97831] = 12'h999;
rom[97832] = 12'h999;
rom[97833] = 12'h999;
rom[97834] = 12'h999;
rom[97835] = 12'h999;
rom[97836] = 12'haaa;
rom[97837] = 12'haaa;
rom[97838] = 12'haaa;
rom[97839] = 12'haaa;
rom[97840] = 12'haaa;
rom[97841] = 12'h999;
rom[97842] = 12'h999;
rom[97843] = 12'h999;
rom[97844] = 12'h999;
rom[97845] = 12'h888;
rom[97846] = 12'h888;
rom[97847] = 12'h888;
rom[97848] = 12'h888;
rom[97849] = 12'h777;
rom[97850] = 12'h777;
rom[97851] = 12'h888;
rom[97852] = 12'h888;
rom[97853] = 12'h888;
rom[97854] = 12'h888;
rom[97855] = 12'h999;
rom[97856] = 12'h999;
rom[97857] = 12'h999;
rom[97858] = 12'h999;
rom[97859] = 12'haaa;
rom[97860] = 12'haaa;
rom[97861] = 12'haaa;
rom[97862] = 12'haaa;
rom[97863] = 12'h999;
rom[97864] = 12'h999;
rom[97865] = 12'h999;
rom[97866] = 12'h888;
rom[97867] = 12'h888;
rom[97868] = 12'h888;
rom[97869] = 12'h888;
rom[97870] = 12'h777;
rom[97871] = 12'h777;
rom[97872] = 12'h888;
rom[97873] = 12'h888;
rom[97874] = 12'h888;
rom[97875] = 12'h888;
rom[97876] = 12'h888;
rom[97877] = 12'h888;
rom[97878] = 12'h888;
rom[97879] = 12'h888;
rom[97880] = 12'h999;
rom[97881] = 12'h999;
rom[97882] = 12'h999;
rom[97883] = 12'haaa;
rom[97884] = 12'hbbb;
rom[97885] = 12'hddd;
rom[97886] = 12'heee;
rom[97887] = 12'hfff;
rom[97888] = 12'hfff;
rom[97889] = 12'heee;
rom[97890] = 12'hddd;
rom[97891] = 12'hccc;
rom[97892] = 12'haaa;
rom[97893] = 12'h999;
rom[97894] = 12'h888;
rom[97895] = 12'h888;
rom[97896] = 12'h999;
rom[97897] = 12'haaa;
rom[97898] = 12'hbbb;
rom[97899] = 12'hddd;
rom[97900] = 12'heee;
rom[97901] = 12'heee;
rom[97902] = 12'hddd;
rom[97903] = 12'hbbb;
rom[97904] = 12'h888;
rom[97905] = 12'h666;
rom[97906] = 12'h555;
rom[97907] = 12'h555;
rom[97908] = 12'h555;
rom[97909] = 12'h555;
rom[97910] = 12'h555;
rom[97911] = 12'h555;
rom[97912] = 12'h666;
rom[97913] = 12'h666;
rom[97914] = 12'h666;
rom[97915] = 12'h777;
rom[97916] = 12'h888;
rom[97917] = 12'h888;
rom[97918] = 12'h777;
rom[97919] = 12'h777;
rom[97920] = 12'h999;
rom[97921] = 12'hbbb;
rom[97922] = 12'hddd;
rom[97923] = 12'hfff;
rom[97924] = 12'hfff;
rom[97925] = 12'hfff;
rom[97926] = 12'heee;
rom[97927] = 12'hccc;
rom[97928] = 12'h999;
rom[97929] = 12'h777;
rom[97930] = 12'h555;
rom[97931] = 12'h444;
rom[97932] = 12'h444;
rom[97933] = 12'h333;
rom[97934] = 12'h333;
rom[97935] = 12'h333;
rom[97936] = 12'h222;
rom[97937] = 12'h222;
rom[97938] = 12'h222;
rom[97939] = 12'h111;
rom[97940] = 12'h111;
rom[97941] = 12'h  0;
rom[97942] = 12'h111;
rom[97943] = 12'h111;
rom[97944] = 12'h111;
rom[97945] = 12'h222;
rom[97946] = 12'h222;
rom[97947] = 12'h222;
rom[97948] = 12'h111;
rom[97949] = 12'h111;
rom[97950] = 12'h111;
rom[97951] = 12'h111;
rom[97952] = 12'h111;
rom[97953] = 12'h111;
rom[97954] = 12'h111;
rom[97955] = 12'h111;
rom[97956] = 12'h111;
rom[97957] = 12'h111;
rom[97958] = 12'h111;
rom[97959] = 12'h111;
rom[97960] = 12'h111;
rom[97961] = 12'h111;
rom[97962] = 12'h111;
rom[97963] = 12'h111;
rom[97964] = 12'h111;
rom[97965] = 12'h111;
rom[97966] = 12'h111;
rom[97967] = 12'h111;
rom[97968] = 12'h111;
rom[97969] = 12'h111;
rom[97970] = 12'h111;
rom[97971] = 12'h111;
rom[97972] = 12'h111;
rom[97973] = 12'h111;
rom[97974] = 12'h111;
rom[97975] = 12'h111;
rom[97976] = 12'h222;
rom[97977] = 12'h222;
rom[97978] = 12'h222;
rom[97979] = 12'h333;
rom[97980] = 12'h333;
rom[97981] = 12'h444;
rom[97982] = 12'h555;
rom[97983] = 12'h555;
rom[97984] = 12'h555;
rom[97985] = 12'h444;
rom[97986] = 12'h444;
rom[97987] = 12'h333;
rom[97988] = 12'h444;
rom[97989] = 12'h444;
rom[97990] = 12'h555;
rom[97991] = 12'h555;
rom[97992] = 12'h666;
rom[97993] = 12'h666;
rom[97994] = 12'h666;
rom[97995] = 12'h666;
rom[97996] = 12'h666;
rom[97997] = 12'h555;
rom[97998] = 12'h555;
rom[97999] = 12'h555;
rom[98000] = 12'hfff;
rom[98001] = 12'hfff;
rom[98002] = 12'hfff;
rom[98003] = 12'hfff;
rom[98004] = 12'hfff;
rom[98005] = 12'hfff;
rom[98006] = 12'hfff;
rom[98007] = 12'hfff;
rom[98008] = 12'hfff;
rom[98009] = 12'hfff;
rom[98010] = 12'hfff;
rom[98011] = 12'hfff;
rom[98012] = 12'hfff;
rom[98013] = 12'hfff;
rom[98014] = 12'hfff;
rom[98015] = 12'hfff;
rom[98016] = 12'hfff;
rom[98017] = 12'hfff;
rom[98018] = 12'hfff;
rom[98019] = 12'hfff;
rom[98020] = 12'hfff;
rom[98021] = 12'hfff;
rom[98022] = 12'hfff;
rom[98023] = 12'hfff;
rom[98024] = 12'hfff;
rom[98025] = 12'hfff;
rom[98026] = 12'hfff;
rom[98027] = 12'hfff;
rom[98028] = 12'hfff;
rom[98029] = 12'hfff;
rom[98030] = 12'hfff;
rom[98031] = 12'hfff;
rom[98032] = 12'hfff;
rom[98033] = 12'hfff;
rom[98034] = 12'hfff;
rom[98035] = 12'hfff;
rom[98036] = 12'hfff;
rom[98037] = 12'hfff;
rom[98038] = 12'hfff;
rom[98039] = 12'hfff;
rom[98040] = 12'hfff;
rom[98041] = 12'hfff;
rom[98042] = 12'hfff;
rom[98043] = 12'hfff;
rom[98044] = 12'hfff;
rom[98045] = 12'hfff;
rom[98046] = 12'hfff;
rom[98047] = 12'hfff;
rom[98048] = 12'hfff;
rom[98049] = 12'hfff;
rom[98050] = 12'hfff;
rom[98051] = 12'hfff;
rom[98052] = 12'hfff;
rom[98053] = 12'hfff;
rom[98054] = 12'hfff;
rom[98055] = 12'hfff;
rom[98056] = 12'hfff;
rom[98057] = 12'hfff;
rom[98058] = 12'hfff;
rom[98059] = 12'hfff;
rom[98060] = 12'hfff;
rom[98061] = 12'hfff;
rom[98062] = 12'hfff;
rom[98063] = 12'hfff;
rom[98064] = 12'hfff;
rom[98065] = 12'hfff;
rom[98066] = 12'hfff;
rom[98067] = 12'hfff;
rom[98068] = 12'hfff;
rom[98069] = 12'hfff;
rom[98070] = 12'hfff;
rom[98071] = 12'hfff;
rom[98072] = 12'hfff;
rom[98073] = 12'hfff;
rom[98074] = 12'hfff;
rom[98075] = 12'hfff;
rom[98076] = 12'hfff;
rom[98077] = 12'hfff;
rom[98078] = 12'hfff;
rom[98079] = 12'hfff;
rom[98080] = 12'hfff;
rom[98081] = 12'hfff;
rom[98082] = 12'hfff;
rom[98083] = 12'hfff;
rom[98084] = 12'hfff;
rom[98085] = 12'hfff;
rom[98086] = 12'hfff;
rom[98087] = 12'hfff;
rom[98088] = 12'hfff;
rom[98089] = 12'hfff;
rom[98090] = 12'hfff;
rom[98091] = 12'hfff;
rom[98092] = 12'hfff;
rom[98093] = 12'hfff;
rom[98094] = 12'hfff;
rom[98095] = 12'hfff;
rom[98096] = 12'hfff;
rom[98097] = 12'hfff;
rom[98098] = 12'hfff;
rom[98099] = 12'hfff;
rom[98100] = 12'hfff;
rom[98101] = 12'hfff;
rom[98102] = 12'hfff;
rom[98103] = 12'hfff;
rom[98104] = 12'hfff;
rom[98105] = 12'hfff;
rom[98106] = 12'hfff;
rom[98107] = 12'hfff;
rom[98108] = 12'hfff;
rom[98109] = 12'hfff;
rom[98110] = 12'hfff;
rom[98111] = 12'hfff;
rom[98112] = 12'hfff;
rom[98113] = 12'hfff;
rom[98114] = 12'hfff;
rom[98115] = 12'hfff;
rom[98116] = 12'hfff;
rom[98117] = 12'hfff;
rom[98118] = 12'hfff;
rom[98119] = 12'hfff;
rom[98120] = 12'hfff;
rom[98121] = 12'hfff;
rom[98122] = 12'hfff;
rom[98123] = 12'hfff;
rom[98124] = 12'hfff;
rom[98125] = 12'hfff;
rom[98126] = 12'hfff;
rom[98127] = 12'hfff;
rom[98128] = 12'hfff;
rom[98129] = 12'hfff;
rom[98130] = 12'hfff;
rom[98131] = 12'hfff;
rom[98132] = 12'hfff;
rom[98133] = 12'hfff;
rom[98134] = 12'hfff;
rom[98135] = 12'hfff;
rom[98136] = 12'hfff;
rom[98137] = 12'hfff;
rom[98138] = 12'hfff;
rom[98139] = 12'hfff;
rom[98140] = 12'hfff;
rom[98141] = 12'hfff;
rom[98142] = 12'hfff;
rom[98143] = 12'hfff;
rom[98144] = 12'hfff;
rom[98145] = 12'hfff;
rom[98146] = 12'hfff;
rom[98147] = 12'hfff;
rom[98148] = 12'hfff;
rom[98149] = 12'heee;
rom[98150] = 12'heee;
rom[98151] = 12'heee;
rom[98152] = 12'heee;
rom[98153] = 12'heee;
rom[98154] = 12'hddd;
rom[98155] = 12'hddd;
rom[98156] = 12'hddd;
rom[98157] = 12'hddd;
rom[98158] = 12'hddd;
rom[98159] = 12'hccc;
rom[98160] = 12'hddd;
rom[98161] = 12'hccc;
rom[98162] = 12'hccc;
rom[98163] = 12'hccc;
rom[98164] = 12'hccc;
rom[98165] = 12'hccc;
rom[98166] = 12'hccc;
rom[98167] = 12'hccc;
rom[98168] = 12'hccc;
rom[98169] = 12'hccc;
rom[98170] = 12'hccc;
rom[98171] = 12'hccc;
rom[98172] = 12'hccc;
rom[98173] = 12'hccc;
rom[98174] = 12'hccc;
rom[98175] = 12'hbbb;
rom[98176] = 12'hbbb;
rom[98177] = 12'hbbb;
rom[98178] = 12'hbbb;
rom[98179] = 12'hbbb;
rom[98180] = 12'haaa;
rom[98181] = 12'haaa;
rom[98182] = 12'haaa;
rom[98183] = 12'haaa;
rom[98184] = 12'haaa;
rom[98185] = 12'haaa;
rom[98186] = 12'haaa;
rom[98187] = 12'haaa;
rom[98188] = 12'h999;
rom[98189] = 12'h999;
rom[98190] = 12'h999;
rom[98191] = 12'h999;
rom[98192] = 12'haaa;
rom[98193] = 12'haaa;
rom[98194] = 12'haaa;
rom[98195] = 12'haaa;
rom[98196] = 12'haaa;
rom[98197] = 12'haaa;
rom[98198] = 12'haaa;
rom[98199] = 12'haaa;
rom[98200] = 12'haaa;
rom[98201] = 12'haaa;
rom[98202] = 12'haaa;
rom[98203] = 12'haaa;
rom[98204] = 12'haaa;
rom[98205] = 12'haaa;
rom[98206] = 12'haaa;
rom[98207] = 12'haaa;
rom[98208] = 12'haaa;
rom[98209] = 12'haaa;
rom[98210] = 12'haaa;
rom[98211] = 12'hbbb;
rom[98212] = 12'hbbb;
rom[98213] = 12'hbbb;
rom[98214] = 12'hbbb;
rom[98215] = 12'hbbb;
rom[98216] = 12'hbbb;
rom[98217] = 12'hbbb;
rom[98218] = 12'hbbb;
rom[98219] = 12'haaa;
rom[98220] = 12'haaa;
rom[98221] = 12'haaa;
rom[98222] = 12'h999;
rom[98223] = 12'h999;
rom[98224] = 12'h888;
rom[98225] = 12'h999;
rom[98226] = 12'h999;
rom[98227] = 12'h888;
rom[98228] = 12'h888;
rom[98229] = 12'h999;
rom[98230] = 12'h999;
rom[98231] = 12'h999;
rom[98232] = 12'haaa;
rom[98233] = 12'haaa;
rom[98234] = 12'haaa;
rom[98235] = 12'haaa;
rom[98236] = 12'haaa;
rom[98237] = 12'haaa;
rom[98238] = 12'haaa;
rom[98239] = 12'haaa;
rom[98240] = 12'haaa;
rom[98241] = 12'haaa;
rom[98242] = 12'h999;
rom[98243] = 12'h999;
rom[98244] = 12'h999;
rom[98245] = 12'h999;
rom[98246] = 12'h888;
rom[98247] = 12'h888;
rom[98248] = 12'h888;
rom[98249] = 12'h888;
rom[98250] = 12'h888;
rom[98251] = 12'h888;
rom[98252] = 12'h888;
rom[98253] = 12'h999;
rom[98254] = 12'h999;
rom[98255] = 12'h999;
rom[98256] = 12'haaa;
rom[98257] = 12'haaa;
rom[98258] = 12'haaa;
rom[98259] = 12'haaa;
rom[98260] = 12'haaa;
rom[98261] = 12'haaa;
rom[98262] = 12'h999;
rom[98263] = 12'h999;
rom[98264] = 12'h999;
rom[98265] = 12'h888;
rom[98266] = 12'h888;
rom[98267] = 12'h888;
rom[98268] = 12'h888;
rom[98269] = 12'h888;
rom[98270] = 12'h888;
rom[98271] = 12'h888;
rom[98272] = 12'h888;
rom[98273] = 12'h888;
rom[98274] = 12'h999;
rom[98275] = 12'h999;
rom[98276] = 12'h999;
rom[98277] = 12'h999;
rom[98278] = 12'h999;
rom[98279] = 12'h999;
rom[98280] = 12'h999;
rom[98281] = 12'haaa;
rom[98282] = 12'hbbb;
rom[98283] = 12'hccc;
rom[98284] = 12'hddd;
rom[98285] = 12'heee;
rom[98286] = 12'hfff;
rom[98287] = 12'hfff;
rom[98288] = 12'heee;
rom[98289] = 12'hddd;
rom[98290] = 12'hccc;
rom[98291] = 12'hbbb;
rom[98292] = 12'haaa;
rom[98293] = 12'h888;
rom[98294] = 12'h777;
rom[98295] = 12'h777;
rom[98296] = 12'h777;
rom[98297] = 12'h777;
rom[98298] = 12'h999;
rom[98299] = 12'haaa;
rom[98300] = 12'hccc;
rom[98301] = 12'heee;
rom[98302] = 12'hfff;
rom[98303] = 12'heee;
rom[98304] = 12'hccc;
rom[98305] = 12'h999;
rom[98306] = 12'h666;
rom[98307] = 12'h555;
rom[98308] = 12'h555;
rom[98309] = 12'h444;
rom[98310] = 12'h444;
rom[98311] = 12'h666;
rom[98312] = 12'h666;
rom[98313] = 12'h666;
rom[98314] = 12'h666;
rom[98315] = 12'h777;
rom[98316] = 12'h888;
rom[98317] = 12'h888;
rom[98318] = 12'h777;
rom[98319] = 12'h666;
rom[98320] = 12'h666;
rom[98321] = 12'h777;
rom[98322] = 12'h999;
rom[98323] = 12'hbbb;
rom[98324] = 12'hddd;
rom[98325] = 12'hfff;
rom[98326] = 12'hfff;
rom[98327] = 12'hfff;
rom[98328] = 12'heee;
rom[98329] = 12'hbbb;
rom[98330] = 12'h888;
rom[98331] = 12'h666;
rom[98332] = 12'h555;
rom[98333] = 12'h444;
rom[98334] = 12'h333;
rom[98335] = 12'h333;
rom[98336] = 12'h222;
rom[98337] = 12'h222;
rom[98338] = 12'h222;
rom[98339] = 12'h222;
rom[98340] = 12'h111;
rom[98341] = 12'h111;
rom[98342] = 12'h111;
rom[98343] = 12'h111;
rom[98344] = 12'h111;
rom[98345] = 12'h111;
rom[98346] = 12'h222;
rom[98347] = 12'h222;
rom[98348] = 12'h222;
rom[98349] = 12'h222;
rom[98350] = 12'h111;
rom[98351] = 12'h111;
rom[98352] = 12'h111;
rom[98353] = 12'h111;
rom[98354] = 12'h111;
rom[98355] = 12'h111;
rom[98356] = 12'h111;
rom[98357] = 12'h111;
rom[98358] = 12'h111;
rom[98359] = 12'h111;
rom[98360] = 12'h111;
rom[98361] = 12'h111;
rom[98362] = 12'h111;
rom[98363] = 12'h111;
rom[98364] = 12'h111;
rom[98365] = 12'h111;
rom[98366] = 12'h111;
rom[98367] = 12'h111;
rom[98368] = 12'h111;
rom[98369] = 12'h111;
rom[98370] = 12'h111;
rom[98371] = 12'h111;
rom[98372] = 12'h111;
rom[98373] = 12'h111;
rom[98374] = 12'h111;
rom[98375] = 12'h111;
rom[98376] = 12'h111;
rom[98377] = 12'h111;
rom[98378] = 12'h222;
rom[98379] = 12'h222;
rom[98380] = 12'h333;
rom[98381] = 12'h333;
rom[98382] = 12'h444;
rom[98383] = 12'h444;
rom[98384] = 12'h555;
rom[98385] = 12'h555;
rom[98386] = 12'h444;
rom[98387] = 12'h333;
rom[98388] = 12'h222;
rom[98389] = 12'h333;
rom[98390] = 12'h333;
rom[98391] = 12'h444;
rom[98392] = 12'h444;
rom[98393] = 12'h444;
rom[98394] = 12'h555;
rom[98395] = 12'h555;
rom[98396] = 12'h555;
rom[98397] = 12'h555;
rom[98398] = 12'h555;
rom[98399] = 12'h555;
rom[98400] = 12'hfff;
rom[98401] = 12'hfff;
rom[98402] = 12'hfff;
rom[98403] = 12'hfff;
rom[98404] = 12'hfff;
rom[98405] = 12'hfff;
rom[98406] = 12'hfff;
rom[98407] = 12'hfff;
rom[98408] = 12'hfff;
rom[98409] = 12'hfff;
rom[98410] = 12'hfff;
rom[98411] = 12'hfff;
rom[98412] = 12'hfff;
rom[98413] = 12'hfff;
rom[98414] = 12'hfff;
rom[98415] = 12'hfff;
rom[98416] = 12'hfff;
rom[98417] = 12'hfff;
rom[98418] = 12'hfff;
rom[98419] = 12'hfff;
rom[98420] = 12'hfff;
rom[98421] = 12'hfff;
rom[98422] = 12'hfff;
rom[98423] = 12'hfff;
rom[98424] = 12'hfff;
rom[98425] = 12'hfff;
rom[98426] = 12'hfff;
rom[98427] = 12'hfff;
rom[98428] = 12'hfff;
rom[98429] = 12'hfff;
rom[98430] = 12'hfff;
rom[98431] = 12'hfff;
rom[98432] = 12'hfff;
rom[98433] = 12'hfff;
rom[98434] = 12'hfff;
rom[98435] = 12'hfff;
rom[98436] = 12'hfff;
rom[98437] = 12'hfff;
rom[98438] = 12'hfff;
rom[98439] = 12'hfff;
rom[98440] = 12'hfff;
rom[98441] = 12'hfff;
rom[98442] = 12'hfff;
rom[98443] = 12'hfff;
rom[98444] = 12'hfff;
rom[98445] = 12'hfff;
rom[98446] = 12'hfff;
rom[98447] = 12'hfff;
rom[98448] = 12'hfff;
rom[98449] = 12'hfff;
rom[98450] = 12'hfff;
rom[98451] = 12'hfff;
rom[98452] = 12'hfff;
rom[98453] = 12'hfff;
rom[98454] = 12'hfff;
rom[98455] = 12'hfff;
rom[98456] = 12'hfff;
rom[98457] = 12'hfff;
rom[98458] = 12'hfff;
rom[98459] = 12'hfff;
rom[98460] = 12'hfff;
rom[98461] = 12'hfff;
rom[98462] = 12'hfff;
rom[98463] = 12'hfff;
rom[98464] = 12'hfff;
rom[98465] = 12'hfff;
rom[98466] = 12'hfff;
rom[98467] = 12'hfff;
rom[98468] = 12'hfff;
rom[98469] = 12'hfff;
rom[98470] = 12'hfff;
rom[98471] = 12'hfff;
rom[98472] = 12'hfff;
rom[98473] = 12'hfff;
rom[98474] = 12'hfff;
rom[98475] = 12'hfff;
rom[98476] = 12'hfff;
rom[98477] = 12'hfff;
rom[98478] = 12'hfff;
rom[98479] = 12'hfff;
rom[98480] = 12'hfff;
rom[98481] = 12'hfff;
rom[98482] = 12'hfff;
rom[98483] = 12'hfff;
rom[98484] = 12'hfff;
rom[98485] = 12'hfff;
rom[98486] = 12'hfff;
rom[98487] = 12'hfff;
rom[98488] = 12'hfff;
rom[98489] = 12'hfff;
rom[98490] = 12'hfff;
rom[98491] = 12'hfff;
rom[98492] = 12'hfff;
rom[98493] = 12'hfff;
rom[98494] = 12'hfff;
rom[98495] = 12'hfff;
rom[98496] = 12'hfff;
rom[98497] = 12'hfff;
rom[98498] = 12'hfff;
rom[98499] = 12'hfff;
rom[98500] = 12'hfff;
rom[98501] = 12'hfff;
rom[98502] = 12'hfff;
rom[98503] = 12'hfff;
rom[98504] = 12'hfff;
rom[98505] = 12'hfff;
rom[98506] = 12'hfff;
rom[98507] = 12'hfff;
rom[98508] = 12'hfff;
rom[98509] = 12'hfff;
rom[98510] = 12'hfff;
rom[98511] = 12'hfff;
rom[98512] = 12'hfff;
rom[98513] = 12'hfff;
rom[98514] = 12'hfff;
rom[98515] = 12'hfff;
rom[98516] = 12'hfff;
rom[98517] = 12'hfff;
rom[98518] = 12'hfff;
rom[98519] = 12'hfff;
rom[98520] = 12'hfff;
rom[98521] = 12'hfff;
rom[98522] = 12'hfff;
rom[98523] = 12'hfff;
rom[98524] = 12'hfff;
rom[98525] = 12'hfff;
rom[98526] = 12'hfff;
rom[98527] = 12'hfff;
rom[98528] = 12'hfff;
rom[98529] = 12'hfff;
rom[98530] = 12'hfff;
rom[98531] = 12'hfff;
rom[98532] = 12'hfff;
rom[98533] = 12'hfff;
rom[98534] = 12'hfff;
rom[98535] = 12'hfff;
rom[98536] = 12'hfff;
rom[98537] = 12'hfff;
rom[98538] = 12'hfff;
rom[98539] = 12'hfff;
rom[98540] = 12'hfff;
rom[98541] = 12'hfff;
rom[98542] = 12'hfff;
rom[98543] = 12'hfff;
rom[98544] = 12'hfff;
rom[98545] = 12'hfff;
rom[98546] = 12'hfff;
rom[98547] = 12'hfff;
rom[98548] = 12'hfff;
rom[98549] = 12'hfff;
rom[98550] = 12'hfff;
rom[98551] = 12'heee;
rom[98552] = 12'heee;
rom[98553] = 12'heee;
rom[98554] = 12'heee;
rom[98555] = 12'hddd;
rom[98556] = 12'hddd;
rom[98557] = 12'hddd;
rom[98558] = 12'hddd;
rom[98559] = 12'hddd;
rom[98560] = 12'hddd;
rom[98561] = 12'hddd;
rom[98562] = 12'hccc;
rom[98563] = 12'hccc;
rom[98564] = 12'hccc;
rom[98565] = 12'hccc;
rom[98566] = 12'hccc;
rom[98567] = 12'hccc;
rom[98568] = 12'hccc;
rom[98569] = 12'hccc;
rom[98570] = 12'hccc;
rom[98571] = 12'hccc;
rom[98572] = 12'hccc;
rom[98573] = 12'hccc;
rom[98574] = 12'hccc;
rom[98575] = 12'hccc;
rom[98576] = 12'hccc;
rom[98577] = 12'hbbb;
rom[98578] = 12'hbbb;
rom[98579] = 12'hbbb;
rom[98580] = 12'hbbb;
rom[98581] = 12'hbbb;
rom[98582] = 12'haaa;
rom[98583] = 12'haaa;
rom[98584] = 12'haaa;
rom[98585] = 12'haaa;
rom[98586] = 12'haaa;
rom[98587] = 12'haaa;
rom[98588] = 12'haaa;
rom[98589] = 12'haaa;
rom[98590] = 12'haaa;
rom[98591] = 12'haaa;
rom[98592] = 12'haaa;
rom[98593] = 12'haaa;
rom[98594] = 12'haaa;
rom[98595] = 12'haaa;
rom[98596] = 12'haaa;
rom[98597] = 12'haaa;
rom[98598] = 12'haaa;
rom[98599] = 12'haaa;
rom[98600] = 12'haaa;
rom[98601] = 12'haaa;
rom[98602] = 12'haaa;
rom[98603] = 12'haaa;
rom[98604] = 12'haaa;
rom[98605] = 12'haaa;
rom[98606] = 12'haaa;
rom[98607] = 12'haaa;
rom[98608] = 12'hbbb;
rom[98609] = 12'hbbb;
rom[98610] = 12'hbbb;
rom[98611] = 12'hbbb;
rom[98612] = 12'hbbb;
rom[98613] = 12'hbbb;
rom[98614] = 12'hbbb;
rom[98615] = 12'hbbb;
rom[98616] = 12'hbbb;
rom[98617] = 12'hbbb;
rom[98618] = 12'hbbb;
rom[98619] = 12'hbbb;
rom[98620] = 12'hbbb;
rom[98621] = 12'hbbb;
rom[98622] = 12'haaa;
rom[98623] = 12'haaa;
rom[98624] = 12'h999;
rom[98625] = 12'h999;
rom[98626] = 12'h999;
rom[98627] = 12'h999;
rom[98628] = 12'h999;
rom[98629] = 12'h999;
rom[98630] = 12'h999;
rom[98631] = 12'haaa;
rom[98632] = 12'haaa;
rom[98633] = 12'haaa;
rom[98634] = 12'haaa;
rom[98635] = 12'haaa;
rom[98636] = 12'haaa;
rom[98637] = 12'hbbb;
rom[98638] = 12'hbbb;
rom[98639] = 12'hbbb;
rom[98640] = 12'haaa;
rom[98641] = 12'haaa;
rom[98642] = 12'haaa;
rom[98643] = 12'haaa;
rom[98644] = 12'haaa;
rom[98645] = 12'h999;
rom[98646] = 12'h999;
rom[98647] = 12'h999;
rom[98648] = 12'h999;
rom[98649] = 12'h999;
rom[98650] = 12'h999;
rom[98651] = 12'h999;
rom[98652] = 12'haaa;
rom[98653] = 12'haaa;
rom[98654] = 12'haaa;
rom[98655] = 12'haaa;
rom[98656] = 12'hbbb;
rom[98657] = 12'hbbb;
rom[98658] = 12'haaa;
rom[98659] = 12'haaa;
rom[98660] = 12'haaa;
rom[98661] = 12'h999;
rom[98662] = 12'h999;
rom[98663] = 12'h999;
rom[98664] = 12'h999;
rom[98665] = 12'h999;
rom[98666] = 12'h999;
rom[98667] = 12'h999;
rom[98668] = 12'h999;
rom[98669] = 12'h888;
rom[98670] = 12'h888;
rom[98671] = 12'h888;
rom[98672] = 12'h999;
rom[98673] = 12'h999;
rom[98674] = 12'h999;
rom[98675] = 12'h999;
rom[98676] = 12'h999;
rom[98677] = 12'h999;
rom[98678] = 12'h999;
rom[98679] = 12'haaa;
rom[98680] = 12'haaa;
rom[98681] = 12'hbbb;
rom[98682] = 12'hddd;
rom[98683] = 12'heee;
rom[98684] = 12'hfff;
rom[98685] = 12'hfff;
rom[98686] = 12'hfff;
rom[98687] = 12'heee;
rom[98688] = 12'hddd;
rom[98689] = 12'hccc;
rom[98690] = 12'hbbb;
rom[98691] = 12'haaa;
rom[98692] = 12'h999;
rom[98693] = 12'h888;
rom[98694] = 12'h777;
rom[98695] = 12'h666;
rom[98696] = 12'h555;
rom[98697] = 12'h555;
rom[98698] = 12'h666;
rom[98699] = 12'h777;
rom[98700] = 12'h888;
rom[98701] = 12'hbbb;
rom[98702] = 12'hddd;
rom[98703] = 12'heee;
rom[98704] = 12'heee;
rom[98705] = 12'hccc;
rom[98706] = 12'haaa;
rom[98707] = 12'h888;
rom[98708] = 12'h666;
rom[98709] = 12'h444;
rom[98710] = 12'h444;
rom[98711] = 12'h555;
rom[98712] = 12'h555;
rom[98713] = 12'h555;
rom[98714] = 12'h555;
rom[98715] = 12'h666;
rom[98716] = 12'h777;
rom[98717] = 12'h777;
rom[98718] = 12'h777;
rom[98719] = 12'h777;
rom[98720] = 12'h555;
rom[98721] = 12'h444;
rom[98722] = 12'h555;
rom[98723] = 12'h666;
rom[98724] = 12'h999;
rom[98725] = 12'hbbb;
rom[98726] = 12'heee;
rom[98727] = 12'hfff;
rom[98728] = 12'hfff;
rom[98729] = 12'heee;
rom[98730] = 12'hccc;
rom[98731] = 12'haaa;
rom[98732] = 12'h888;
rom[98733] = 12'h666;
rom[98734] = 12'h444;
rom[98735] = 12'h333;
rom[98736] = 12'h333;
rom[98737] = 12'h333;
rom[98738] = 12'h222;
rom[98739] = 12'h222;
rom[98740] = 12'h222;
rom[98741] = 12'h111;
rom[98742] = 12'h111;
rom[98743] = 12'h111;
rom[98744] = 12'h111;
rom[98745] = 12'h111;
rom[98746] = 12'h111;
rom[98747] = 12'h111;
rom[98748] = 12'h222;
rom[98749] = 12'h222;
rom[98750] = 12'h111;
rom[98751] = 12'h111;
rom[98752] = 12'h111;
rom[98753] = 12'h111;
rom[98754] = 12'h111;
rom[98755] = 12'h111;
rom[98756] = 12'h111;
rom[98757] = 12'h111;
rom[98758] = 12'h111;
rom[98759] = 12'h111;
rom[98760] = 12'h111;
rom[98761] = 12'h111;
rom[98762] = 12'h111;
rom[98763] = 12'h111;
rom[98764] = 12'h111;
rom[98765] = 12'h111;
rom[98766] = 12'h111;
rom[98767] = 12'h111;
rom[98768] = 12'h111;
rom[98769] = 12'h111;
rom[98770] = 12'h111;
rom[98771] = 12'h111;
rom[98772] = 12'h111;
rom[98773] = 12'h111;
rom[98774] = 12'h111;
rom[98775] = 12'h111;
rom[98776] = 12'h111;
rom[98777] = 12'h111;
rom[98778] = 12'h111;
rom[98779] = 12'h222;
rom[98780] = 12'h222;
rom[98781] = 12'h222;
rom[98782] = 12'h333;
rom[98783] = 12'h333;
rom[98784] = 12'h444;
rom[98785] = 12'h444;
rom[98786] = 12'h444;
rom[98787] = 12'h333;
rom[98788] = 12'h333;
rom[98789] = 12'h222;
rom[98790] = 12'h222;
rom[98791] = 12'h222;
rom[98792] = 12'h333;
rom[98793] = 12'h333;
rom[98794] = 12'h333;
rom[98795] = 12'h333;
rom[98796] = 12'h444;
rom[98797] = 12'h444;
rom[98798] = 12'h444;
rom[98799] = 12'h555;
rom[98800] = 12'hfff;
rom[98801] = 12'hfff;
rom[98802] = 12'hfff;
rom[98803] = 12'hfff;
rom[98804] = 12'hfff;
rom[98805] = 12'hfff;
rom[98806] = 12'hfff;
rom[98807] = 12'hfff;
rom[98808] = 12'hfff;
rom[98809] = 12'hfff;
rom[98810] = 12'hfff;
rom[98811] = 12'hfff;
rom[98812] = 12'hfff;
rom[98813] = 12'hfff;
rom[98814] = 12'hfff;
rom[98815] = 12'hfff;
rom[98816] = 12'hfff;
rom[98817] = 12'hfff;
rom[98818] = 12'hfff;
rom[98819] = 12'hfff;
rom[98820] = 12'hfff;
rom[98821] = 12'hfff;
rom[98822] = 12'hfff;
rom[98823] = 12'hfff;
rom[98824] = 12'hfff;
rom[98825] = 12'hfff;
rom[98826] = 12'hfff;
rom[98827] = 12'hfff;
rom[98828] = 12'hfff;
rom[98829] = 12'hfff;
rom[98830] = 12'hfff;
rom[98831] = 12'hfff;
rom[98832] = 12'hfff;
rom[98833] = 12'hfff;
rom[98834] = 12'hfff;
rom[98835] = 12'hfff;
rom[98836] = 12'hfff;
rom[98837] = 12'hfff;
rom[98838] = 12'hfff;
rom[98839] = 12'hfff;
rom[98840] = 12'hfff;
rom[98841] = 12'hfff;
rom[98842] = 12'hfff;
rom[98843] = 12'hfff;
rom[98844] = 12'hfff;
rom[98845] = 12'hfff;
rom[98846] = 12'hfff;
rom[98847] = 12'hfff;
rom[98848] = 12'hfff;
rom[98849] = 12'hfff;
rom[98850] = 12'hfff;
rom[98851] = 12'hfff;
rom[98852] = 12'hfff;
rom[98853] = 12'hfff;
rom[98854] = 12'hfff;
rom[98855] = 12'hfff;
rom[98856] = 12'hfff;
rom[98857] = 12'hfff;
rom[98858] = 12'hfff;
rom[98859] = 12'hfff;
rom[98860] = 12'hfff;
rom[98861] = 12'hfff;
rom[98862] = 12'hfff;
rom[98863] = 12'hfff;
rom[98864] = 12'hfff;
rom[98865] = 12'hfff;
rom[98866] = 12'hfff;
rom[98867] = 12'hfff;
rom[98868] = 12'hfff;
rom[98869] = 12'hfff;
rom[98870] = 12'hfff;
rom[98871] = 12'hfff;
rom[98872] = 12'hfff;
rom[98873] = 12'hfff;
rom[98874] = 12'hfff;
rom[98875] = 12'hfff;
rom[98876] = 12'hfff;
rom[98877] = 12'hfff;
rom[98878] = 12'hfff;
rom[98879] = 12'hfff;
rom[98880] = 12'hfff;
rom[98881] = 12'hfff;
rom[98882] = 12'hfff;
rom[98883] = 12'hfff;
rom[98884] = 12'hfff;
rom[98885] = 12'hfff;
rom[98886] = 12'hfff;
rom[98887] = 12'hfff;
rom[98888] = 12'hfff;
rom[98889] = 12'hfff;
rom[98890] = 12'hfff;
rom[98891] = 12'hfff;
rom[98892] = 12'hfff;
rom[98893] = 12'hfff;
rom[98894] = 12'hfff;
rom[98895] = 12'hfff;
rom[98896] = 12'hfff;
rom[98897] = 12'hfff;
rom[98898] = 12'hfff;
rom[98899] = 12'hfff;
rom[98900] = 12'hfff;
rom[98901] = 12'hfff;
rom[98902] = 12'hfff;
rom[98903] = 12'hfff;
rom[98904] = 12'hfff;
rom[98905] = 12'hfff;
rom[98906] = 12'hfff;
rom[98907] = 12'hfff;
rom[98908] = 12'hfff;
rom[98909] = 12'hfff;
rom[98910] = 12'hfff;
rom[98911] = 12'hfff;
rom[98912] = 12'hfff;
rom[98913] = 12'hfff;
rom[98914] = 12'hfff;
rom[98915] = 12'hfff;
rom[98916] = 12'hfff;
rom[98917] = 12'hfff;
rom[98918] = 12'hfff;
rom[98919] = 12'hfff;
rom[98920] = 12'hfff;
rom[98921] = 12'hfff;
rom[98922] = 12'hfff;
rom[98923] = 12'hfff;
rom[98924] = 12'hfff;
rom[98925] = 12'hfff;
rom[98926] = 12'hfff;
rom[98927] = 12'hfff;
rom[98928] = 12'hfff;
rom[98929] = 12'hfff;
rom[98930] = 12'hfff;
rom[98931] = 12'hfff;
rom[98932] = 12'hfff;
rom[98933] = 12'hfff;
rom[98934] = 12'hfff;
rom[98935] = 12'hfff;
rom[98936] = 12'hfff;
rom[98937] = 12'hfff;
rom[98938] = 12'hfff;
rom[98939] = 12'hfff;
rom[98940] = 12'hfff;
rom[98941] = 12'hfff;
rom[98942] = 12'hfff;
rom[98943] = 12'hfff;
rom[98944] = 12'hfff;
rom[98945] = 12'hfff;
rom[98946] = 12'hfff;
rom[98947] = 12'hfff;
rom[98948] = 12'hfff;
rom[98949] = 12'hfff;
rom[98950] = 12'hfff;
rom[98951] = 12'hfff;
rom[98952] = 12'heee;
rom[98953] = 12'heee;
rom[98954] = 12'heee;
rom[98955] = 12'heee;
rom[98956] = 12'hddd;
rom[98957] = 12'hddd;
rom[98958] = 12'hddd;
rom[98959] = 12'hddd;
rom[98960] = 12'hddd;
rom[98961] = 12'hddd;
rom[98962] = 12'hddd;
rom[98963] = 12'hddd;
rom[98964] = 12'hddd;
rom[98965] = 12'hddd;
rom[98966] = 12'hddd;
rom[98967] = 12'hddd;
rom[98968] = 12'hddd;
rom[98969] = 12'hccc;
rom[98970] = 12'hccc;
rom[98971] = 12'hccc;
rom[98972] = 12'hccc;
rom[98973] = 12'hccc;
rom[98974] = 12'hccc;
rom[98975] = 12'hccc;
rom[98976] = 12'hccc;
rom[98977] = 12'hccc;
rom[98978] = 12'hccc;
rom[98979] = 12'hbbb;
rom[98980] = 12'hbbb;
rom[98981] = 12'hbbb;
rom[98982] = 12'hbbb;
rom[98983] = 12'haaa;
rom[98984] = 12'hbbb;
rom[98985] = 12'haaa;
rom[98986] = 12'haaa;
rom[98987] = 12'haaa;
rom[98988] = 12'haaa;
rom[98989] = 12'haaa;
rom[98990] = 12'haaa;
rom[98991] = 12'haaa;
rom[98992] = 12'haaa;
rom[98993] = 12'haaa;
rom[98994] = 12'haaa;
rom[98995] = 12'haaa;
rom[98996] = 12'haaa;
rom[98997] = 12'haaa;
rom[98998] = 12'haaa;
rom[98999] = 12'haaa;
rom[99000] = 12'haaa;
rom[99001] = 12'haaa;
rom[99002] = 12'haaa;
rom[99003] = 12'haaa;
rom[99004] = 12'haaa;
rom[99005] = 12'haaa;
rom[99006] = 12'hbbb;
rom[99007] = 12'hbbb;
rom[99008] = 12'hbbb;
rom[99009] = 12'hbbb;
rom[99010] = 12'hbbb;
rom[99011] = 12'hbbb;
rom[99012] = 12'hbbb;
rom[99013] = 12'hbbb;
rom[99014] = 12'hbbb;
rom[99015] = 12'hbbb;
rom[99016] = 12'hccc;
rom[99017] = 12'hccc;
rom[99018] = 12'hccc;
rom[99019] = 12'hccc;
rom[99020] = 12'hccc;
rom[99021] = 12'hccc;
rom[99022] = 12'hbbb;
rom[99023] = 12'hbbb;
rom[99024] = 12'haaa;
rom[99025] = 12'haaa;
rom[99026] = 12'haaa;
rom[99027] = 12'h999;
rom[99028] = 12'h999;
rom[99029] = 12'h999;
rom[99030] = 12'h999;
rom[99031] = 12'haaa;
rom[99032] = 12'haaa;
rom[99033] = 12'haaa;
rom[99034] = 12'haaa;
rom[99035] = 12'haaa;
rom[99036] = 12'hbbb;
rom[99037] = 12'hbbb;
rom[99038] = 12'hbbb;
rom[99039] = 12'hbbb;
rom[99040] = 12'hbbb;
rom[99041] = 12'haaa;
rom[99042] = 12'haaa;
rom[99043] = 12'haaa;
rom[99044] = 12'haaa;
rom[99045] = 12'haaa;
rom[99046] = 12'haaa;
rom[99047] = 12'h999;
rom[99048] = 12'h999;
rom[99049] = 12'h999;
rom[99050] = 12'haaa;
rom[99051] = 12'haaa;
rom[99052] = 12'hbbb;
rom[99053] = 12'hbbb;
rom[99054] = 12'hbbb;
rom[99055] = 12'hbbb;
rom[99056] = 12'haaa;
rom[99057] = 12'haaa;
rom[99058] = 12'haaa;
rom[99059] = 12'haaa;
rom[99060] = 12'haaa;
rom[99061] = 12'h999;
rom[99062] = 12'h999;
rom[99063] = 12'h999;
rom[99064] = 12'h999;
rom[99065] = 12'h999;
rom[99066] = 12'h999;
rom[99067] = 12'h999;
rom[99068] = 12'h999;
rom[99069] = 12'h999;
rom[99070] = 12'h999;
rom[99071] = 12'h999;
rom[99072] = 12'h999;
rom[99073] = 12'h999;
rom[99074] = 12'h999;
rom[99075] = 12'h999;
rom[99076] = 12'h999;
rom[99077] = 12'haaa;
rom[99078] = 12'haaa;
rom[99079] = 12'haaa;
rom[99080] = 12'hbbb;
rom[99081] = 12'hccc;
rom[99082] = 12'heee;
rom[99083] = 12'hfff;
rom[99084] = 12'hfff;
rom[99085] = 12'hfff;
rom[99086] = 12'heee;
rom[99087] = 12'hddd;
rom[99088] = 12'hccc;
rom[99089] = 12'hbbb;
rom[99090] = 12'haaa;
rom[99091] = 12'h999;
rom[99092] = 12'h888;
rom[99093] = 12'h777;
rom[99094] = 12'h666;
rom[99095] = 12'h666;
rom[99096] = 12'h555;
rom[99097] = 12'h555;
rom[99098] = 12'h555;
rom[99099] = 12'h444;
rom[99100] = 12'h555;
rom[99101] = 12'h777;
rom[99102] = 12'haaa;
rom[99103] = 12'hccc;
rom[99104] = 12'hfff;
rom[99105] = 12'hfff;
rom[99106] = 12'hddd;
rom[99107] = 12'hbbb;
rom[99108] = 12'h888;
rom[99109] = 12'h666;
rom[99110] = 12'h555;
rom[99111] = 12'h444;
rom[99112] = 12'h555;
rom[99113] = 12'h555;
rom[99114] = 12'h555;
rom[99115] = 12'h555;
rom[99116] = 12'h666;
rom[99117] = 12'h666;
rom[99118] = 12'h777;
rom[99119] = 12'h888;
rom[99120] = 12'h777;
rom[99121] = 12'h555;
rom[99122] = 12'h333;
rom[99123] = 12'h333;
rom[99124] = 12'h555;
rom[99125] = 12'h777;
rom[99126] = 12'haaa;
rom[99127] = 12'hccc;
rom[99128] = 12'heee;
rom[99129] = 12'hfff;
rom[99130] = 12'hfff;
rom[99131] = 12'heee;
rom[99132] = 12'hbbb;
rom[99133] = 12'h888;
rom[99134] = 12'h666;
rom[99135] = 12'h555;
rom[99136] = 12'h555;
rom[99137] = 12'h444;
rom[99138] = 12'h333;
rom[99139] = 12'h222;
rom[99140] = 12'h222;
rom[99141] = 12'h111;
rom[99142] = 12'h111;
rom[99143] = 12'h111;
rom[99144] = 12'h111;
rom[99145] = 12'h111;
rom[99146] = 12'h111;
rom[99147] = 12'h111;
rom[99148] = 12'h222;
rom[99149] = 12'h222;
rom[99150] = 12'h222;
rom[99151] = 12'h111;
rom[99152] = 12'h111;
rom[99153] = 12'h111;
rom[99154] = 12'h111;
rom[99155] = 12'h111;
rom[99156] = 12'h111;
rom[99157] = 12'h111;
rom[99158] = 12'h111;
rom[99159] = 12'h111;
rom[99160] = 12'h111;
rom[99161] = 12'h111;
rom[99162] = 12'h111;
rom[99163] = 12'h111;
rom[99164] = 12'h111;
rom[99165] = 12'h111;
rom[99166] = 12'h111;
rom[99167] = 12'h111;
rom[99168] = 12'h111;
rom[99169] = 12'h111;
rom[99170] = 12'h111;
rom[99171] = 12'h111;
rom[99172] = 12'h111;
rom[99173] = 12'h111;
rom[99174] = 12'h111;
rom[99175] = 12'h111;
rom[99176] = 12'h111;
rom[99177] = 12'h111;
rom[99178] = 12'h111;
rom[99179] = 12'h111;
rom[99180] = 12'h111;
rom[99181] = 12'h222;
rom[99182] = 12'h222;
rom[99183] = 12'h333;
rom[99184] = 12'h333;
rom[99185] = 12'h444;
rom[99186] = 12'h444;
rom[99187] = 12'h444;
rom[99188] = 12'h333;
rom[99189] = 12'h333;
rom[99190] = 12'h222;
rom[99191] = 12'h222;
rom[99192] = 12'h222;
rom[99193] = 12'h222;
rom[99194] = 12'h222;
rom[99195] = 12'h222;
rom[99196] = 12'h333;
rom[99197] = 12'h333;
rom[99198] = 12'h333;
rom[99199] = 12'h444;
rom[99200] = 12'hfff;
rom[99201] = 12'hfff;
rom[99202] = 12'hfff;
rom[99203] = 12'hfff;
rom[99204] = 12'hfff;
rom[99205] = 12'hfff;
rom[99206] = 12'hfff;
rom[99207] = 12'hfff;
rom[99208] = 12'hfff;
rom[99209] = 12'hfff;
rom[99210] = 12'hfff;
rom[99211] = 12'hfff;
rom[99212] = 12'hfff;
rom[99213] = 12'hfff;
rom[99214] = 12'hfff;
rom[99215] = 12'hfff;
rom[99216] = 12'hfff;
rom[99217] = 12'hfff;
rom[99218] = 12'hfff;
rom[99219] = 12'hfff;
rom[99220] = 12'hfff;
rom[99221] = 12'hfff;
rom[99222] = 12'hfff;
rom[99223] = 12'hfff;
rom[99224] = 12'hfff;
rom[99225] = 12'hfff;
rom[99226] = 12'hfff;
rom[99227] = 12'hfff;
rom[99228] = 12'hfff;
rom[99229] = 12'hfff;
rom[99230] = 12'hfff;
rom[99231] = 12'hfff;
rom[99232] = 12'hfff;
rom[99233] = 12'hfff;
rom[99234] = 12'hfff;
rom[99235] = 12'hfff;
rom[99236] = 12'hfff;
rom[99237] = 12'hfff;
rom[99238] = 12'hfff;
rom[99239] = 12'hfff;
rom[99240] = 12'hfff;
rom[99241] = 12'hfff;
rom[99242] = 12'hfff;
rom[99243] = 12'hfff;
rom[99244] = 12'hfff;
rom[99245] = 12'hfff;
rom[99246] = 12'hfff;
rom[99247] = 12'hfff;
rom[99248] = 12'hfff;
rom[99249] = 12'hfff;
rom[99250] = 12'hfff;
rom[99251] = 12'hfff;
rom[99252] = 12'hfff;
rom[99253] = 12'hfff;
rom[99254] = 12'hfff;
rom[99255] = 12'hfff;
rom[99256] = 12'hfff;
rom[99257] = 12'hfff;
rom[99258] = 12'hfff;
rom[99259] = 12'hfff;
rom[99260] = 12'hfff;
rom[99261] = 12'hfff;
rom[99262] = 12'hfff;
rom[99263] = 12'hfff;
rom[99264] = 12'hfff;
rom[99265] = 12'hfff;
rom[99266] = 12'hfff;
rom[99267] = 12'hfff;
rom[99268] = 12'hfff;
rom[99269] = 12'hfff;
rom[99270] = 12'hfff;
rom[99271] = 12'hfff;
rom[99272] = 12'hfff;
rom[99273] = 12'hfff;
rom[99274] = 12'hfff;
rom[99275] = 12'hfff;
rom[99276] = 12'hfff;
rom[99277] = 12'hfff;
rom[99278] = 12'hfff;
rom[99279] = 12'hfff;
rom[99280] = 12'hfff;
rom[99281] = 12'hfff;
rom[99282] = 12'hfff;
rom[99283] = 12'heee;
rom[99284] = 12'hfff;
rom[99285] = 12'hfff;
rom[99286] = 12'hfff;
rom[99287] = 12'hfff;
rom[99288] = 12'hfff;
rom[99289] = 12'hfff;
rom[99290] = 12'hfff;
rom[99291] = 12'hfff;
rom[99292] = 12'hfff;
rom[99293] = 12'hfff;
rom[99294] = 12'hfff;
rom[99295] = 12'hfff;
rom[99296] = 12'hfff;
rom[99297] = 12'hfff;
rom[99298] = 12'hfff;
rom[99299] = 12'hfff;
rom[99300] = 12'hfff;
rom[99301] = 12'hfff;
rom[99302] = 12'hfff;
rom[99303] = 12'hfff;
rom[99304] = 12'hfff;
rom[99305] = 12'hfff;
rom[99306] = 12'hfff;
rom[99307] = 12'hfff;
rom[99308] = 12'hfff;
rom[99309] = 12'hfff;
rom[99310] = 12'hfff;
rom[99311] = 12'hfff;
rom[99312] = 12'hfff;
rom[99313] = 12'hfff;
rom[99314] = 12'hfff;
rom[99315] = 12'hfff;
rom[99316] = 12'hfff;
rom[99317] = 12'hfff;
rom[99318] = 12'hfff;
rom[99319] = 12'hfff;
rom[99320] = 12'hfff;
rom[99321] = 12'hfff;
rom[99322] = 12'hfff;
rom[99323] = 12'hfff;
rom[99324] = 12'hfff;
rom[99325] = 12'hfff;
rom[99326] = 12'hfff;
rom[99327] = 12'hfff;
rom[99328] = 12'hfff;
rom[99329] = 12'hfff;
rom[99330] = 12'hfff;
rom[99331] = 12'hfff;
rom[99332] = 12'hfff;
rom[99333] = 12'hfff;
rom[99334] = 12'hfff;
rom[99335] = 12'hfff;
rom[99336] = 12'hfff;
rom[99337] = 12'hfff;
rom[99338] = 12'hfff;
rom[99339] = 12'hfff;
rom[99340] = 12'hfff;
rom[99341] = 12'hfff;
rom[99342] = 12'hfff;
rom[99343] = 12'hfff;
rom[99344] = 12'hfff;
rom[99345] = 12'hfff;
rom[99346] = 12'hfff;
rom[99347] = 12'hfff;
rom[99348] = 12'hfff;
rom[99349] = 12'hfff;
rom[99350] = 12'hfff;
rom[99351] = 12'hfff;
rom[99352] = 12'hfff;
rom[99353] = 12'hfff;
rom[99354] = 12'hfff;
rom[99355] = 12'heee;
rom[99356] = 12'heee;
rom[99357] = 12'heee;
rom[99358] = 12'heee;
rom[99359] = 12'hddd;
rom[99360] = 12'hddd;
rom[99361] = 12'hddd;
rom[99362] = 12'hddd;
rom[99363] = 12'hddd;
rom[99364] = 12'hddd;
rom[99365] = 12'hddd;
rom[99366] = 12'hddd;
rom[99367] = 12'hddd;
rom[99368] = 12'hddd;
rom[99369] = 12'hddd;
rom[99370] = 12'hccc;
rom[99371] = 12'hccc;
rom[99372] = 12'hccc;
rom[99373] = 12'hccc;
rom[99374] = 12'hccc;
rom[99375] = 12'hccc;
rom[99376] = 12'hccc;
rom[99377] = 12'hccc;
rom[99378] = 12'hccc;
rom[99379] = 12'hccc;
rom[99380] = 12'hbbb;
rom[99381] = 12'hbbb;
rom[99382] = 12'hbbb;
rom[99383] = 12'hbbb;
rom[99384] = 12'hbbb;
rom[99385] = 12'hbbb;
rom[99386] = 12'hbbb;
rom[99387] = 12'hbbb;
rom[99388] = 12'hbbb;
rom[99389] = 12'hbbb;
rom[99390] = 12'hbbb;
rom[99391] = 12'hbbb;
rom[99392] = 12'hbbb;
rom[99393] = 12'hbbb;
rom[99394] = 12'hbbb;
rom[99395] = 12'hbbb;
rom[99396] = 12'hbbb;
rom[99397] = 12'hbbb;
rom[99398] = 12'hbbb;
rom[99399] = 12'hbbb;
rom[99400] = 12'hbbb;
rom[99401] = 12'hbbb;
rom[99402] = 12'hbbb;
rom[99403] = 12'hbbb;
rom[99404] = 12'hbbb;
rom[99405] = 12'hbbb;
rom[99406] = 12'hbbb;
rom[99407] = 12'hbbb;
rom[99408] = 12'hbbb;
rom[99409] = 12'hbbb;
rom[99410] = 12'hbbb;
rom[99411] = 12'hbbb;
rom[99412] = 12'hbbb;
rom[99413] = 12'hbbb;
rom[99414] = 12'hbbb;
rom[99415] = 12'hccc;
rom[99416] = 12'hccc;
rom[99417] = 12'hccc;
rom[99418] = 12'hccc;
rom[99419] = 12'hccc;
rom[99420] = 12'hccc;
rom[99421] = 12'hccc;
rom[99422] = 12'hccc;
rom[99423] = 12'hccc;
rom[99424] = 12'hccc;
rom[99425] = 12'hbbb;
rom[99426] = 12'hbbb;
rom[99427] = 12'haaa;
rom[99428] = 12'haaa;
rom[99429] = 12'haaa;
rom[99430] = 12'haaa;
rom[99431] = 12'haaa;
rom[99432] = 12'hbbb;
rom[99433] = 12'hbbb;
rom[99434] = 12'haaa;
rom[99435] = 12'haaa;
rom[99436] = 12'hbbb;
rom[99437] = 12'hbbb;
rom[99438] = 12'hbbb;
rom[99439] = 12'hbbb;
rom[99440] = 12'hbbb;
rom[99441] = 12'hbbb;
rom[99442] = 12'haaa;
rom[99443] = 12'haaa;
rom[99444] = 12'hbbb;
rom[99445] = 12'hbbb;
rom[99446] = 12'hbbb;
rom[99447] = 12'hbbb;
rom[99448] = 12'hbbb;
rom[99449] = 12'hbbb;
rom[99450] = 12'hbbb;
rom[99451] = 12'hbbb;
rom[99452] = 12'hbbb;
rom[99453] = 12'hbbb;
rom[99454] = 12'hbbb;
rom[99455] = 12'hbbb;
rom[99456] = 12'haaa;
rom[99457] = 12'haaa;
rom[99458] = 12'haaa;
rom[99459] = 12'haaa;
rom[99460] = 12'h999;
rom[99461] = 12'h999;
rom[99462] = 12'h999;
rom[99463] = 12'h999;
rom[99464] = 12'h999;
rom[99465] = 12'h999;
rom[99466] = 12'haaa;
rom[99467] = 12'haaa;
rom[99468] = 12'haaa;
rom[99469] = 12'h999;
rom[99470] = 12'h999;
rom[99471] = 12'h999;
rom[99472] = 12'h999;
rom[99473] = 12'haaa;
rom[99474] = 12'haaa;
rom[99475] = 12'haaa;
rom[99476] = 12'haaa;
rom[99477] = 12'hbbb;
rom[99478] = 12'hccc;
rom[99479] = 12'hccc;
rom[99480] = 12'heee;
rom[99481] = 12'heee;
rom[99482] = 12'hfff;
rom[99483] = 12'hfff;
rom[99484] = 12'hfff;
rom[99485] = 12'heee;
rom[99486] = 12'hccc;
rom[99487] = 12'hbbb;
rom[99488] = 12'haaa;
rom[99489] = 12'haaa;
rom[99490] = 12'haaa;
rom[99491] = 12'h999;
rom[99492] = 12'h888;
rom[99493] = 12'h777;
rom[99494] = 12'h666;
rom[99495] = 12'h555;
rom[99496] = 12'h555;
rom[99497] = 12'h444;
rom[99498] = 12'h444;
rom[99499] = 12'h444;
rom[99500] = 12'h444;
rom[99501] = 12'h444;
rom[99502] = 12'h555;
rom[99503] = 12'h777;
rom[99504] = 12'haaa;
rom[99505] = 12'hddd;
rom[99506] = 12'heee;
rom[99507] = 12'heee;
rom[99508] = 12'hccc;
rom[99509] = 12'haaa;
rom[99510] = 12'h777;
rom[99511] = 12'h555;
rom[99512] = 12'h444;
rom[99513] = 12'h444;
rom[99514] = 12'h555;
rom[99515] = 12'h555;
rom[99516] = 12'h666;
rom[99517] = 12'h666;
rom[99518] = 12'h777;
rom[99519] = 12'h888;
rom[99520] = 12'h666;
rom[99521] = 12'h666;
rom[99522] = 12'h444;
rom[99523] = 12'h333;
rom[99524] = 12'h333;
rom[99525] = 12'h444;
rom[99526] = 12'h555;
rom[99527] = 12'h777;
rom[99528] = 12'h999;
rom[99529] = 12'hccc;
rom[99530] = 12'hfff;
rom[99531] = 12'hfff;
rom[99532] = 12'hfff;
rom[99533] = 12'hddd;
rom[99534] = 12'hbbb;
rom[99535] = 12'h888;
rom[99536] = 12'h666;
rom[99537] = 12'h555;
rom[99538] = 12'h444;
rom[99539] = 12'h333;
rom[99540] = 12'h333;
rom[99541] = 12'h222;
rom[99542] = 12'h222;
rom[99543] = 12'h222;
rom[99544] = 12'h111;
rom[99545] = 12'h111;
rom[99546] = 12'h111;
rom[99547] = 12'h  0;
rom[99548] = 12'h  0;
rom[99549] = 12'h111;
rom[99550] = 12'h111;
rom[99551] = 12'h222;
rom[99552] = 12'h111;
rom[99553] = 12'h111;
rom[99554] = 12'h111;
rom[99555] = 12'h111;
rom[99556] = 12'h111;
rom[99557] = 12'h111;
rom[99558] = 12'h111;
rom[99559] = 12'h111;
rom[99560] = 12'h111;
rom[99561] = 12'h111;
rom[99562] = 12'h111;
rom[99563] = 12'h111;
rom[99564] = 12'h111;
rom[99565] = 12'h111;
rom[99566] = 12'h111;
rom[99567] = 12'h111;
rom[99568] = 12'h111;
rom[99569] = 12'h111;
rom[99570] = 12'h111;
rom[99571] = 12'h111;
rom[99572] = 12'h111;
rom[99573] = 12'h111;
rom[99574] = 12'h111;
rom[99575] = 12'h111;
rom[99576] = 12'h111;
rom[99577] = 12'h111;
rom[99578] = 12'h111;
rom[99579] = 12'h111;
rom[99580] = 12'h111;
rom[99581] = 12'h111;
rom[99582] = 12'h111;
rom[99583] = 12'h222;
rom[99584] = 12'h333;
rom[99585] = 12'h333;
rom[99586] = 12'h333;
rom[99587] = 12'h444;
rom[99588] = 12'h444;
rom[99589] = 12'h333;
rom[99590] = 12'h222;
rom[99591] = 12'h111;
rom[99592] = 12'h111;
rom[99593] = 12'h111;
rom[99594] = 12'h111;
rom[99595] = 12'h111;
rom[99596] = 12'h222;
rom[99597] = 12'h222;
rom[99598] = 12'h222;
rom[99599] = 12'h222;
rom[99600] = 12'hfff;
rom[99601] = 12'hfff;
rom[99602] = 12'hfff;
rom[99603] = 12'hfff;
rom[99604] = 12'hfff;
rom[99605] = 12'hfff;
rom[99606] = 12'hfff;
rom[99607] = 12'hfff;
rom[99608] = 12'hfff;
rom[99609] = 12'hfff;
rom[99610] = 12'hfff;
rom[99611] = 12'hfff;
rom[99612] = 12'hfff;
rom[99613] = 12'hfff;
rom[99614] = 12'hfff;
rom[99615] = 12'hfff;
rom[99616] = 12'hfff;
rom[99617] = 12'hfff;
rom[99618] = 12'hfff;
rom[99619] = 12'hfff;
rom[99620] = 12'hfff;
rom[99621] = 12'hfff;
rom[99622] = 12'hfff;
rom[99623] = 12'hfff;
rom[99624] = 12'hfff;
rom[99625] = 12'hfff;
rom[99626] = 12'hfff;
rom[99627] = 12'hfff;
rom[99628] = 12'hfff;
rom[99629] = 12'hfff;
rom[99630] = 12'hfff;
rom[99631] = 12'hfff;
rom[99632] = 12'hfff;
rom[99633] = 12'hfff;
rom[99634] = 12'hfff;
rom[99635] = 12'hfff;
rom[99636] = 12'hfff;
rom[99637] = 12'hfff;
rom[99638] = 12'hfff;
rom[99639] = 12'hfff;
rom[99640] = 12'hfff;
rom[99641] = 12'hfff;
rom[99642] = 12'hfff;
rom[99643] = 12'hfff;
rom[99644] = 12'hfff;
rom[99645] = 12'hfff;
rom[99646] = 12'hfff;
rom[99647] = 12'hfff;
rom[99648] = 12'hfff;
rom[99649] = 12'hfff;
rom[99650] = 12'hfff;
rom[99651] = 12'hfff;
rom[99652] = 12'hfff;
rom[99653] = 12'hfff;
rom[99654] = 12'hfff;
rom[99655] = 12'hfff;
rom[99656] = 12'hfff;
rom[99657] = 12'hfff;
rom[99658] = 12'hfff;
rom[99659] = 12'hfff;
rom[99660] = 12'hfff;
rom[99661] = 12'hfff;
rom[99662] = 12'hfff;
rom[99663] = 12'hfff;
rom[99664] = 12'hfff;
rom[99665] = 12'hfff;
rom[99666] = 12'hfff;
rom[99667] = 12'hfff;
rom[99668] = 12'hfff;
rom[99669] = 12'hfff;
rom[99670] = 12'hfff;
rom[99671] = 12'hfff;
rom[99672] = 12'hfff;
rom[99673] = 12'hfff;
rom[99674] = 12'hfff;
rom[99675] = 12'hfff;
rom[99676] = 12'hfff;
rom[99677] = 12'hfff;
rom[99678] = 12'hfff;
rom[99679] = 12'hfff;
rom[99680] = 12'hfff;
rom[99681] = 12'hfff;
rom[99682] = 12'hfff;
rom[99683] = 12'heee;
rom[99684] = 12'hfff;
rom[99685] = 12'hfff;
rom[99686] = 12'hfff;
rom[99687] = 12'hfff;
rom[99688] = 12'hfff;
rom[99689] = 12'hfff;
rom[99690] = 12'hfff;
rom[99691] = 12'hfff;
rom[99692] = 12'hfff;
rom[99693] = 12'hfff;
rom[99694] = 12'hfff;
rom[99695] = 12'hfff;
rom[99696] = 12'hfff;
rom[99697] = 12'hfff;
rom[99698] = 12'hfff;
rom[99699] = 12'hfff;
rom[99700] = 12'hfff;
rom[99701] = 12'hfff;
rom[99702] = 12'hfff;
rom[99703] = 12'hfff;
rom[99704] = 12'hfff;
rom[99705] = 12'hfff;
rom[99706] = 12'hfff;
rom[99707] = 12'hfff;
rom[99708] = 12'hfff;
rom[99709] = 12'hfff;
rom[99710] = 12'hfff;
rom[99711] = 12'hfff;
rom[99712] = 12'hfff;
rom[99713] = 12'hfff;
rom[99714] = 12'hfff;
rom[99715] = 12'hfff;
rom[99716] = 12'hfff;
rom[99717] = 12'hfff;
rom[99718] = 12'hfff;
rom[99719] = 12'hfff;
rom[99720] = 12'hfff;
rom[99721] = 12'hfff;
rom[99722] = 12'hfff;
rom[99723] = 12'hfff;
rom[99724] = 12'hfff;
rom[99725] = 12'hfff;
rom[99726] = 12'hfff;
rom[99727] = 12'hfff;
rom[99728] = 12'hfff;
rom[99729] = 12'hfff;
rom[99730] = 12'hfff;
rom[99731] = 12'hfff;
rom[99732] = 12'hfff;
rom[99733] = 12'hfff;
rom[99734] = 12'hfff;
rom[99735] = 12'hfff;
rom[99736] = 12'hfff;
rom[99737] = 12'hfff;
rom[99738] = 12'hfff;
rom[99739] = 12'hfff;
rom[99740] = 12'hfff;
rom[99741] = 12'hfff;
rom[99742] = 12'hfff;
rom[99743] = 12'hfff;
rom[99744] = 12'hfff;
rom[99745] = 12'hfff;
rom[99746] = 12'hfff;
rom[99747] = 12'hfff;
rom[99748] = 12'hfff;
rom[99749] = 12'hfff;
rom[99750] = 12'hfff;
rom[99751] = 12'hfff;
rom[99752] = 12'hfff;
rom[99753] = 12'hfff;
rom[99754] = 12'hfff;
rom[99755] = 12'hfff;
rom[99756] = 12'heee;
rom[99757] = 12'heee;
rom[99758] = 12'heee;
rom[99759] = 12'heee;
rom[99760] = 12'hddd;
rom[99761] = 12'hddd;
rom[99762] = 12'hddd;
rom[99763] = 12'hddd;
rom[99764] = 12'hddd;
rom[99765] = 12'hddd;
rom[99766] = 12'hddd;
rom[99767] = 12'hddd;
rom[99768] = 12'hddd;
rom[99769] = 12'hddd;
rom[99770] = 12'hddd;
rom[99771] = 12'hccc;
rom[99772] = 12'hccc;
rom[99773] = 12'hccc;
rom[99774] = 12'hccc;
rom[99775] = 12'hccc;
rom[99776] = 12'hccc;
rom[99777] = 12'hccc;
rom[99778] = 12'hccc;
rom[99779] = 12'hccc;
rom[99780] = 12'hccc;
rom[99781] = 12'hccc;
rom[99782] = 12'hccc;
rom[99783] = 12'hccc;
rom[99784] = 12'hccc;
rom[99785] = 12'hbbb;
rom[99786] = 12'hbbb;
rom[99787] = 12'hbbb;
rom[99788] = 12'hbbb;
rom[99789] = 12'hbbb;
rom[99790] = 12'hbbb;
rom[99791] = 12'hbbb;
rom[99792] = 12'hbbb;
rom[99793] = 12'hbbb;
rom[99794] = 12'hbbb;
rom[99795] = 12'hbbb;
rom[99796] = 12'hbbb;
rom[99797] = 12'hbbb;
rom[99798] = 12'hbbb;
rom[99799] = 12'hbbb;
rom[99800] = 12'hbbb;
rom[99801] = 12'hbbb;
rom[99802] = 12'hbbb;
rom[99803] = 12'hbbb;
rom[99804] = 12'hbbb;
rom[99805] = 12'hbbb;
rom[99806] = 12'hbbb;
rom[99807] = 12'hbbb;
rom[99808] = 12'hbbb;
rom[99809] = 12'hbbb;
rom[99810] = 12'hbbb;
rom[99811] = 12'hbbb;
rom[99812] = 12'hccc;
rom[99813] = 12'hccc;
rom[99814] = 12'hccc;
rom[99815] = 12'hccc;
rom[99816] = 12'hccc;
rom[99817] = 12'hccc;
rom[99818] = 12'hccc;
rom[99819] = 12'hccc;
rom[99820] = 12'hccc;
rom[99821] = 12'hccc;
rom[99822] = 12'hccc;
rom[99823] = 12'hccc;
rom[99824] = 12'hccc;
rom[99825] = 12'hccc;
rom[99826] = 12'hccc;
rom[99827] = 12'hbbb;
rom[99828] = 12'hbbb;
rom[99829] = 12'hbbb;
rom[99830] = 12'hbbb;
rom[99831] = 12'hbbb;
rom[99832] = 12'hbbb;
rom[99833] = 12'hbbb;
rom[99834] = 12'hbbb;
rom[99835] = 12'hbbb;
rom[99836] = 12'hbbb;
rom[99837] = 12'hbbb;
rom[99838] = 12'hbbb;
rom[99839] = 12'hbbb;
rom[99840] = 12'hbbb;
rom[99841] = 12'hbbb;
rom[99842] = 12'hbbb;
rom[99843] = 12'hbbb;
rom[99844] = 12'hccc;
rom[99845] = 12'hccc;
rom[99846] = 12'hccc;
rom[99847] = 12'hccc;
rom[99848] = 12'hccc;
rom[99849] = 12'hccc;
rom[99850] = 12'hccc;
rom[99851] = 12'hbbb;
rom[99852] = 12'hbbb;
rom[99853] = 12'hbbb;
rom[99854] = 12'hbbb;
rom[99855] = 12'haaa;
rom[99856] = 12'haaa;
rom[99857] = 12'haaa;
rom[99858] = 12'haaa;
rom[99859] = 12'haaa;
rom[99860] = 12'h999;
rom[99861] = 12'h999;
rom[99862] = 12'h999;
rom[99863] = 12'h999;
rom[99864] = 12'haaa;
rom[99865] = 12'haaa;
rom[99866] = 12'haaa;
rom[99867] = 12'haaa;
rom[99868] = 12'haaa;
rom[99869] = 12'haaa;
rom[99870] = 12'haaa;
rom[99871] = 12'haaa;
rom[99872] = 12'haaa;
rom[99873] = 12'haaa;
rom[99874] = 12'haaa;
rom[99875] = 12'hbbb;
rom[99876] = 12'hbbb;
rom[99877] = 12'hccc;
rom[99878] = 12'hddd;
rom[99879] = 12'heee;
rom[99880] = 12'hfff;
rom[99881] = 12'hfff;
rom[99882] = 12'hfff;
rom[99883] = 12'heee;
rom[99884] = 12'heee;
rom[99885] = 12'hddd;
rom[99886] = 12'hccc;
rom[99887] = 12'hbbb;
rom[99888] = 12'haaa;
rom[99889] = 12'haaa;
rom[99890] = 12'h999;
rom[99891] = 12'h999;
rom[99892] = 12'h888;
rom[99893] = 12'h777;
rom[99894] = 12'h666;
rom[99895] = 12'h555;
rom[99896] = 12'h444;
rom[99897] = 12'h444;
rom[99898] = 12'h333;
rom[99899] = 12'h333;
rom[99900] = 12'h333;
rom[99901] = 12'h333;
rom[99902] = 12'h333;
rom[99903] = 12'h444;
rom[99904] = 12'h666;
rom[99905] = 12'h888;
rom[99906] = 12'hbbb;
rom[99907] = 12'hddd;
rom[99908] = 12'heee;
rom[99909] = 12'heee;
rom[99910] = 12'hbbb;
rom[99911] = 12'h888;
rom[99912] = 12'h555;
rom[99913] = 12'h444;
rom[99914] = 12'h555;
rom[99915] = 12'h555;
rom[99916] = 12'h666;
rom[99917] = 12'h666;
rom[99918] = 12'h666;
rom[99919] = 12'h777;
rom[99920] = 12'h666;
rom[99921] = 12'h666;
rom[99922] = 12'h555;
rom[99923] = 12'h555;
rom[99924] = 12'h444;
rom[99925] = 12'h444;
rom[99926] = 12'h333;
rom[99927] = 12'h333;
rom[99928] = 12'h666;
rom[99929] = 12'h888;
rom[99930] = 12'haaa;
rom[99931] = 12'hddd;
rom[99932] = 12'heee;
rom[99933] = 12'hfff;
rom[99934] = 12'heee;
rom[99935] = 12'hccc;
rom[99936] = 12'h999;
rom[99937] = 12'h777;
rom[99938] = 12'h555;
rom[99939] = 12'h444;
rom[99940] = 12'h333;
rom[99941] = 12'h333;
rom[99942] = 12'h222;
rom[99943] = 12'h222;
rom[99944] = 12'h111;
rom[99945] = 12'h111;
rom[99946] = 12'h111;
rom[99947] = 12'h111;
rom[99948] = 12'h111;
rom[99949] = 12'h111;
rom[99950] = 12'h111;
rom[99951] = 12'h111;
rom[99952] = 12'h111;
rom[99953] = 12'h111;
rom[99954] = 12'h111;
rom[99955] = 12'h111;
rom[99956] = 12'h111;
rom[99957] = 12'h111;
rom[99958] = 12'h111;
rom[99959] = 12'h111;
rom[99960] = 12'h111;
rom[99961] = 12'h111;
rom[99962] = 12'h111;
rom[99963] = 12'h111;
rom[99964] = 12'h111;
rom[99965] = 12'h111;
rom[99966] = 12'h111;
rom[99967] = 12'h111;
rom[99968] = 12'h111;
rom[99969] = 12'h111;
rom[99970] = 12'h111;
rom[99971] = 12'h111;
rom[99972] = 12'h111;
rom[99973] = 12'h111;
rom[99974] = 12'h111;
rom[99975] = 12'h111;
rom[99976] = 12'h  0;
rom[99977] = 12'h  0;
rom[99978] = 12'h  0;
rom[99979] = 12'h111;
rom[99980] = 12'h111;
rom[99981] = 12'h111;
rom[99982] = 12'h111;
rom[99983] = 12'h111;
rom[99984] = 12'h222;
rom[99985] = 12'h222;
rom[99986] = 12'h333;
rom[99987] = 12'h333;
rom[99988] = 12'h444;
rom[99989] = 12'h333;
rom[99990] = 12'h222;
rom[99991] = 12'h222;
rom[99992] = 12'h111;
rom[99993] = 12'h111;
rom[99994] = 12'h111;
rom[99995] = 12'h111;
rom[99996] = 12'h222;
rom[99997] = 12'h222;
rom[99998] = 12'h222;
rom[99999] = 12'h222;
rom[100000] = 12'hfff;
rom[100001] = 12'hfff;
rom[100002] = 12'hfff;
rom[100003] = 12'hfff;
rom[100004] = 12'hfff;
rom[100005] = 12'hfff;
rom[100006] = 12'hfff;
rom[100007] = 12'hfff;
rom[100008] = 12'hfff;
rom[100009] = 12'hfff;
rom[100010] = 12'hfff;
rom[100011] = 12'hfff;
rom[100012] = 12'hfff;
rom[100013] = 12'hfff;
rom[100014] = 12'hfff;
rom[100015] = 12'hfff;
rom[100016] = 12'hfff;
rom[100017] = 12'hfff;
rom[100018] = 12'hfff;
rom[100019] = 12'hfff;
rom[100020] = 12'hfff;
rom[100021] = 12'hfff;
rom[100022] = 12'hfff;
rom[100023] = 12'hfff;
rom[100024] = 12'hfff;
rom[100025] = 12'hfff;
rom[100026] = 12'hfff;
rom[100027] = 12'hfff;
rom[100028] = 12'hfff;
rom[100029] = 12'hfff;
rom[100030] = 12'hfff;
rom[100031] = 12'hfff;
rom[100032] = 12'hfff;
rom[100033] = 12'hfff;
rom[100034] = 12'hfff;
rom[100035] = 12'hfff;
rom[100036] = 12'hfff;
rom[100037] = 12'hfff;
rom[100038] = 12'hfff;
rom[100039] = 12'hfff;
rom[100040] = 12'hfff;
rom[100041] = 12'hfff;
rom[100042] = 12'hfff;
rom[100043] = 12'hfff;
rom[100044] = 12'hfff;
rom[100045] = 12'hfff;
rom[100046] = 12'hfff;
rom[100047] = 12'hfff;
rom[100048] = 12'hfff;
rom[100049] = 12'hfff;
rom[100050] = 12'hfff;
rom[100051] = 12'hfff;
rom[100052] = 12'hfff;
rom[100053] = 12'hfff;
rom[100054] = 12'hfff;
rom[100055] = 12'hfff;
rom[100056] = 12'hfff;
rom[100057] = 12'hfff;
rom[100058] = 12'hfff;
rom[100059] = 12'hfff;
rom[100060] = 12'hfff;
rom[100061] = 12'hfff;
rom[100062] = 12'hfff;
rom[100063] = 12'hfff;
rom[100064] = 12'hfff;
rom[100065] = 12'hfff;
rom[100066] = 12'hfff;
rom[100067] = 12'hfff;
rom[100068] = 12'hfff;
rom[100069] = 12'hfff;
rom[100070] = 12'hfff;
rom[100071] = 12'hfff;
rom[100072] = 12'hfff;
rom[100073] = 12'hfff;
rom[100074] = 12'hfff;
rom[100075] = 12'hfff;
rom[100076] = 12'hfff;
rom[100077] = 12'hfff;
rom[100078] = 12'hfff;
rom[100079] = 12'hfff;
rom[100080] = 12'hfff;
rom[100081] = 12'hfff;
rom[100082] = 12'heee;
rom[100083] = 12'heee;
rom[100084] = 12'hfff;
rom[100085] = 12'hfff;
rom[100086] = 12'hfff;
rom[100087] = 12'hfff;
rom[100088] = 12'hfff;
rom[100089] = 12'hfff;
rom[100090] = 12'hfff;
rom[100091] = 12'hfff;
rom[100092] = 12'hfff;
rom[100093] = 12'hfff;
rom[100094] = 12'hfff;
rom[100095] = 12'hfff;
rom[100096] = 12'hfff;
rom[100097] = 12'hfff;
rom[100098] = 12'hfff;
rom[100099] = 12'hfff;
rom[100100] = 12'hfff;
rom[100101] = 12'hfff;
rom[100102] = 12'heee;
rom[100103] = 12'heee;
rom[100104] = 12'hfff;
rom[100105] = 12'hfff;
rom[100106] = 12'hfff;
rom[100107] = 12'hfff;
rom[100108] = 12'hfff;
rom[100109] = 12'hfff;
rom[100110] = 12'hfff;
rom[100111] = 12'hfff;
rom[100112] = 12'hfff;
rom[100113] = 12'hfff;
rom[100114] = 12'hfff;
rom[100115] = 12'hfff;
rom[100116] = 12'hfff;
rom[100117] = 12'hfff;
rom[100118] = 12'hfff;
rom[100119] = 12'hfff;
rom[100120] = 12'hfff;
rom[100121] = 12'hfff;
rom[100122] = 12'hfff;
rom[100123] = 12'hfff;
rom[100124] = 12'hfff;
rom[100125] = 12'hfff;
rom[100126] = 12'hfff;
rom[100127] = 12'hfff;
rom[100128] = 12'hfff;
rom[100129] = 12'hfff;
rom[100130] = 12'hfff;
rom[100131] = 12'hfff;
rom[100132] = 12'hfff;
rom[100133] = 12'hfff;
rom[100134] = 12'hfff;
rom[100135] = 12'hfff;
rom[100136] = 12'hfff;
rom[100137] = 12'hfff;
rom[100138] = 12'hfff;
rom[100139] = 12'hfff;
rom[100140] = 12'hfff;
rom[100141] = 12'hfff;
rom[100142] = 12'hfff;
rom[100143] = 12'hfff;
rom[100144] = 12'hfff;
rom[100145] = 12'hfff;
rom[100146] = 12'hfff;
rom[100147] = 12'hfff;
rom[100148] = 12'hfff;
rom[100149] = 12'hfff;
rom[100150] = 12'hfff;
rom[100151] = 12'hfff;
rom[100152] = 12'hfff;
rom[100153] = 12'hfff;
rom[100154] = 12'hfff;
rom[100155] = 12'hfff;
rom[100156] = 12'hfff;
rom[100157] = 12'hfff;
rom[100158] = 12'hfff;
rom[100159] = 12'hfff;
rom[100160] = 12'heee;
rom[100161] = 12'heee;
rom[100162] = 12'heee;
rom[100163] = 12'hddd;
rom[100164] = 12'hddd;
rom[100165] = 12'hddd;
rom[100166] = 12'hddd;
rom[100167] = 12'hddd;
rom[100168] = 12'hddd;
rom[100169] = 12'hddd;
rom[100170] = 12'hddd;
rom[100171] = 12'hddd;
rom[100172] = 12'hddd;
rom[100173] = 12'hccc;
rom[100174] = 12'hddd;
rom[100175] = 12'hddd;
rom[100176] = 12'hccc;
rom[100177] = 12'hccc;
rom[100178] = 12'hccc;
rom[100179] = 12'hccc;
rom[100180] = 12'hccc;
rom[100181] = 12'hccc;
rom[100182] = 12'hccc;
rom[100183] = 12'hccc;
rom[100184] = 12'hccc;
rom[100185] = 12'hccc;
rom[100186] = 12'hccc;
rom[100187] = 12'hccc;
rom[100188] = 12'hccc;
rom[100189] = 12'hbbb;
rom[100190] = 12'hbbb;
rom[100191] = 12'hbbb;
rom[100192] = 12'hbbb;
rom[100193] = 12'hbbb;
rom[100194] = 12'hbbb;
rom[100195] = 12'hbbb;
rom[100196] = 12'hbbb;
rom[100197] = 12'hbbb;
rom[100198] = 12'hbbb;
rom[100199] = 12'hbbb;
rom[100200] = 12'hbbb;
rom[100201] = 12'hbbb;
rom[100202] = 12'hbbb;
rom[100203] = 12'hccc;
rom[100204] = 12'hccc;
rom[100205] = 12'hccc;
rom[100206] = 12'hccc;
rom[100207] = 12'hccc;
rom[100208] = 12'hccc;
rom[100209] = 12'hccc;
rom[100210] = 12'hccc;
rom[100211] = 12'hccc;
rom[100212] = 12'hccc;
rom[100213] = 12'hccc;
rom[100214] = 12'hccc;
rom[100215] = 12'hccc;
rom[100216] = 12'hccc;
rom[100217] = 12'hccc;
rom[100218] = 12'hccc;
rom[100219] = 12'hddd;
rom[100220] = 12'hddd;
rom[100221] = 12'hddd;
rom[100222] = 12'hddd;
rom[100223] = 12'hddd;
rom[100224] = 12'hddd;
rom[100225] = 12'hddd;
rom[100226] = 12'hddd;
rom[100227] = 12'hccc;
rom[100228] = 12'hccc;
rom[100229] = 12'hccc;
rom[100230] = 12'hccc;
rom[100231] = 12'hccc;
rom[100232] = 12'hccc;
rom[100233] = 12'hccc;
rom[100234] = 12'hccc;
rom[100235] = 12'hccc;
rom[100236] = 12'hccc;
rom[100237] = 12'hccc;
rom[100238] = 12'hccc;
rom[100239] = 12'hccc;
rom[100240] = 12'hccc;
rom[100241] = 12'hccc;
rom[100242] = 12'hccc;
rom[100243] = 12'hccc;
rom[100244] = 12'hddd;
rom[100245] = 12'hddd;
rom[100246] = 12'hddd;
rom[100247] = 12'hccc;
rom[100248] = 12'hddd;
rom[100249] = 12'hccc;
rom[100250] = 12'hccc;
rom[100251] = 12'hccc;
rom[100252] = 12'hccc;
rom[100253] = 12'hbbb;
rom[100254] = 12'hbbb;
rom[100255] = 12'haaa;
rom[100256] = 12'haaa;
rom[100257] = 12'haaa;
rom[100258] = 12'haaa;
rom[100259] = 12'haaa;
rom[100260] = 12'haaa;
rom[100261] = 12'haaa;
rom[100262] = 12'haaa;
rom[100263] = 12'haaa;
rom[100264] = 12'haaa;
rom[100265] = 12'haaa;
rom[100266] = 12'haaa;
rom[100267] = 12'haaa;
rom[100268] = 12'haaa;
rom[100269] = 12'haaa;
rom[100270] = 12'haaa;
rom[100271] = 12'haaa;
rom[100272] = 12'haaa;
rom[100273] = 12'hbbb;
rom[100274] = 12'hbbb;
rom[100275] = 12'hccc;
rom[100276] = 12'hddd;
rom[100277] = 12'hddd;
rom[100278] = 12'heee;
rom[100279] = 12'hfff;
rom[100280] = 12'hfff;
rom[100281] = 12'hfff;
rom[100282] = 12'heee;
rom[100283] = 12'hddd;
rom[100284] = 12'hccc;
rom[100285] = 12'hccc;
rom[100286] = 12'hbbb;
rom[100287] = 12'hbbb;
rom[100288] = 12'hbbb;
rom[100289] = 12'haaa;
rom[100290] = 12'h999;
rom[100291] = 12'h999;
rom[100292] = 12'h888;
rom[100293] = 12'h888;
rom[100294] = 12'h666;
rom[100295] = 12'h555;
rom[100296] = 12'h444;
rom[100297] = 12'h444;
rom[100298] = 12'h444;
rom[100299] = 12'h333;
rom[100300] = 12'h333;
rom[100301] = 12'h333;
rom[100302] = 12'h222;
rom[100303] = 12'h222;
rom[100304] = 12'h222;
rom[100305] = 12'h444;
rom[100306] = 12'h666;
rom[100307] = 12'h999;
rom[100308] = 12'hddd;
rom[100309] = 12'hfff;
rom[100310] = 12'heee;
rom[100311] = 12'hccc;
rom[100312] = 12'h888;
rom[100313] = 12'h666;
rom[100314] = 12'h444;
rom[100315] = 12'h444;
rom[100316] = 12'h555;
rom[100317] = 12'h666;
rom[100318] = 12'h666;
rom[100319] = 12'h666;
rom[100320] = 12'h777;
rom[100321] = 12'h666;
rom[100322] = 12'h555;
rom[100323] = 12'h444;
rom[100324] = 12'h444;
rom[100325] = 12'h444;
rom[100326] = 12'h333;
rom[100327] = 12'h333;
rom[100328] = 12'h333;
rom[100329] = 12'h444;
rom[100330] = 12'h666;
rom[100331] = 12'h999;
rom[100332] = 12'hbbb;
rom[100333] = 12'heee;
rom[100334] = 12'hfff;
rom[100335] = 12'hfff;
rom[100336] = 12'hddd;
rom[100337] = 12'hbbb;
rom[100338] = 12'h888;
rom[100339] = 12'h555;
rom[100340] = 12'h444;
rom[100341] = 12'h333;
rom[100342] = 12'h333;
rom[100343] = 12'h222;
rom[100344] = 12'h222;
rom[100345] = 12'h222;
rom[100346] = 12'h222;
rom[100347] = 12'h111;
rom[100348] = 12'h111;
rom[100349] = 12'h111;
rom[100350] = 12'h111;
rom[100351] = 12'h111;
rom[100352] = 12'h111;
rom[100353] = 12'h111;
rom[100354] = 12'h111;
rom[100355] = 12'h111;
rom[100356] = 12'h111;
rom[100357] = 12'h111;
rom[100358] = 12'h111;
rom[100359] = 12'h111;
rom[100360] = 12'h111;
rom[100361] = 12'h111;
rom[100362] = 12'h111;
rom[100363] = 12'h111;
rom[100364] = 12'h111;
rom[100365] = 12'h111;
rom[100366] = 12'h111;
rom[100367] = 12'h111;
rom[100368] = 12'h  0;
rom[100369] = 12'h  0;
rom[100370] = 12'h  0;
rom[100371] = 12'h  0;
rom[100372] = 12'h  0;
rom[100373] = 12'h  0;
rom[100374] = 12'h  0;
rom[100375] = 12'h  0;
rom[100376] = 12'h  0;
rom[100377] = 12'h  0;
rom[100378] = 12'h  0;
rom[100379] = 12'h  0;
rom[100380] = 12'h111;
rom[100381] = 12'h111;
rom[100382] = 12'h111;
rom[100383] = 12'h111;
rom[100384] = 12'h111;
rom[100385] = 12'h111;
rom[100386] = 12'h222;
rom[100387] = 12'h333;
rom[100388] = 12'h333;
rom[100389] = 12'h333;
rom[100390] = 12'h333;
rom[100391] = 12'h222;
rom[100392] = 12'h111;
rom[100393] = 12'h111;
rom[100394] = 12'h111;
rom[100395] = 12'h111;
rom[100396] = 12'h111;
rom[100397] = 12'h111;
rom[100398] = 12'h111;
rom[100399] = 12'h111;
rom[100400] = 12'hfff;
rom[100401] = 12'hfff;
rom[100402] = 12'hfff;
rom[100403] = 12'hfff;
rom[100404] = 12'hfff;
rom[100405] = 12'hfff;
rom[100406] = 12'hfff;
rom[100407] = 12'hfff;
rom[100408] = 12'hfff;
rom[100409] = 12'hfff;
rom[100410] = 12'hfff;
rom[100411] = 12'hfff;
rom[100412] = 12'hfff;
rom[100413] = 12'hfff;
rom[100414] = 12'hfff;
rom[100415] = 12'hfff;
rom[100416] = 12'hfff;
rom[100417] = 12'hfff;
rom[100418] = 12'hfff;
rom[100419] = 12'hfff;
rom[100420] = 12'hfff;
rom[100421] = 12'hfff;
rom[100422] = 12'hfff;
rom[100423] = 12'hfff;
rom[100424] = 12'hfff;
rom[100425] = 12'hfff;
rom[100426] = 12'hfff;
rom[100427] = 12'hfff;
rom[100428] = 12'hfff;
rom[100429] = 12'hfff;
rom[100430] = 12'hfff;
rom[100431] = 12'hfff;
rom[100432] = 12'hfff;
rom[100433] = 12'hfff;
rom[100434] = 12'hfff;
rom[100435] = 12'hfff;
rom[100436] = 12'hfff;
rom[100437] = 12'hfff;
rom[100438] = 12'hfff;
rom[100439] = 12'hfff;
rom[100440] = 12'hfff;
rom[100441] = 12'hfff;
rom[100442] = 12'hfff;
rom[100443] = 12'hfff;
rom[100444] = 12'hfff;
rom[100445] = 12'hfff;
rom[100446] = 12'hfff;
rom[100447] = 12'hfff;
rom[100448] = 12'hfff;
rom[100449] = 12'hfff;
rom[100450] = 12'hfff;
rom[100451] = 12'hfff;
rom[100452] = 12'hfff;
rom[100453] = 12'hfff;
rom[100454] = 12'hfff;
rom[100455] = 12'hfff;
rom[100456] = 12'hfff;
rom[100457] = 12'hfff;
rom[100458] = 12'hfff;
rom[100459] = 12'hfff;
rom[100460] = 12'hfff;
rom[100461] = 12'hfff;
rom[100462] = 12'hfff;
rom[100463] = 12'hfff;
rom[100464] = 12'hfff;
rom[100465] = 12'hfff;
rom[100466] = 12'hfff;
rom[100467] = 12'hfff;
rom[100468] = 12'hfff;
rom[100469] = 12'hfff;
rom[100470] = 12'hfff;
rom[100471] = 12'hfff;
rom[100472] = 12'hfff;
rom[100473] = 12'hfff;
rom[100474] = 12'hfff;
rom[100475] = 12'hfff;
rom[100476] = 12'hfff;
rom[100477] = 12'hfff;
rom[100478] = 12'hfff;
rom[100479] = 12'hfff;
rom[100480] = 12'heee;
rom[100481] = 12'heee;
rom[100482] = 12'heee;
rom[100483] = 12'heee;
rom[100484] = 12'hfff;
rom[100485] = 12'hfff;
rom[100486] = 12'hfff;
rom[100487] = 12'heee;
rom[100488] = 12'hfff;
rom[100489] = 12'hfff;
rom[100490] = 12'hfff;
rom[100491] = 12'hfff;
rom[100492] = 12'hfff;
rom[100493] = 12'hfff;
rom[100494] = 12'hfff;
rom[100495] = 12'hfff;
rom[100496] = 12'hfff;
rom[100497] = 12'hfff;
rom[100498] = 12'hfff;
rom[100499] = 12'hfff;
rom[100500] = 12'heee;
rom[100501] = 12'heee;
rom[100502] = 12'heee;
rom[100503] = 12'heee;
rom[100504] = 12'heee;
rom[100505] = 12'heee;
rom[100506] = 12'hfff;
rom[100507] = 12'hfff;
rom[100508] = 12'hfff;
rom[100509] = 12'hfff;
rom[100510] = 12'hfff;
rom[100511] = 12'hfff;
rom[100512] = 12'hfff;
rom[100513] = 12'hfff;
rom[100514] = 12'hfff;
rom[100515] = 12'hfff;
rom[100516] = 12'hfff;
rom[100517] = 12'hfff;
rom[100518] = 12'hfff;
rom[100519] = 12'hfff;
rom[100520] = 12'hfff;
rom[100521] = 12'hfff;
rom[100522] = 12'hfff;
rom[100523] = 12'hfff;
rom[100524] = 12'hfff;
rom[100525] = 12'hfff;
rom[100526] = 12'hfff;
rom[100527] = 12'hfff;
rom[100528] = 12'hfff;
rom[100529] = 12'hfff;
rom[100530] = 12'hfff;
rom[100531] = 12'hfff;
rom[100532] = 12'hfff;
rom[100533] = 12'hfff;
rom[100534] = 12'hfff;
rom[100535] = 12'hfff;
rom[100536] = 12'hfff;
rom[100537] = 12'hfff;
rom[100538] = 12'hfff;
rom[100539] = 12'hfff;
rom[100540] = 12'hfff;
rom[100541] = 12'hfff;
rom[100542] = 12'hfff;
rom[100543] = 12'hfff;
rom[100544] = 12'hfff;
rom[100545] = 12'hfff;
rom[100546] = 12'hfff;
rom[100547] = 12'hfff;
rom[100548] = 12'hfff;
rom[100549] = 12'hfff;
rom[100550] = 12'hfff;
rom[100551] = 12'hfff;
rom[100552] = 12'hfff;
rom[100553] = 12'hfff;
rom[100554] = 12'hfff;
rom[100555] = 12'hfff;
rom[100556] = 12'hfff;
rom[100557] = 12'hfff;
rom[100558] = 12'hfff;
rom[100559] = 12'hfff;
rom[100560] = 12'hfff;
rom[100561] = 12'hfff;
rom[100562] = 12'heee;
rom[100563] = 12'heee;
rom[100564] = 12'heee;
rom[100565] = 12'heee;
rom[100566] = 12'heee;
rom[100567] = 12'heee;
rom[100568] = 12'hddd;
rom[100569] = 12'hddd;
rom[100570] = 12'hddd;
rom[100571] = 12'hddd;
rom[100572] = 12'hddd;
rom[100573] = 12'hddd;
rom[100574] = 12'hddd;
rom[100575] = 12'hddd;
rom[100576] = 12'hddd;
rom[100577] = 12'hccc;
rom[100578] = 12'hccc;
rom[100579] = 12'hccc;
rom[100580] = 12'hccc;
rom[100581] = 12'hccc;
rom[100582] = 12'hccc;
rom[100583] = 12'hccc;
rom[100584] = 12'hccc;
rom[100585] = 12'hccc;
rom[100586] = 12'hccc;
rom[100587] = 12'hccc;
rom[100588] = 12'hccc;
rom[100589] = 12'hccc;
rom[100590] = 12'hccc;
rom[100591] = 12'hccc;
rom[100592] = 12'hccc;
rom[100593] = 12'hccc;
rom[100594] = 12'hccc;
rom[100595] = 12'hccc;
rom[100596] = 12'hccc;
rom[100597] = 12'hccc;
rom[100598] = 12'hccc;
rom[100599] = 12'hccc;
rom[100600] = 12'hccc;
rom[100601] = 12'hccc;
rom[100602] = 12'hccc;
rom[100603] = 12'hccc;
rom[100604] = 12'hccc;
rom[100605] = 12'hccc;
rom[100606] = 12'hccc;
rom[100607] = 12'hccc;
rom[100608] = 12'hccc;
rom[100609] = 12'hccc;
rom[100610] = 12'hccc;
rom[100611] = 12'hccc;
rom[100612] = 12'hccc;
rom[100613] = 12'hccc;
rom[100614] = 12'hddd;
rom[100615] = 12'hddd;
rom[100616] = 12'hccc;
rom[100617] = 12'hddd;
rom[100618] = 12'hddd;
rom[100619] = 12'hddd;
rom[100620] = 12'hddd;
rom[100621] = 12'hddd;
rom[100622] = 12'hddd;
rom[100623] = 12'hddd;
rom[100624] = 12'hddd;
rom[100625] = 12'hddd;
rom[100626] = 12'hddd;
rom[100627] = 12'hddd;
rom[100628] = 12'hddd;
rom[100629] = 12'hddd;
rom[100630] = 12'hddd;
rom[100631] = 12'hddd;
rom[100632] = 12'hddd;
rom[100633] = 12'hddd;
rom[100634] = 12'hddd;
rom[100635] = 12'hddd;
rom[100636] = 12'hddd;
rom[100637] = 12'hddd;
rom[100638] = 12'hddd;
rom[100639] = 12'hddd;
rom[100640] = 12'hddd;
rom[100641] = 12'hddd;
rom[100642] = 12'hddd;
rom[100643] = 12'hddd;
rom[100644] = 12'hddd;
rom[100645] = 12'hddd;
rom[100646] = 12'hddd;
rom[100647] = 12'hccc;
rom[100648] = 12'hccc;
rom[100649] = 12'hccc;
rom[100650] = 12'hccc;
rom[100651] = 12'hccc;
rom[100652] = 12'hccc;
rom[100653] = 12'hbbb;
rom[100654] = 12'hbbb;
rom[100655] = 12'hbbb;
rom[100656] = 12'haaa;
rom[100657] = 12'haaa;
rom[100658] = 12'haaa;
rom[100659] = 12'haaa;
rom[100660] = 12'haaa;
rom[100661] = 12'haaa;
rom[100662] = 12'haaa;
rom[100663] = 12'haaa;
rom[100664] = 12'haaa;
rom[100665] = 12'haaa;
rom[100666] = 12'haaa;
rom[100667] = 12'haaa;
rom[100668] = 12'haaa;
rom[100669] = 12'haaa;
rom[100670] = 12'hbbb;
rom[100671] = 12'hbbb;
rom[100672] = 12'hccc;
rom[100673] = 12'hccc;
rom[100674] = 12'hddd;
rom[100675] = 12'hddd;
rom[100676] = 12'heee;
rom[100677] = 12'hfff;
rom[100678] = 12'hfff;
rom[100679] = 12'hfff;
rom[100680] = 12'hfff;
rom[100681] = 12'heee;
rom[100682] = 12'hddd;
rom[100683] = 12'hddd;
rom[100684] = 12'hccc;
rom[100685] = 12'hccc;
rom[100686] = 12'hccc;
rom[100687] = 12'hccc;
rom[100688] = 12'hbbb;
rom[100689] = 12'haaa;
rom[100690] = 12'h999;
rom[100691] = 12'h999;
rom[100692] = 12'h999;
rom[100693] = 12'h888;
rom[100694] = 12'h777;
rom[100695] = 12'h666;
rom[100696] = 12'h555;
rom[100697] = 12'h555;
rom[100698] = 12'h444;
rom[100699] = 12'h333;
rom[100700] = 12'h333;
rom[100701] = 12'h333;
rom[100702] = 12'h333;
rom[100703] = 12'h333;
rom[100704] = 12'h333;
rom[100705] = 12'h333;
rom[100706] = 12'h444;
rom[100707] = 12'h555;
rom[100708] = 12'h777;
rom[100709] = 12'haaa;
rom[100710] = 12'hccc;
rom[100711] = 12'heee;
rom[100712] = 12'hddd;
rom[100713] = 12'haaa;
rom[100714] = 12'h666;
rom[100715] = 12'h444;
rom[100716] = 12'h444;
rom[100717] = 12'h555;
rom[100718] = 12'h666;
rom[100719] = 12'h666;
rom[100720] = 12'h888;
rom[100721] = 12'h666;
rom[100722] = 12'h555;
rom[100723] = 12'h444;
rom[100724] = 12'h333;
rom[100725] = 12'h444;
rom[100726] = 12'h444;
rom[100727] = 12'h444;
rom[100728] = 12'h333;
rom[100729] = 12'h333;
rom[100730] = 12'h444;
rom[100731] = 12'h555;
rom[100732] = 12'h777;
rom[100733] = 12'h999;
rom[100734] = 12'hccc;
rom[100735] = 12'hfff;
rom[100736] = 12'hfff;
rom[100737] = 12'heee;
rom[100738] = 12'hccc;
rom[100739] = 12'h999;
rom[100740] = 12'h666;
rom[100741] = 12'h555;
rom[100742] = 12'h444;
rom[100743] = 12'h333;
rom[100744] = 12'h222;
rom[100745] = 12'h222;
rom[100746] = 12'h222;
rom[100747] = 12'h222;
rom[100748] = 12'h222;
rom[100749] = 12'h111;
rom[100750] = 12'h111;
rom[100751] = 12'h111;
rom[100752] = 12'h111;
rom[100753] = 12'h111;
rom[100754] = 12'h111;
rom[100755] = 12'h111;
rom[100756] = 12'h111;
rom[100757] = 12'h111;
rom[100758] = 12'h111;
rom[100759] = 12'h111;
rom[100760] = 12'h111;
rom[100761] = 12'h111;
rom[100762] = 12'h111;
rom[100763] = 12'h111;
rom[100764] = 12'h111;
rom[100765] = 12'h  0;
rom[100766] = 12'h  0;
rom[100767] = 12'h111;
rom[100768] = 12'h  0;
rom[100769] = 12'h  0;
rom[100770] = 12'h  0;
rom[100771] = 12'h  0;
rom[100772] = 12'h  0;
rom[100773] = 12'h  0;
rom[100774] = 12'h  0;
rom[100775] = 12'h  0;
rom[100776] = 12'h  0;
rom[100777] = 12'h  0;
rom[100778] = 12'h  0;
rom[100779] = 12'h  0;
rom[100780] = 12'h  0;
rom[100781] = 12'h111;
rom[100782] = 12'h111;
rom[100783] = 12'h111;
rom[100784] = 12'h111;
rom[100785] = 12'h111;
rom[100786] = 12'h111;
rom[100787] = 12'h222;
rom[100788] = 12'h333;
rom[100789] = 12'h333;
rom[100790] = 12'h333;
rom[100791] = 12'h222;
rom[100792] = 12'h111;
rom[100793] = 12'h111;
rom[100794] = 12'h111;
rom[100795] = 12'h111;
rom[100796] = 12'h111;
rom[100797] = 12'h111;
rom[100798] = 12'h111;
rom[100799] = 12'h111;
rom[100800] = 12'hfff;
rom[100801] = 12'hfff;
rom[100802] = 12'hfff;
rom[100803] = 12'hfff;
rom[100804] = 12'hfff;
rom[100805] = 12'hfff;
rom[100806] = 12'hfff;
rom[100807] = 12'hfff;
rom[100808] = 12'hfff;
rom[100809] = 12'hfff;
rom[100810] = 12'hfff;
rom[100811] = 12'hfff;
rom[100812] = 12'hfff;
rom[100813] = 12'hfff;
rom[100814] = 12'hfff;
rom[100815] = 12'hfff;
rom[100816] = 12'hfff;
rom[100817] = 12'hfff;
rom[100818] = 12'hfff;
rom[100819] = 12'hfff;
rom[100820] = 12'hfff;
rom[100821] = 12'hfff;
rom[100822] = 12'hfff;
rom[100823] = 12'hfff;
rom[100824] = 12'hfff;
rom[100825] = 12'hfff;
rom[100826] = 12'hfff;
rom[100827] = 12'hfff;
rom[100828] = 12'hfff;
rom[100829] = 12'hfff;
rom[100830] = 12'hfff;
rom[100831] = 12'hfff;
rom[100832] = 12'hfff;
rom[100833] = 12'hfff;
rom[100834] = 12'hfff;
rom[100835] = 12'hfff;
rom[100836] = 12'hfff;
rom[100837] = 12'hfff;
rom[100838] = 12'hfff;
rom[100839] = 12'hfff;
rom[100840] = 12'hfff;
rom[100841] = 12'hfff;
rom[100842] = 12'hfff;
rom[100843] = 12'hfff;
rom[100844] = 12'hfff;
rom[100845] = 12'hfff;
rom[100846] = 12'hfff;
rom[100847] = 12'hfff;
rom[100848] = 12'hfff;
rom[100849] = 12'hfff;
rom[100850] = 12'hfff;
rom[100851] = 12'hfff;
rom[100852] = 12'hfff;
rom[100853] = 12'hfff;
rom[100854] = 12'hfff;
rom[100855] = 12'hfff;
rom[100856] = 12'hfff;
rom[100857] = 12'hfff;
rom[100858] = 12'hfff;
rom[100859] = 12'hfff;
rom[100860] = 12'hfff;
rom[100861] = 12'hfff;
rom[100862] = 12'hfff;
rom[100863] = 12'hfff;
rom[100864] = 12'hfff;
rom[100865] = 12'hfff;
rom[100866] = 12'hfff;
rom[100867] = 12'hfff;
rom[100868] = 12'hfff;
rom[100869] = 12'hfff;
rom[100870] = 12'hfff;
rom[100871] = 12'hfff;
rom[100872] = 12'heee;
rom[100873] = 12'hfff;
rom[100874] = 12'hfff;
rom[100875] = 12'hfff;
rom[100876] = 12'hfff;
rom[100877] = 12'hfff;
rom[100878] = 12'hfff;
rom[100879] = 12'heee;
rom[100880] = 12'heee;
rom[100881] = 12'heee;
rom[100882] = 12'heee;
rom[100883] = 12'heee;
rom[100884] = 12'heee;
rom[100885] = 12'heee;
rom[100886] = 12'heee;
rom[100887] = 12'heee;
rom[100888] = 12'hfff;
rom[100889] = 12'hfff;
rom[100890] = 12'hfff;
rom[100891] = 12'hfff;
rom[100892] = 12'hfff;
rom[100893] = 12'hfff;
rom[100894] = 12'hfff;
rom[100895] = 12'hfff;
rom[100896] = 12'heee;
rom[100897] = 12'heee;
rom[100898] = 12'heee;
rom[100899] = 12'heee;
rom[100900] = 12'heee;
rom[100901] = 12'heee;
rom[100902] = 12'heee;
rom[100903] = 12'heee;
rom[100904] = 12'heee;
rom[100905] = 12'heee;
rom[100906] = 12'hfff;
rom[100907] = 12'hfff;
rom[100908] = 12'hfff;
rom[100909] = 12'hfff;
rom[100910] = 12'hfff;
rom[100911] = 12'hfff;
rom[100912] = 12'hfff;
rom[100913] = 12'hfff;
rom[100914] = 12'hfff;
rom[100915] = 12'hfff;
rom[100916] = 12'hfff;
rom[100917] = 12'hfff;
rom[100918] = 12'hfff;
rom[100919] = 12'hfff;
rom[100920] = 12'hfff;
rom[100921] = 12'hfff;
rom[100922] = 12'hfff;
rom[100923] = 12'hfff;
rom[100924] = 12'hfff;
rom[100925] = 12'hfff;
rom[100926] = 12'hfff;
rom[100927] = 12'hfff;
rom[100928] = 12'hfff;
rom[100929] = 12'hfff;
rom[100930] = 12'hfff;
rom[100931] = 12'hfff;
rom[100932] = 12'hfff;
rom[100933] = 12'hfff;
rom[100934] = 12'hfff;
rom[100935] = 12'hfff;
rom[100936] = 12'hfff;
rom[100937] = 12'hfff;
rom[100938] = 12'hfff;
rom[100939] = 12'hfff;
rom[100940] = 12'hfff;
rom[100941] = 12'hfff;
rom[100942] = 12'hfff;
rom[100943] = 12'hfff;
rom[100944] = 12'hfff;
rom[100945] = 12'hfff;
rom[100946] = 12'hfff;
rom[100947] = 12'hfff;
rom[100948] = 12'hfff;
rom[100949] = 12'hfff;
rom[100950] = 12'hfff;
rom[100951] = 12'hfff;
rom[100952] = 12'hfff;
rom[100953] = 12'hfff;
rom[100954] = 12'hfff;
rom[100955] = 12'hfff;
rom[100956] = 12'hfff;
rom[100957] = 12'hfff;
rom[100958] = 12'hfff;
rom[100959] = 12'hfff;
rom[100960] = 12'hfff;
rom[100961] = 12'hfff;
rom[100962] = 12'hfff;
rom[100963] = 12'hfff;
rom[100964] = 12'heee;
rom[100965] = 12'heee;
rom[100966] = 12'heee;
rom[100967] = 12'heee;
rom[100968] = 12'heee;
rom[100969] = 12'heee;
rom[100970] = 12'heee;
rom[100971] = 12'hddd;
rom[100972] = 12'hddd;
rom[100973] = 12'hddd;
rom[100974] = 12'hddd;
rom[100975] = 12'hddd;
rom[100976] = 12'hddd;
rom[100977] = 12'hddd;
rom[100978] = 12'hddd;
rom[100979] = 12'hccc;
rom[100980] = 12'hccc;
rom[100981] = 12'hccc;
rom[100982] = 12'hccc;
rom[100983] = 12'hccc;
rom[100984] = 12'hccc;
rom[100985] = 12'hccc;
rom[100986] = 12'hccc;
rom[100987] = 12'hccc;
rom[100988] = 12'hccc;
rom[100989] = 12'hccc;
rom[100990] = 12'hccc;
rom[100991] = 12'hccc;
rom[100992] = 12'hccc;
rom[100993] = 12'hccc;
rom[100994] = 12'hccc;
rom[100995] = 12'hccc;
rom[100996] = 12'hccc;
rom[100997] = 12'hccc;
rom[100998] = 12'hccc;
rom[100999] = 12'hccc;
rom[101000] = 12'hccc;
rom[101001] = 12'hccc;
rom[101002] = 12'hccc;
rom[101003] = 12'hccc;
rom[101004] = 12'hccc;
rom[101005] = 12'hccc;
rom[101006] = 12'hccc;
rom[101007] = 12'hccc;
rom[101008] = 12'hccc;
rom[101009] = 12'hccc;
rom[101010] = 12'hccc;
rom[101011] = 12'hccc;
rom[101012] = 12'hddd;
rom[101013] = 12'hddd;
rom[101014] = 12'hddd;
rom[101015] = 12'hddd;
rom[101016] = 12'hddd;
rom[101017] = 12'hddd;
rom[101018] = 12'hddd;
rom[101019] = 12'hddd;
rom[101020] = 12'hddd;
rom[101021] = 12'hddd;
rom[101022] = 12'heee;
rom[101023] = 12'heee;
rom[101024] = 12'hddd;
rom[101025] = 12'hddd;
rom[101026] = 12'hddd;
rom[101027] = 12'hddd;
rom[101028] = 12'hddd;
rom[101029] = 12'heee;
rom[101030] = 12'heee;
rom[101031] = 12'heee;
rom[101032] = 12'heee;
rom[101033] = 12'heee;
rom[101034] = 12'heee;
rom[101035] = 12'hddd;
rom[101036] = 12'hddd;
rom[101037] = 12'hddd;
rom[101038] = 12'hddd;
rom[101039] = 12'hddd;
rom[101040] = 12'heee;
rom[101041] = 12'hddd;
rom[101042] = 12'hddd;
rom[101043] = 12'hddd;
rom[101044] = 12'hddd;
rom[101045] = 12'hddd;
rom[101046] = 12'hddd;
rom[101047] = 12'hccc;
rom[101048] = 12'hccc;
rom[101049] = 12'hccc;
rom[101050] = 12'hccc;
rom[101051] = 12'hccc;
rom[101052] = 12'hccc;
rom[101053] = 12'hbbb;
rom[101054] = 12'hbbb;
rom[101055] = 12'hbbb;
rom[101056] = 12'haaa;
rom[101057] = 12'haaa;
rom[101058] = 12'haaa;
rom[101059] = 12'haaa;
rom[101060] = 12'haaa;
rom[101061] = 12'haaa;
rom[101062] = 12'haaa;
rom[101063] = 12'haaa;
rom[101064] = 12'haaa;
rom[101065] = 12'haaa;
rom[101066] = 12'haaa;
rom[101067] = 12'haaa;
rom[101068] = 12'haaa;
rom[101069] = 12'hbbb;
rom[101070] = 12'hbbb;
rom[101071] = 12'hccc;
rom[101072] = 12'hddd;
rom[101073] = 12'hddd;
rom[101074] = 12'heee;
rom[101075] = 12'hfff;
rom[101076] = 12'hfff;
rom[101077] = 12'hfff;
rom[101078] = 12'hfff;
rom[101079] = 12'hfff;
rom[101080] = 12'heee;
rom[101081] = 12'hddd;
rom[101082] = 12'hccc;
rom[101083] = 12'hccc;
rom[101084] = 12'hccc;
rom[101085] = 12'hddd;
rom[101086] = 12'hddd;
rom[101087] = 12'hddd;
rom[101088] = 12'hccc;
rom[101089] = 12'hbbb;
rom[101090] = 12'haaa;
rom[101091] = 12'haaa;
rom[101092] = 12'h999;
rom[101093] = 12'h888;
rom[101094] = 12'h777;
rom[101095] = 12'h666;
rom[101096] = 12'h555;
rom[101097] = 12'h555;
rom[101098] = 12'h444;
rom[101099] = 12'h333;
rom[101100] = 12'h333;
rom[101101] = 12'h333;
rom[101102] = 12'h333;
rom[101103] = 12'h333;
rom[101104] = 12'h444;
rom[101105] = 12'h333;
rom[101106] = 12'h333;
rom[101107] = 12'h333;
rom[101108] = 12'h333;
rom[101109] = 12'h444;
rom[101110] = 12'h888;
rom[101111] = 12'hbbb;
rom[101112] = 12'heee;
rom[101113] = 12'hddd;
rom[101114] = 12'hbbb;
rom[101115] = 12'h888;
rom[101116] = 12'h666;
rom[101117] = 12'h555;
rom[101118] = 12'h555;
rom[101119] = 12'h555;
rom[101120] = 12'h777;
rom[101121] = 12'h666;
rom[101122] = 12'h666;
rom[101123] = 12'h555;
rom[101124] = 12'h444;
rom[101125] = 12'h333;
rom[101126] = 12'h333;
rom[101127] = 12'h333;
rom[101128] = 12'h444;
rom[101129] = 12'h333;
rom[101130] = 12'h333;
rom[101131] = 12'h333;
rom[101132] = 12'h444;
rom[101133] = 12'h555;
rom[101134] = 12'h777;
rom[101135] = 12'haaa;
rom[101136] = 12'hddd;
rom[101137] = 12'heee;
rom[101138] = 12'hfff;
rom[101139] = 12'hddd;
rom[101140] = 12'haaa;
rom[101141] = 12'h777;
rom[101142] = 12'h555;
rom[101143] = 12'h444;
rom[101144] = 12'h333;
rom[101145] = 12'h222;
rom[101146] = 12'h222;
rom[101147] = 12'h222;
rom[101148] = 12'h222;
rom[101149] = 12'h222;
rom[101150] = 12'h111;
rom[101151] = 12'h111;
rom[101152] = 12'h111;
rom[101153] = 12'h111;
rom[101154] = 12'h111;
rom[101155] = 12'h111;
rom[101156] = 12'h111;
rom[101157] = 12'h111;
rom[101158] = 12'h111;
rom[101159] = 12'h111;
rom[101160] = 12'h111;
rom[101161] = 12'h111;
rom[101162] = 12'h111;
rom[101163] = 12'h111;
rom[101164] = 12'h  0;
rom[101165] = 12'h  0;
rom[101166] = 12'h  0;
rom[101167] = 12'h  0;
rom[101168] = 12'h  0;
rom[101169] = 12'h  0;
rom[101170] = 12'h  0;
rom[101171] = 12'h  0;
rom[101172] = 12'h  0;
rom[101173] = 12'h  0;
rom[101174] = 12'h  0;
rom[101175] = 12'h  0;
rom[101176] = 12'h  0;
rom[101177] = 12'h  0;
rom[101178] = 12'h  0;
rom[101179] = 12'h  0;
rom[101180] = 12'h  0;
rom[101181] = 12'h111;
rom[101182] = 12'h111;
rom[101183] = 12'h111;
rom[101184] = 12'h111;
rom[101185] = 12'h111;
rom[101186] = 12'h  0;
rom[101187] = 12'h111;
rom[101188] = 12'h222;
rom[101189] = 12'h333;
rom[101190] = 12'h333;
rom[101191] = 12'h333;
rom[101192] = 12'h222;
rom[101193] = 12'h111;
rom[101194] = 12'h111;
rom[101195] = 12'h111;
rom[101196] = 12'h111;
rom[101197] = 12'h111;
rom[101198] = 12'h  0;
rom[101199] = 12'h  0;
rom[101200] = 12'hfff;
rom[101201] = 12'hfff;
rom[101202] = 12'hfff;
rom[101203] = 12'hfff;
rom[101204] = 12'hfff;
rom[101205] = 12'hfff;
rom[101206] = 12'hfff;
rom[101207] = 12'hfff;
rom[101208] = 12'hfff;
rom[101209] = 12'hfff;
rom[101210] = 12'hfff;
rom[101211] = 12'hfff;
rom[101212] = 12'hfff;
rom[101213] = 12'hfff;
rom[101214] = 12'hfff;
rom[101215] = 12'hfff;
rom[101216] = 12'hfff;
rom[101217] = 12'hfff;
rom[101218] = 12'hfff;
rom[101219] = 12'hfff;
rom[101220] = 12'hfff;
rom[101221] = 12'hfff;
rom[101222] = 12'hfff;
rom[101223] = 12'hfff;
rom[101224] = 12'hfff;
rom[101225] = 12'hfff;
rom[101226] = 12'hfff;
rom[101227] = 12'hfff;
rom[101228] = 12'hfff;
rom[101229] = 12'hfff;
rom[101230] = 12'hfff;
rom[101231] = 12'hfff;
rom[101232] = 12'hfff;
rom[101233] = 12'hfff;
rom[101234] = 12'hfff;
rom[101235] = 12'hfff;
rom[101236] = 12'hfff;
rom[101237] = 12'hfff;
rom[101238] = 12'hfff;
rom[101239] = 12'hfff;
rom[101240] = 12'hfff;
rom[101241] = 12'hfff;
rom[101242] = 12'hfff;
rom[101243] = 12'hfff;
rom[101244] = 12'hfff;
rom[101245] = 12'hfff;
rom[101246] = 12'hfff;
rom[101247] = 12'hfff;
rom[101248] = 12'hfff;
rom[101249] = 12'hfff;
rom[101250] = 12'hfff;
rom[101251] = 12'hfff;
rom[101252] = 12'hfff;
rom[101253] = 12'hfff;
rom[101254] = 12'hfff;
rom[101255] = 12'hfff;
rom[101256] = 12'hfff;
rom[101257] = 12'hfff;
rom[101258] = 12'hfff;
rom[101259] = 12'hfff;
rom[101260] = 12'hfff;
rom[101261] = 12'hfff;
rom[101262] = 12'hfff;
rom[101263] = 12'hfff;
rom[101264] = 12'hfff;
rom[101265] = 12'hfff;
rom[101266] = 12'hfff;
rom[101267] = 12'hfff;
rom[101268] = 12'hfff;
rom[101269] = 12'hfff;
rom[101270] = 12'hfff;
rom[101271] = 12'hfff;
rom[101272] = 12'heee;
rom[101273] = 12'hfff;
rom[101274] = 12'hfff;
rom[101275] = 12'hfff;
rom[101276] = 12'hfff;
rom[101277] = 12'hfff;
rom[101278] = 12'heee;
rom[101279] = 12'heee;
rom[101280] = 12'heee;
rom[101281] = 12'heee;
rom[101282] = 12'heee;
rom[101283] = 12'heee;
rom[101284] = 12'heee;
rom[101285] = 12'heee;
rom[101286] = 12'heee;
rom[101287] = 12'heee;
rom[101288] = 12'hfff;
rom[101289] = 12'hfff;
rom[101290] = 12'hfff;
rom[101291] = 12'hfff;
rom[101292] = 12'hfff;
rom[101293] = 12'hfff;
rom[101294] = 12'hfff;
rom[101295] = 12'hfff;
rom[101296] = 12'heee;
rom[101297] = 12'heee;
rom[101298] = 12'heee;
rom[101299] = 12'heee;
rom[101300] = 12'heee;
rom[101301] = 12'heee;
rom[101302] = 12'heee;
rom[101303] = 12'heee;
rom[101304] = 12'heee;
rom[101305] = 12'heee;
rom[101306] = 12'hfff;
rom[101307] = 12'hfff;
rom[101308] = 12'hfff;
rom[101309] = 12'heee;
rom[101310] = 12'hfff;
rom[101311] = 12'hfff;
rom[101312] = 12'hfff;
rom[101313] = 12'hfff;
rom[101314] = 12'hfff;
rom[101315] = 12'hfff;
rom[101316] = 12'hfff;
rom[101317] = 12'hfff;
rom[101318] = 12'hfff;
rom[101319] = 12'hfff;
rom[101320] = 12'hfff;
rom[101321] = 12'hfff;
rom[101322] = 12'hfff;
rom[101323] = 12'hfff;
rom[101324] = 12'hfff;
rom[101325] = 12'hfff;
rom[101326] = 12'hfff;
rom[101327] = 12'hfff;
rom[101328] = 12'hfff;
rom[101329] = 12'hfff;
rom[101330] = 12'hfff;
rom[101331] = 12'hfff;
rom[101332] = 12'hfff;
rom[101333] = 12'hfff;
rom[101334] = 12'hfff;
rom[101335] = 12'hfff;
rom[101336] = 12'hfff;
rom[101337] = 12'hfff;
rom[101338] = 12'hfff;
rom[101339] = 12'hfff;
rom[101340] = 12'hfff;
rom[101341] = 12'hfff;
rom[101342] = 12'hfff;
rom[101343] = 12'hfff;
rom[101344] = 12'hfff;
rom[101345] = 12'hfff;
rom[101346] = 12'hfff;
rom[101347] = 12'hfff;
rom[101348] = 12'hfff;
rom[101349] = 12'hfff;
rom[101350] = 12'hfff;
rom[101351] = 12'hfff;
rom[101352] = 12'hfff;
rom[101353] = 12'hfff;
rom[101354] = 12'hfff;
rom[101355] = 12'hfff;
rom[101356] = 12'hfff;
rom[101357] = 12'hfff;
rom[101358] = 12'hfff;
rom[101359] = 12'hfff;
rom[101360] = 12'hfff;
rom[101361] = 12'hfff;
rom[101362] = 12'hfff;
rom[101363] = 12'hfff;
rom[101364] = 12'hfff;
rom[101365] = 12'hfff;
rom[101366] = 12'hfff;
rom[101367] = 12'hfff;
rom[101368] = 12'heee;
rom[101369] = 12'heee;
rom[101370] = 12'heee;
rom[101371] = 12'heee;
rom[101372] = 12'heee;
rom[101373] = 12'heee;
rom[101374] = 12'hddd;
rom[101375] = 12'hddd;
rom[101376] = 12'hddd;
rom[101377] = 12'hddd;
rom[101378] = 12'hddd;
rom[101379] = 12'hddd;
rom[101380] = 12'hddd;
rom[101381] = 12'hddd;
rom[101382] = 12'hddd;
rom[101383] = 12'hddd;
rom[101384] = 12'hddd;
rom[101385] = 12'hddd;
rom[101386] = 12'hddd;
rom[101387] = 12'hddd;
rom[101388] = 12'hddd;
rom[101389] = 12'hddd;
rom[101390] = 12'hddd;
rom[101391] = 12'hddd;
rom[101392] = 12'hccc;
rom[101393] = 12'hccc;
rom[101394] = 12'hccc;
rom[101395] = 12'hccc;
rom[101396] = 12'hccc;
rom[101397] = 12'hccc;
rom[101398] = 12'hccc;
rom[101399] = 12'hccc;
rom[101400] = 12'hccc;
rom[101401] = 12'hccc;
rom[101402] = 12'hccc;
rom[101403] = 12'hccc;
rom[101404] = 12'hccc;
rom[101405] = 12'hddd;
rom[101406] = 12'hddd;
rom[101407] = 12'hddd;
rom[101408] = 12'hddd;
rom[101409] = 12'hddd;
rom[101410] = 12'hddd;
rom[101411] = 12'hddd;
rom[101412] = 12'hddd;
rom[101413] = 12'hddd;
rom[101414] = 12'hddd;
rom[101415] = 12'hddd;
rom[101416] = 12'hddd;
rom[101417] = 12'hddd;
rom[101418] = 12'heee;
rom[101419] = 12'heee;
rom[101420] = 12'heee;
rom[101421] = 12'heee;
rom[101422] = 12'heee;
rom[101423] = 12'heee;
rom[101424] = 12'heee;
rom[101425] = 12'heee;
rom[101426] = 12'heee;
rom[101427] = 12'heee;
rom[101428] = 12'heee;
rom[101429] = 12'heee;
rom[101430] = 12'heee;
rom[101431] = 12'heee;
rom[101432] = 12'heee;
rom[101433] = 12'heee;
rom[101434] = 12'heee;
rom[101435] = 12'heee;
rom[101436] = 12'heee;
rom[101437] = 12'heee;
rom[101438] = 12'heee;
rom[101439] = 12'heee;
rom[101440] = 12'heee;
rom[101441] = 12'hddd;
rom[101442] = 12'hddd;
rom[101443] = 12'hddd;
rom[101444] = 12'hddd;
rom[101445] = 12'hddd;
rom[101446] = 12'hddd;
rom[101447] = 12'hccc;
rom[101448] = 12'hccc;
rom[101449] = 12'hccc;
rom[101450] = 12'hccc;
rom[101451] = 12'hccc;
rom[101452] = 12'hccc;
rom[101453] = 12'hbbb;
rom[101454] = 12'hbbb;
rom[101455] = 12'hbbb;
rom[101456] = 12'haaa;
rom[101457] = 12'haaa;
rom[101458] = 12'haaa;
rom[101459] = 12'haaa;
rom[101460] = 12'haaa;
rom[101461] = 12'haaa;
rom[101462] = 12'haaa;
rom[101463] = 12'haaa;
rom[101464] = 12'haaa;
rom[101465] = 12'hbbb;
rom[101466] = 12'hbbb;
rom[101467] = 12'hbbb;
rom[101468] = 12'hbbb;
rom[101469] = 12'hccc;
rom[101470] = 12'hddd;
rom[101471] = 12'hddd;
rom[101472] = 12'heee;
rom[101473] = 12'heee;
rom[101474] = 12'hfff;
rom[101475] = 12'hfff;
rom[101476] = 12'hfff;
rom[101477] = 12'hfff;
rom[101478] = 12'hfff;
rom[101479] = 12'heee;
rom[101480] = 12'hccc;
rom[101481] = 12'hccc;
rom[101482] = 12'hbbb;
rom[101483] = 12'hbbb;
rom[101484] = 12'hccc;
rom[101485] = 12'hddd;
rom[101486] = 12'hddd;
rom[101487] = 12'hddd;
rom[101488] = 12'hddd;
rom[101489] = 12'hccc;
rom[101490] = 12'hbbb;
rom[101491] = 12'haaa;
rom[101492] = 12'haaa;
rom[101493] = 12'h999;
rom[101494] = 12'h777;
rom[101495] = 12'h777;
rom[101496] = 12'h555;
rom[101497] = 12'h555;
rom[101498] = 12'h444;
rom[101499] = 12'h333;
rom[101500] = 12'h333;
rom[101501] = 12'h333;
rom[101502] = 12'h333;
rom[101503] = 12'h333;
rom[101504] = 12'h333;
rom[101505] = 12'h222;
rom[101506] = 12'h222;
rom[101507] = 12'h333;
rom[101508] = 12'h333;
rom[101509] = 12'h333;
rom[101510] = 12'h444;
rom[101511] = 12'h666;
rom[101512] = 12'haaa;
rom[101513] = 12'hccc;
rom[101514] = 12'heee;
rom[101515] = 12'hccc;
rom[101516] = 12'h888;
rom[101517] = 12'h666;
rom[101518] = 12'h555;
rom[101519] = 12'h555;
rom[101520] = 12'h666;
rom[101521] = 12'h666;
rom[101522] = 12'h666;
rom[101523] = 12'h555;
rom[101524] = 12'h444;
rom[101525] = 12'h333;
rom[101526] = 12'h333;
rom[101527] = 12'h333;
rom[101528] = 12'h444;
rom[101529] = 12'h333;
rom[101530] = 12'h222;
rom[101531] = 12'h333;
rom[101532] = 12'h444;
rom[101533] = 12'h444;
rom[101534] = 12'h444;
rom[101535] = 12'h555;
rom[101536] = 12'h999;
rom[101537] = 12'hccc;
rom[101538] = 12'hfff;
rom[101539] = 12'hfff;
rom[101540] = 12'heee;
rom[101541] = 12'hbbb;
rom[101542] = 12'h888;
rom[101543] = 12'h666;
rom[101544] = 12'h444;
rom[101545] = 12'h333;
rom[101546] = 12'h333;
rom[101547] = 12'h222;
rom[101548] = 12'h222;
rom[101549] = 12'h222;
rom[101550] = 12'h111;
rom[101551] = 12'h222;
rom[101552] = 12'h111;
rom[101553] = 12'h111;
rom[101554] = 12'h111;
rom[101555] = 12'h111;
rom[101556] = 12'h111;
rom[101557] = 12'h111;
rom[101558] = 12'h111;
rom[101559] = 12'h111;
rom[101560] = 12'h111;
rom[101561] = 12'h111;
rom[101562] = 12'h111;
rom[101563] = 12'h111;
rom[101564] = 12'h  0;
rom[101565] = 12'h  0;
rom[101566] = 12'h  0;
rom[101567] = 12'h  0;
rom[101568] = 12'h  0;
rom[101569] = 12'h  0;
rom[101570] = 12'h  0;
rom[101571] = 12'h  0;
rom[101572] = 12'h  0;
rom[101573] = 12'h  0;
rom[101574] = 12'h  0;
rom[101575] = 12'h  0;
rom[101576] = 12'h  0;
rom[101577] = 12'h  0;
rom[101578] = 12'h  0;
rom[101579] = 12'h  0;
rom[101580] = 12'h  0;
rom[101581] = 12'h  0;
rom[101582] = 12'h  0;
rom[101583] = 12'h111;
rom[101584] = 12'h111;
rom[101585] = 12'h111;
rom[101586] = 12'h  0;
rom[101587] = 12'h111;
rom[101588] = 12'h111;
rom[101589] = 12'h222;
rom[101590] = 12'h222;
rom[101591] = 12'h222;
rom[101592] = 12'h222;
rom[101593] = 12'h222;
rom[101594] = 12'h111;
rom[101595] = 12'h111;
rom[101596] = 12'h  0;
rom[101597] = 12'h  0;
rom[101598] = 12'h  0;
rom[101599] = 12'h  0;
rom[101600] = 12'hfff;
rom[101601] = 12'hfff;
rom[101602] = 12'hfff;
rom[101603] = 12'hfff;
rom[101604] = 12'hfff;
rom[101605] = 12'hfff;
rom[101606] = 12'hfff;
rom[101607] = 12'hfff;
rom[101608] = 12'hfff;
rom[101609] = 12'hfff;
rom[101610] = 12'hfff;
rom[101611] = 12'hfff;
rom[101612] = 12'hfff;
rom[101613] = 12'hfff;
rom[101614] = 12'hfff;
rom[101615] = 12'hfff;
rom[101616] = 12'hfff;
rom[101617] = 12'hfff;
rom[101618] = 12'hfff;
rom[101619] = 12'hfff;
rom[101620] = 12'hfff;
rom[101621] = 12'hfff;
rom[101622] = 12'hfff;
rom[101623] = 12'hfff;
rom[101624] = 12'hfff;
rom[101625] = 12'hfff;
rom[101626] = 12'hfff;
rom[101627] = 12'hfff;
rom[101628] = 12'hfff;
rom[101629] = 12'hfff;
rom[101630] = 12'hfff;
rom[101631] = 12'hfff;
rom[101632] = 12'hfff;
rom[101633] = 12'hfff;
rom[101634] = 12'hfff;
rom[101635] = 12'hfff;
rom[101636] = 12'hfff;
rom[101637] = 12'hfff;
rom[101638] = 12'hfff;
rom[101639] = 12'hfff;
rom[101640] = 12'hfff;
rom[101641] = 12'hfff;
rom[101642] = 12'hfff;
rom[101643] = 12'hfff;
rom[101644] = 12'hfff;
rom[101645] = 12'hfff;
rom[101646] = 12'hfff;
rom[101647] = 12'hfff;
rom[101648] = 12'hfff;
rom[101649] = 12'hfff;
rom[101650] = 12'hfff;
rom[101651] = 12'hfff;
rom[101652] = 12'hfff;
rom[101653] = 12'hfff;
rom[101654] = 12'hfff;
rom[101655] = 12'hfff;
rom[101656] = 12'hfff;
rom[101657] = 12'hfff;
rom[101658] = 12'hfff;
rom[101659] = 12'hfff;
rom[101660] = 12'hfff;
rom[101661] = 12'hfff;
rom[101662] = 12'hfff;
rom[101663] = 12'hfff;
rom[101664] = 12'hfff;
rom[101665] = 12'hfff;
rom[101666] = 12'heee;
rom[101667] = 12'heee;
rom[101668] = 12'heee;
rom[101669] = 12'heee;
rom[101670] = 12'heee;
rom[101671] = 12'heee;
rom[101672] = 12'hfff;
rom[101673] = 12'hfff;
rom[101674] = 12'hfff;
rom[101675] = 12'hfff;
rom[101676] = 12'hfff;
rom[101677] = 12'heee;
rom[101678] = 12'heee;
rom[101679] = 12'heee;
rom[101680] = 12'heee;
rom[101681] = 12'heee;
rom[101682] = 12'heee;
rom[101683] = 12'heee;
rom[101684] = 12'heee;
rom[101685] = 12'heee;
rom[101686] = 12'heee;
rom[101687] = 12'heee;
rom[101688] = 12'hfff;
rom[101689] = 12'hfff;
rom[101690] = 12'hfff;
rom[101691] = 12'hfff;
rom[101692] = 12'hfff;
rom[101693] = 12'hfff;
rom[101694] = 12'heee;
rom[101695] = 12'heee;
rom[101696] = 12'heee;
rom[101697] = 12'heee;
rom[101698] = 12'heee;
rom[101699] = 12'heee;
rom[101700] = 12'heee;
rom[101701] = 12'heee;
rom[101702] = 12'heee;
rom[101703] = 12'heee;
rom[101704] = 12'heee;
rom[101705] = 12'hfff;
rom[101706] = 12'hfff;
rom[101707] = 12'hfff;
rom[101708] = 12'heee;
rom[101709] = 12'heee;
rom[101710] = 12'heee;
rom[101711] = 12'heee;
rom[101712] = 12'hfff;
rom[101713] = 12'hfff;
rom[101714] = 12'hfff;
rom[101715] = 12'hfff;
rom[101716] = 12'hfff;
rom[101717] = 12'hfff;
rom[101718] = 12'hfff;
rom[101719] = 12'hfff;
rom[101720] = 12'hfff;
rom[101721] = 12'hfff;
rom[101722] = 12'hfff;
rom[101723] = 12'hfff;
rom[101724] = 12'hfff;
rom[101725] = 12'hfff;
rom[101726] = 12'hfff;
rom[101727] = 12'hfff;
rom[101728] = 12'hfff;
rom[101729] = 12'hfff;
rom[101730] = 12'hfff;
rom[101731] = 12'hfff;
rom[101732] = 12'hfff;
rom[101733] = 12'hfff;
rom[101734] = 12'hfff;
rom[101735] = 12'hfff;
rom[101736] = 12'hfff;
rom[101737] = 12'hfff;
rom[101738] = 12'hfff;
rom[101739] = 12'hfff;
rom[101740] = 12'hfff;
rom[101741] = 12'hfff;
rom[101742] = 12'hfff;
rom[101743] = 12'hfff;
rom[101744] = 12'hfff;
rom[101745] = 12'hfff;
rom[101746] = 12'hfff;
rom[101747] = 12'hfff;
rom[101748] = 12'hfff;
rom[101749] = 12'hfff;
rom[101750] = 12'hfff;
rom[101751] = 12'hfff;
rom[101752] = 12'hfff;
rom[101753] = 12'hfff;
rom[101754] = 12'hfff;
rom[101755] = 12'hfff;
rom[101756] = 12'hfff;
rom[101757] = 12'hfff;
rom[101758] = 12'hfff;
rom[101759] = 12'hfff;
rom[101760] = 12'hfff;
rom[101761] = 12'hfff;
rom[101762] = 12'hfff;
rom[101763] = 12'hfff;
rom[101764] = 12'hfff;
rom[101765] = 12'hfff;
rom[101766] = 12'hfff;
rom[101767] = 12'hfff;
rom[101768] = 12'hfff;
rom[101769] = 12'hfff;
rom[101770] = 12'hfff;
rom[101771] = 12'hfff;
rom[101772] = 12'hfff;
rom[101773] = 12'heee;
rom[101774] = 12'heee;
rom[101775] = 12'heee;
rom[101776] = 12'heee;
rom[101777] = 12'heee;
rom[101778] = 12'heee;
rom[101779] = 12'heee;
rom[101780] = 12'hddd;
rom[101781] = 12'hddd;
rom[101782] = 12'hddd;
rom[101783] = 12'hddd;
rom[101784] = 12'hddd;
rom[101785] = 12'hddd;
rom[101786] = 12'hddd;
rom[101787] = 12'hddd;
rom[101788] = 12'hddd;
rom[101789] = 12'hddd;
rom[101790] = 12'hddd;
rom[101791] = 12'hddd;
rom[101792] = 12'hddd;
rom[101793] = 12'hddd;
rom[101794] = 12'hddd;
rom[101795] = 12'hddd;
rom[101796] = 12'hddd;
rom[101797] = 12'hddd;
rom[101798] = 12'hddd;
rom[101799] = 12'hddd;
rom[101800] = 12'hddd;
rom[101801] = 12'hddd;
rom[101802] = 12'hddd;
rom[101803] = 12'hddd;
rom[101804] = 12'hddd;
rom[101805] = 12'hddd;
rom[101806] = 12'hddd;
rom[101807] = 12'hddd;
rom[101808] = 12'hddd;
rom[101809] = 12'hddd;
rom[101810] = 12'hddd;
rom[101811] = 12'hddd;
rom[101812] = 12'hddd;
rom[101813] = 12'hddd;
rom[101814] = 12'heee;
rom[101815] = 12'heee;
rom[101816] = 12'heee;
rom[101817] = 12'heee;
rom[101818] = 12'heee;
rom[101819] = 12'heee;
rom[101820] = 12'heee;
rom[101821] = 12'heee;
rom[101822] = 12'heee;
rom[101823] = 12'heee;
rom[101824] = 12'hfff;
rom[101825] = 12'heee;
rom[101826] = 12'heee;
rom[101827] = 12'heee;
rom[101828] = 12'heee;
rom[101829] = 12'hfff;
rom[101830] = 12'hfff;
rom[101831] = 12'hfff;
rom[101832] = 12'heee;
rom[101833] = 12'heee;
rom[101834] = 12'heee;
rom[101835] = 12'heee;
rom[101836] = 12'heee;
rom[101837] = 12'heee;
rom[101838] = 12'heee;
rom[101839] = 12'heee;
rom[101840] = 12'heee;
rom[101841] = 12'heee;
rom[101842] = 12'hddd;
rom[101843] = 12'hddd;
rom[101844] = 12'hddd;
rom[101845] = 12'hddd;
rom[101846] = 12'hddd;
rom[101847] = 12'hddd;
rom[101848] = 12'hddd;
rom[101849] = 12'hccc;
rom[101850] = 12'hccc;
rom[101851] = 12'hccc;
rom[101852] = 12'hccc;
rom[101853] = 12'hccc;
rom[101854] = 12'hbbb;
rom[101855] = 12'hbbb;
rom[101856] = 12'hbbb;
rom[101857] = 12'hbbb;
rom[101858] = 12'hbbb;
rom[101859] = 12'hbbb;
rom[101860] = 12'hbbb;
rom[101861] = 12'hbbb;
rom[101862] = 12'hbbb;
rom[101863] = 12'hbbb;
rom[101864] = 12'hbbb;
rom[101865] = 12'hccc;
rom[101866] = 12'hccc;
rom[101867] = 12'hccc;
rom[101868] = 12'hddd;
rom[101869] = 12'hddd;
rom[101870] = 12'heee;
rom[101871] = 12'heee;
rom[101872] = 12'hfff;
rom[101873] = 12'hfff;
rom[101874] = 12'hfff;
rom[101875] = 12'hfff;
rom[101876] = 12'hfff;
rom[101877] = 12'heee;
rom[101878] = 12'hddd;
rom[101879] = 12'hccc;
rom[101880] = 12'hbbb;
rom[101881] = 12'haaa;
rom[101882] = 12'haaa;
rom[101883] = 12'haaa;
rom[101884] = 12'hbbb;
rom[101885] = 12'hccc;
rom[101886] = 12'hddd;
rom[101887] = 12'hddd;
rom[101888] = 12'hddd;
rom[101889] = 12'hddd;
rom[101890] = 12'hccc;
rom[101891] = 12'hbbb;
rom[101892] = 12'haaa;
rom[101893] = 12'h999;
rom[101894] = 12'h888;
rom[101895] = 12'h888;
rom[101896] = 12'h666;
rom[101897] = 12'h555;
rom[101898] = 12'h444;
rom[101899] = 12'h444;
rom[101900] = 12'h333;
rom[101901] = 12'h333;
rom[101902] = 12'h222;
rom[101903] = 12'h222;
rom[101904] = 12'h222;
rom[101905] = 12'h333;
rom[101906] = 12'h333;
rom[101907] = 12'h333;
rom[101908] = 12'h333;
rom[101909] = 12'h333;
rom[101910] = 12'h333;
rom[101911] = 12'h333;
rom[101912] = 12'h555;
rom[101913] = 12'h999;
rom[101914] = 12'hccc;
rom[101915] = 12'hddd;
rom[101916] = 12'hccc;
rom[101917] = 12'h999;
rom[101918] = 12'h777;
rom[101919] = 12'h666;
rom[101920] = 12'h666;
rom[101921] = 12'h666;
rom[101922] = 12'h666;
rom[101923] = 12'h555;
rom[101924] = 12'h444;
rom[101925] = 12'h333;
rom[101926] = 12'h333;
rom[101927] = 12'h444;
rom[101928] = 12'h333;
rom[101929] = 12'h222;
rom[101930] = 12'h222;
rom[101931] = 12'h333;
rom[101932] = 12'h333;
rom[101933] = 12'h444;
rom[101934] = 12'h333;
rom[101935] = 12'h333;
rom[101936] = 12'h555;
rom[101937] = 12'h777;
rom[101938] = 12'haaa;
rom[101939] = 12'hddd;
rom[101940] = 12'heee;
rom[101941] = 12'heee;
rom[101942] = 12'hccc;
rom[101943] = 12'haaa;
rom[101944] = 12'h777;
rom[101945] = 12'h555;
rom[101946] = 12'h444;
rom[101947] = 12'h333;
rom[101948] = 12'h333;
rom[101949] = 12'h222;
rom[101950] = 12'h222;
rom[101951] = 12'h222;
rom[101952] = 12'h111;
rom[101953] = 12'h111;
rom[101954] = 12'h111;
rom[101955] = 12'h111;
rom[101956] = 12'h111;
rom[101957] = 12'h111;
rom[101958] = 12'h111;
rom[101959] = 12'h111;
rom[101960] = 12'h111;
rom[101961] = 12'h111;
rom[101962] = 12'h111;
rom[101963] = 12'h  0;
rom[101964] = 12'h  0;
rom[101965] = 12'h  0;
rom[101966] = 12'h  0;
rom[101967] = 12'h  0;
rom[101968] = 12'h  0;
rom[101969] = 12'h  0;
rom[101970] = 12'h  0;
rom[101971] = 12'h  0;
rom[101972] = 12'h  0;
rom[101973] = 12'h  0;
rom[101974] = 12'h  0;
rom[101975] = 12'h  0;
rom[101976] = 12'h  0;
rom[101977] = 12'h  0;
rom[101978] = 12'h  0;
rom[101979] = 12'h  0;
rom[101980] = 12'h  0;
rom[101981] = 12'h  0;
rom[101982] = 12'h  0;
rom[101983] = 12'h  0;
rom[101984] = 12'h  0;
rom[101985] = 12'h  0;
rom[101986] = 12'h  0;
rom[101987] = 12'h111;
rom[101988] = 12'h111;
rom[101989] = 12'h111;
rom[101990] = 12'h222;
rom[101991] = 12'h222;
rom[101992] = 12'h222;
rom[101993] = 12'h222;
rom[101994] = 12'h111;
rom[101995] = 12'h111;
rom[101996] = 12'h  0;
rom[101997] = 12'h  0;
rom[101998] = 12'h  0;
rom[101999] = 12'h  0;
rom[102000] = 12'hfff;
rom[102001] = 12'hfff;
rom[102002] = 12'hfff;
rom[102003] = 12'hfff;
rom[102004] = 12'hfff;
rom[102005] = 12'hfff;
rom[102006] = 12'hfff;
rom[102007] = 12'hfff;
rom[102008] = 12'hfff;
rom[102009] = 12'hfff;
rom[102010] = 12'hfff;
rom[102011] = 12'hfff;
rom[102012] = 12'hfff;
rom[102013] = 12'hfff;
rom[102014] = 12'hfff;
rom[102015] = 12'hfff;
rom[102016] = 12'hfff;
rom[102017] = 12'hfff;
rom[102018] = 12'hfff;
rom[102019] = 12'hfff;
rom[102020] = 12'hfff;
rom[102021] = 12'hfff;
rom[102022] = 12'hfff;
rom[102023] = 12'hfff;
rom[102024] = 12'hfff;
rom[102025] = 12'hfff;
rom[102026] = 12'hfff;
rom[102027] = 12'hfff;
rom[102028] = 12'hfff;
rom[102029] = 12'hfff;
rom[102030] = 12'hfff;
rom[102031] = 12'hfff;
rom[102032] = 12'hfff;
rom[102033] = 12'hfff;
rom[102034] = 12'hfff;
rom[102035] = 12'hfff;
rom[102036] = 12'hfff;
rom[102037] = 12'hfff;
rom[102038] = 12'hfff;
rom[102039] = 12'hfff;
rom[102040] = 12'hfff;
rom[102041] = 12'hfff;
rom[102042] = 12'hfff;
rom[102043] = 12'hfff;
rom[102044] = 12'hfff;
rom[102045] = 12'hfff;
rom[102046] = 12'hfff;
rom[102047] = 12'hfff;
rom[102048] = 12'hfff;
rom[102049] = 12'hfff;
rom[102050] = 12'hfff;
rom[102051] = 12'hfff;
rom[102052] = 12'hfff;
rom[102053] = 12'hfff;
rom[102054] = 12'hfff;
rom[102055] = 12'hfff;
rom[102056] = 12'hfff;
rom[102057] = 12'hfff;
rom[102058] = 12'hfff;
rom[102059] = 12'hfff;
rom[102060] = 12'hfff;
rom[102061] = 12'hfff;
rom[102062] = 12'hfff;
rom[102063] = 12'hfff;
rom[102064] = 12'heee;
rom[102065] = 12'heee;
rom[102066] = 12'heee;
rom[102067] = 12'heee;
rom[102068] = 12'heee;
rom[102069] = 12'heee;
rom[102070] = 12'heee;
rom[102071] = 12'heee;
rom[102072] = 12'hfff;
rom[102073] = 12'hfff;
rom[102074] = 12'hfff;
rom[102075] = 12'hfff;
rom[102076] = 12'hfff;
rom[102077] = 12'heee;
rom[102078] = 12'heee;
rom[102079] = 12'heee;
rom[102080] = 12'heee;
rom[102081] = 12'heee;
rom[102082] = 12'heee;
rom[102083] = 12'heee;
rom[102084] = 12'heee;
rom[102085] = 12'heee;
rom[102086] = 12'heee;
rom[102087] = 12'heee;
rom[102088] = 12'hfff;
rom[102089] = 12'hfff;
rom[102090] = 12'hfff;
rom[102091] = 12'hfff;
rom[102092] = 12'hfff;
rom[102093] = 12'heee;
rom[102094] = 12'heee;
rom[102095] = 12'heee;
rom[102096] = 12'hddd;
rom[102097] = 12'hddd;
rom[102098] = 12'heee;
rom[102099] = 12'heee;
rom[102100] = 12'heee;
rom[102101] = 12'heee;
rom[102102] = 12'heee;
rom[102103] = 12'heee;
rom[102104] = 12'hfff;
rom[102105] = 12'hfff;
rom[102106] = 12'hfff;
rom[102107] = 12'hfff;
rom[102108] = 12'heee;
rom[102109] = 12'heee;
rom[102110] = 12'heee;
rom[102111] = 12'heee;
rom[102112] = 12'hfff;
rom[102113] = 12'hfff;
rom[102114] = 12'hfff;
rom[102115] = 12'hfff;
rom[102116] = 12'hfff;
rom[102117] = 12'hfff;
rom[102118] = 12'hfff;
rom[102119] = 12'hfff;
rom[102120] = 12'hfff;
rom[102121] = 12'hfff;
rom[102122] = 12'hfff;
rom[102123] = 12'hfff;
rom[102124] = 12'hfff;
rom[102125] = 12'hfff;
rom[102126] = 12'hfff;
rom[102127] = 12'hfff;
rom[102128] = 12'hfff;
rom[102129] = 12'hfff;
rom[102130] = 12'hfff;
rom[102131] = 12'hfff;
rom[102132] = 12'hfff;
rom[102133] = 12'hfff;
rom[102134] = 12'hfff;
rom[102135] = 12'hfff;
rom[102136] = 12'hfff;
rom[102137] = 12'hfff;
rom[102138] = 12'hfff;
rom[102139] = 12'hfff;
rom[102140] = 12'hfff;
rom[102141] = 12'hfff;
rom[102142] = 12'hfff;
rom[102143] = 12'hfff;
rom[102144] = 12'hfff;
rom[102145] = 12'hfff;
rom[102146] = 12'hfff;
rom[102147] = 12'hfff;
rom[102148] = 12'hfff;
rom[102149] = 12'hfff;
rom[102150] = 12'hfff;
rom[102151] = 12'hfff;
rom[102152] = 12'hfff;
rom[102153] = 12'hfff;
rom[102154] = 12'hfff;
rom[102155] = 12'hfff;
rom[102156] = 12'hfff;
rom[102157] = 12'hfff;
rom[102158] = 12'hfff;
rom[102159] = 12'hfff;
rom[102160] = 12'hfff;
rom[102161] = 12'hfff;
rom[102162] = 12'hfff;
rom[102163] = 12'hfff;
rom[102164] = 12'hfff;
rom[102165] = 12'hfff;
rom[102166] = 12'hfff;
rom[102167] = 12'hfff;
rom[102168] = 12'hfff;
rom[102169] = 12'hfff;
rom[102170] = 12'hfff;
rom[102171] = 12'hfff;
rom[102172] = 12'hfff;
rom[102173] = 12'hfff;
rom[102174] = 12'hfff;
rom[102175] = 12'hfff;
rom[102176] = 12'heee;
rom[102177] = 12'heee;
rom[102178] = 12'heee;
rom[102179] = 12'heee;
rom[102180] = 12'heee;
rom[102181] = 12'heee;
rom[102182] = 12'heee;
rom[102183] = 12'heee;
rom[102184] = 12'hddd;
rom[102185] = 12'hddd;
rom[102186] = 12'hddd;
rom[102187] = 12'hddd;
rom[102188] = 12'hddd;
rom[102189] = 12'hddd;
rom[102190] = 12'hddd;
rom[102191] = 12'hddd;
rom[102192] = 12'hddd;
rom[102193] = 12'hddd;
rom[102194] = 12'hddd;
rom[102195] = 12'hddd;
rom[102196] = 12'hddd;
rom[102197] = 12'hddd;
rom[102198] = 12'hddd;
rom[102199] = 12'hddd;
rom[102200] = 12'hddd;
rom[102201] = 12'hddd;
rom[102202] = 12'hddd;
rom[102203] = 12'hddd;
rom[102204] = 12'hddd;
rom[102205] = 12'hddd;
rom[102206] = 12'hddd;
rom[102207] = 12'hddd;
rom[102208] = 12'heee;
rom[102209] = 12'heee;
rom[102210] = 12'heee;
rom[102211] = 12'heee;
rom[102212] = 12'heee;
rom[102213] = 12'heee;
rom[102214] = 12'heee;
rom[102215] = 12'heee;
rom[102216] = 12'heee;
rom[102217] = 12'heee;
rom[102218] = 12'heee;
rom[102219] = 12'hfff;
rom[102220] = 12'hfff;
rom[102221] = 12'hfff;
rom[102222] = 12'hfff;
rom[102223] = 12'hfff;
rom[102224] = 12'hfff;
rom[102225] = 12'hfff;
rom[102226] = 12'hfff;
rom[102227] = 12'hfff;
rom[102228] = 12'hfff;
rom[102229] = 12'hfff;
rom[102230] = 12'hfff;
rom[102231] = 12'hfff;
rom[102232] = 12'hfff;
rom[102233] = 12'hfff;
rom[102234] = 12'hfff;
rom[102235] = 12'hfff;
rom[102236] = 12'heee;
rom[102237] = 12'heee;
rom[102238] = 12'heee;
rom[102239] = 12'heee;
rom[102240] = 12'heee;
rom[102241] = 12'heee;
rom[102242] = 12'heee;
rom[102243] = 12'hddd;
rom[102244] = 12'hddd;
rom[102245] = 12'hddd;
rom[102246] = 12'hddd;
rom[102247] = 12'hddd;
rom[102248] = 12'hddd;
rom[102249] = 12'hddd;
rom[102250] = 12'hddd;
rom[102251] = 12'hddd;
rom[102252] = 12'hddd;
rom[102253] = 12'hccc;
rom[102254] = 12'hccc;
rom[102255] = 12'hccc;
rom[102256] = 12'hccc;
rom[102257] = 12'hccc;
rom[102258] = 12'hccc;
rom[102259] = 12'hccc;
rom[102260] = 12'hccc;
rom[102261] = 12'hccc;
rom[102262] = 12'hccc;
rom[102263] = 12'hccc;
rom[102264] = 12'hccc;
rom[102265] = 12'hddd;
rom[102266] = 12'hddd;
rom[102267] = 12'hddd;
rom[102268] = 12'heee;
rom[102269] = 12'heee;
rom[102270] = 12'hfff;
rom[102271] = 12'hfff;
rom[102272] = 12'hfff;
rom[102273] = 12'hfff;
rom[102274] = 12'hfff;
rom[102275] = 12'hfff;
rom[102276] = 12'heee;
rom[102277] = 12'hddd;
rom[102278] = 12'hccc;
rom[102279] = 12'hbbb;
rom[102280] = 12'haaa;
rom[102281] = 12'h999;
rom[102282] = 12'h999;
rom[102283] = 12'h999;
rom[102284] = 12'haaa;
rom[102285] = 12'hbbb;
rom[102286] = 12'hddd;
rom[102287] = 12'heee;
rom[102288] = 12'heee;
rom[102289] = 12'heee;
rom[102290] = 12'hddd;
rom[102291] = 12'hccc;
rom[102292] = 12'hbbb;
rom[102293] = 12'haaa;
rom[102294] = 12'h999;
rom[102295] = 12'h999;
rom[102296] = 12'h777;
rom[102297] = 12'h555;
rom[102298] = 12'h333;
rom[102299] = 12'h333;
rom[102300] = 12'h333;
rom[102301] = 12'h333;
rom[102302] = 12'h333;
rom[102303] = 12'h333;
rom[102304] = 12'h222;
rom[102305] = 12'h444;
rom[102306] = 12'h444;
rom[102307] = 12'h222;
rom[102308] = 12'h222;
rom[102309] = 12'h333;
rom[102310] = 12'h333;
rom[102311] = 12'h333;
rom[102312] = 12'h333;
rom[102313] = 12'h555;
rom[102314] = 12'h888;
rom[102315] = 12'hbbb;
rom[102316] = 12'hddd;
rom[102317] = 12'hddd;
rom[102318] = 12'haaa;
rom[102319] = 12'h777;
rom[102320] = 12'h555;
rom[102321] = 12'h666;
rom[102322] = 12'h666;
rom[102323] = 12'h666;
rom[102324] = 12'h555;
rom[102325] = 12'h333;
rom[102326] = 12'h222;
rom[102327] = 12'h222;
rom[102328] = 12'h222;
rom[102329] = 12'h333;
rom[102330] = 12'h333;
rom[102331] = 12'h222;
rom[102332] = 12'h222;
rom[102333] = 12'h333;
rom[102334] = 12'h333;
rom[102335] = 12'h333;
rom[102336] = 12'h333;
rom[102337] = 12'h444;
rom[102338] = 12'h666;
rom[102339] = 12'h999;
rom[102340] = 12'hddd;
rom[102341] = 12'hfff;
rom[102342] = 12'heee;
rom[102343] = 12'hccc;
rom[102344] = 12'h999;
rom[102345] = 12'h777;
rom[102346] = 12'h555;
rom[102347] = 12'h444;
rom[102348] = 12'h333;
rom[102349] = 12'h222;
rom[102350] = 12'h222;
rom[102351] = 12'h222;
rom[102352] = 12'h222;
rom[102353] = 12'h222;
rom[102354] = 12'h111;
rom[102355] = 12'h111;
rom[102356] = 12'h111;
rom[102357] = 12'h111;
rom[102358] = 12'h111;
rom[102359] = 12'h111;
rom[102360] = 12'h111;
rom[102361] = 12'h111;
rom[102362] = 12'h111;
rom[102363] = 12'h  0;
rom[102364] = 12'h  0;
rom[102365] = 12'h  0;
rom[102366] = 12'h  0;
rom[102367] = 12'h  0;
rom[102368] = 12'h  0;
rom[102369] = 12'h  0;
rom[102370] = 12'h  0;
rom[102371] = 12'h  0;
rom[102372] = 12'h  0;
rom[102373] = 12'h  0;
rom[102374] = 12'h  0;
rom[102375] = 12'h  0;
rom[102376] = 12'h  0;
rom[102377] = 12'h  0;
rom[102378] = 12'h  0;
rom[102379] = 12'h  0;
rom[102380] = 12'h  0;
rom[102381] = 12'h  0;
rom[102382] = 12'h  0;
rom[102383] = 12'h  0;
rom[102384] = 12'h  0;
rom[102385] = 12'h  0;
rom[102386] = 12'h  0;
rom[102387] = 12'h111;
rom[102388] = 12'h111;
rom[102389] = 12'h111;
rom[102390] = 12'h111;
rom[102391] = 12'h111;
rom[102392] = 12'h222;
rom[102393] = 12'h222;
rom[102394] = 12'h111;
rom[102395] = 12'h111;
rom[102396] = 12'h  0;
rom[102397] = 12'h  0;
rom[102398] = 12'h  0;
rom[102399] = 12'h  0;
rom[102400] = 12'hfff;
rom[102401] = 12'hfff;
rom[102402] = 12'hfff;
rom[102403] = 12'hfff;
rom[102404] = 12'hfff;
rom[102405] = 12'hfff;
rom[102406] = 12'hfff;
rom[102407] = 12'hfff;
rom[102408] = 12'hfff;
rom[102409] = 12'hfff;
rom[102410] = 12'hfff;
rom[102411] = 12'hfff;
rom[102412] = 12'hfff;
rom[102413] = 12'hfff;
rom[102414] = 12'hfff;
rom[102415] = 12'hfff;
rom[102416] = 12'hfff;
rom[102417] = 12'hfff;
rom[102418] = 12'hfff;
rom[102419] = 12'hfff;
rom[102420] = 12'hfff;
rom[102421] = 12'hfff;
rom[102422] = 12'hfff;
rom[102423] = 12'hfff;
rom[102424] = 12'hfff;
rom[102425] = 12'hfff;
rom[102426] = 12'hfff;
rom[102427] = 12'hfff;
rom[102428] = 12'hfff;
rom[102429] = 12'hfff;
rom[102430] = 12'hfff;
rom[102431] = 12'hfff;
rom[102432] = 12'hfff;
rom[102433] = 12'hfff;
rom[102434] = 12'hfff;
rom[102435] = 12'hfff;
rom[102436] = 12'hfff;
rom[102437] = 12'hfff;
rom[102438] = 12'hfff;
rom[102439] = 12'hfff;
rom[102440] = 12'hfff;
rom[102441] = 12'hfff;
rom[102442] = 12'hfff;
rom[102443] = 12'hfff;
rom[102444] = 12'hfff;
rom[102445] = 12'hfff;
rom[102446] = 12'hfff;
rom[102447] = 12'hfff;
rom[102448] = 12'hfff;
rom[102449] = 12'hfff;
rom[102450] = 12'hfff;
rom[102451] = 12'hfff;
rom[102452] = 12'hfff;
rom[102453] = 12'hfff;
rom[102454] = 12'hfff;
rom[102455] = 12'hfff;
rom[102456] = 12'hfff;
rom[102457] = 12'hfff;
rom[102458] = 12'hfff;
rom[102459] = 12'hfff;
rom[102460] = 12'hfff;
rom[102461] = 12'hfff;
rom[102462] = 12'hfff;
rom[102463] = 12'heee;
rom[102464] = 12'hfff;
rom[102465] = 12'heee;
rom[102466] = 12'heee;
rom[102467] = 12'heee;
rom[102468] = 12'heee;
rom[102469] = 12'heee;
rom[102470] = 12'heee;
rom[102471] = 12'heee;
rom[102472] = 12'hfff;
rom[102473] = 12'hfff;
rom[102474] = 12'hfff;
rom[102475] = 12'heee;
rom[102476] = 12'heee;
rom[102477] = 12'heee;
rom[102478] = 12'heee;
rom[102479] = 12'heee;
rom[102480] = 12'heee;
rom[102481] = 12'heee;
rom[102482] = 12'heee;
rom[102483] = 12'heee;
rom[102484] = 12'heee;
rom[102485] = 12'heee;
rom[102486] = 12'heee;
rom[102487] = 12'hfff;
rom[102488] = 12'hfff;
rom[102489] = 12'hfff;
rom[102490] = 12'hfff;
rom[102491] = 12'heee;
rom[102492] = 12'heee;
rom[102493] = 12'heee;
rom[102494] = 12'heee;
rom[102495] = 12'heee;
rom[102496] = 12'heee;
rom[102497] = 12'heee;
rom[102498] = 12'heee;
rom[102499] = 12'hddd;
rom[102500] = 12'hddd;
rom[102501] = 12'hddd;
rom[102502] = 12'heee;
rom[102503] = 12'hfff;
rom[102504] = 12'hfff;
rom[102505] = 12'heee;
rom[102506] = 12'heee;
rom[102507] = 12'heee;
rom[102508] = 12'heee;
rom[102509] = 12'heee;
rom[102510] = 12'heee;
rom[102511] = 12'heee;
rom[102512] = 12'hfff;
rom[102513] = 12'hfff;
rom[102514] = 12'hfff;
rom[102515] = 12'hfff;
rom[102516] = 12'heee;
rom[102517] = 12'heee;
rom[102518] = 12'hfff;
rom[102519] = 12'hfff;
rom[102520] = 12'hfff;
rom[102521] = 12'hfff;
rom[102522] = 12'hfff;
rom[102523] = 12'hfff;
rom[102524] = 12'hfff;
rom[102525] = 12'hfff;
rom[102526] = 12'hfff;
rom[102527] = 12'hfff;
rom[102528] = 12'hfff;
rom[102529] = 12'hfff;
rom[102530] = 12'hfff;
rom[102531] = 12'hfff;
rom[102532] = 12'hfff;
rom[102533] = 12'hfff;
rom[102534] = 12'hfff;
rom[102535] = 12'hfff;
rom[102536] = 12'hfff;
rom[102537] = 12'hfff;
rom[102538] = 12'hfff;
rom[102539] = 12'hfff;
rom[102540] = 12'hfff;
rom[102541] = 12'hfff;
rom[102542] = 12'hfff;
rom[102543] = 12'hfff;
rom[102544] = 12'hfff;
rom[102545] = 12'hfff;
rom[102546] = 12'hfff;
rom[102547] = 12'hfff;
rom[102548] = 12'hfff;
rom[102549] = 12'hfff;
rom[102550] = 12'hfff;
rom[102551] = 12'hfff;
rom[102552] = 12'hfff;
rom[102553] = 12'hfff;
rom[102554] = 12'hfff;
rom[102555] = 12'hfff;
rom[102556] = 12'hfff;
rom[102557] = 12'hfff;
rom[102558] = 12'hfff;
rom[102559] = 12'hfff;
rom[102560] = 12'hfff;
rom[102561] = 12'hfff;
rom[102562] = 12'hfff;
rom[102563] = 12'hfff;
rom[102564] = 12'hfff;
rom[102565] = 12'hfff;
rom[102566] = 12'hfff;
rom[102567] = 12'hfff;
rom[102568] = 12'hfff;
rom[102569] = 12'hfff;
rom[102570] = 12'hfff;
rom[102571] = 12'hfff;
rom[102572] = 12'hfff;
rom[102573] = 12'hfff;
rom[102574] = 12'hfff;
rom[102575] = 12'hfff;
rom[102576] = 12'hfff;
rom[102577] = 12'hfff;
rom[102578] = 12'hfff;
rom[102579] = 12'hfff;
rom[102580] = 12'hfff;
rom[102581] = 12'hfff;
rom[102582] = 12'heee;
rom[102583] = 12'heee;
rom[102584] = 12'heee;
rom[102585] = 12'heee;
rom[102586] = 12'heee;
rom[102587] = 12'heee;
rom[102588] = 12'heee;
rom[102589] = 12'heee;
rom[102590] = 12'heee;
rom[102591] = 12'heee;
rom[102592] = 12'heee;
rom[102593] = 12'heee;
rom[102594] = 12'heee;
rom[102595] = 12'heee;
rom[102596] = 12'heee;
rom[102597] = 12'heee;
rom[102598] = 12'heee;
rom[102599] = 12'heee;
rom[102600] = 12'heee;
rom[102601] = 12'heee;
rom[102602] = 12'heee;
rom[102603] = 12'heee;
rom[102604] = 12'heee;
rom[102605] = 12'heee;
rom[102606] = 12'heee;
rom[102607] = 12'heee;
rom[102608] = 12'heee;
rom[102609] = 12'heee;
rom[102610] = 12'heee;
rom[102611] = 12'heee;
rom[102612] = 12'heee;
rom[102613] = 12'heee;
rom[102614] = 12'heee;
rom[102615] = 12'heee;
rom[102616] = 12'hfff;
rom[102617] = 12'hfff;
rom[102618] = 12'hfff;
rom[102619] = 12'hfff;
rom[102620] = 12'hfff;
rom[102621] = 12'hfff;
rom[102622] = 12'hfff;
rom[102623] = 12'hfff;
rom[102624] = 12'hfff;
rom[102625] = 12'hfff;
rom[102626] = 12'hfff;
rom[102627] = 12'hfff;
rom[102628] = 12'hfff;
rom[102629] = 12'hfff;
rom[102630] = 12'hfff;
rom[102631] = 12'hfff;
rom[102632] = 12'hfff;
rom[102633] = 12'hfff;
rom[102634] = 12'hfff;
rom[102635] = 12'hfff;
rom[102636] = 12'hfff;
rom[102637] = 12'hfff;
rom[102638] = 12'hfff;
rom[102639] = 12'hfff;
rom[102640] = 12'hfff;
rom[102641] = 12'hfff;
rom[102642] = 12'hfff;
rom[102643] = 12'hfff;
rom[102644] = 12'hfff;
rom[102645] = 12'heee;
rom[102646] = 12'heee;
rom[102647] = 12'heee;
rom[102648] = 12'hddd;
rom[102649] = 12'hddd;
rom[102650] = 12'hddd;
rom[102651] = 12'hddd;
rom[102652] = 12'hddd;
rom[102653] = 12'hddd;
rom[102654] = 12'hddd;
rom[102655] = 12'hddd;
rom[102656] = 12'hddd;
rom[102657] = 12'hddd;
rom[102658] = 12'hddd;
rom[102659] = 12'hddd;
rom[102660] = 12'hddd;
rom[102661] = 12'hddd;
rom[102662] = 12'hddd;
rom[102663] = 12'hddd;
rom[102664] = 12'hddd;
rom[102665] = 12'hddd;
rom[102666] = 12'hddd;
rom[102667] = 12'heee;
rom[102668] = 12'hfff;
rom[102669] = 12'hfff;
rom[102670] = 12'hfff;
rom[102671] = 12'hfff;
rom[102672] = 12'hfff;
rom[102673] = 12'hfff;
rom[102674] = 12'hfff;
rom[102675] = 12'heee;
rom[102676] = 12'hddd;
rom[102677] = 12'hbbb;
rom[102678] = 12'haaa;
rom[102679] = 12'hbbb;
rom[102680] = 12'haaa;
rom[102681] = 12'h999;
rom[102682] = 12'h888;
rom[102683] = 12'h888;
rom[102684] = 12'h999;
rom[102685] = 12'haaa;
rom[102686] = 12'hccc;
rom[102687] = 12'hddd;
rom[102688] = 12'heee;
rom[102689] = 12'heee;
rom[102690] = 12'heee;
rom[102691] = 12'heee;
rom[102692] = 12'hddd;
rom[102693] = 12'hbbb;
rom[102694] = 12'haaa;
rom[102695] = 12'h999;
rom[102696] = 12'h888;
rom[102697] = 12'h666;
rom[102698] = 12'h444;
rom[102699] = 12'h333;
rom[102700] = 12'h333;
rom[102701] = 12'h333;
rom[102702] = 12'h333;
rom[102703] = 12'h333;
rom[102704] = 12'h333;
rom[102705] = 12'h333;
rom[102706] = 12'h333;
rom[102707] = 12'h333;
rom[102708] = 12'h222;
rom[102709] = 12'h222;
rom[102710] = 12'h222;
rom[102711] = 12'h333;
rom[102712] = 12'h333;
rom[102713] = 12'h333;
rom[102714] = 12'h333;
rom[102715] = 12'h666;
rom[102716] = 12'haaa;
rom[102717] = 12'hccc;
rom[102718] = 12'hccc;
rom[102719] = 12'hbbb;
rom[102720] = 12'h777;
rom[102721] = 12'h666;
rom[102722] = 12'h666;
rom[102723] = 12'h666;
rom[102724] = 12'h555;
rom[102725] = 12'h444;
rom[102726] = 12'h222;
rom[102727] = 12'h222;
rom[102728] = 12'h222;
rom[102729] = 12'h222;
rom[102730] = 12'h222;
rom[102731] = 12'h222;
rom[102732] = 12'h222;
rom[102733] = 12'h222;
rom[102734] = 12'h222;
rom[102735] = 12'h222;
rom[102736] = 12'h222;
rom[102737] = 12'h222;
rom[102738] = 12'h333;
rom[102739] = 12'h555;
rom[102740] = 12'h888;
rom[102741] = 12'hbbb;
rom[102742] = 12'heee;
rom[102743] = 12'hfff;
rom[102744] = 12'heee;
rom[102745] = 12'hbbb;
rom[102746] = 12'h888;
rom[102747] = 12'h666;
rom[102748] = 12'h444;
rom[102749] = 12'h333;
rom[102750] = 12'h333;
rom[102751] = 12'h333;
rom[102752] = 12'h222;
rom[102753] = 12'h222;
rom[102754] = 12'h111;
rom[102755] = 12'h111;
rom[102756] = 12'h111;
rom[102757] = 12'h111;
rom[102758] = 12'h111;
rom[102759] = 12'h  0;
rom[102760] = 12'h111;
rom[102761] = 12'h111;
rom[102762] = 12'h111;
rom[102763] = 12'h111;
rom[102764] = 12'h  0;
rom[102765] = 12'h  0;
rom[102766] = 12'h  0;
rom[102767] = 12'h  0;
rom[102768] = 12'h  0;
rom[102769] = 12'h  0;
rom[102770] = 12'h  0;
rom[102771] = 12'h  0;
rom[102772] = 12'h  0;
rom[102773] = 12'h  0;
rom[102774] = 12'h  0;
rom[102775] = 12'h  0;
rom[102776] = 12'h  0;
rom[102777] = 12'h  0;
rom[102778] = 12'h  0;
rom[102779] = 12'h  0;
rom[102780] = 12'h  0;
rom[102781] = 12'h  0;
rom[102782] = 12'h  0;
rom[102783] = 12'h  0;
rom[102784] = 12'h  0;
rom[102785] = 12'h  0;
rom[102786] = 12'h  0;
rom[102787] = 12'h  0;
rom[102788] = 12'h  0;
rom[102789] = 12'h111;
rom[102790] = 12'h111;
rom[102791] = 12'h111;
rom[102792] = 12'h111;
rom[102793] = 12'h222;
rom[102794] = 12'h222;
rom[102795] = 12'h111;
rom[102796] = 12'h111;
rom[102797] = 12'h  0;
rom[102798] = 12'h  0;
rom[102799] = 12'h  0;
rom[102800] = 12'hfff;
rom[102801] = 12'hfff;
rom[102802] = 12'hfff;
rom[102803] = 12'hfff;
rom[102804] = 12'hfff;
rom[102805] = 12'hfff;
rom[102806] = 12'hfff;
rom[102807] = 12'hfff;
rom[102808] = 12'hfff;
rom[102809] = 12'hfff;
rom[102810] = 12'hfff;
rom[102811] = 12'hfff;
rom[102812] = 12'hfff;
rom[102813] = 12'hfff;
rom[102814] = 12'hfff;
rom[102815] = 12'hfff;
rom[102816] = 12'hfff;
rom[102817] = 12'hfff;
rom[102818] = 12'hfff;
rom[102819] = 12'hfff;
rom[102820] = 12'hfff;
rom[102821] = 12'hfff;
rom[102822] = 12'hfff;
rom[102823] = 12'hfff;
rom[102824] = 12'hfff;
rom[102825] = 12'hfff;
rom[102826] = 12'hfff;
rom[102827] = 12'hfff;
rom[102828] = 12'hfff;
rom[102829] = 12'hfff;
rom[102830] = 12'hfff;
rom[102831] = 12'hfff;
rom[102832] = 12'hfff;
rom[102833] = 12'hfff;
rom[102834] = 12'hfff;
rom[102835] = 12'hfff;
rom[102836] = 12'hfff;
rom[102837] = 12'hfff;
rom[102838] = 12'hfff;
rom[102839] = 12'hfff;
rom[102840] = 12'hfff;
rom[102841] = 12'hfff;
rom[102842] = 12'hfff;
rom[102843] = 12'hfff;
rom[102844] = 12'hfff;
rom[102845] = 12'hfff;
rom[102846] = 12'hfff;
rom[102847] = 12'hfff;
rom[102848] = 12'hfff;
rom[102849] = 12'hfff;
rom[102850] = 12'hfff;
rom[102851] = 12'hfff;
rom[102852] = 12'hfff;
rom[102853] = 12'hfff;
rom[102854] = 12'hfff;
rom[102855] = 12'hfff;
rom[102856] = 12'hfff;
rom[102857] = 12'hfff;
rom[102858] = 12'hfff;
rom[102859] = 12'hfff;
rom[102860] = 12'hfff;
rom[102861] = 12'hfff;
rom[102862] = 12'heee;
rom[102863] = 12'heee;
rom[102864] = 12'heee;
rom[102865] = 12'heee;
rom[102866] = 12'heee;
rom[102867] = 12'heee;
rom[102868] = 12'heee;
rom[102869] = 12'heee;
rom[102870] = 12'heee;
rom[102871] = 12'hfff;
rom[102872] = 12'hfff;
rom[102873] = 12'hfff;
rom[102874] = 12'hfff;
rom[102875] = 12'heee;
rom[102876] = 12'heee;
rom[102877] = 12'heee;
rom[102878] = 12'heee;
rom[102879] = 12'heee;
rom[102880] = 12'heee;
rom[102881] = 12'heee;
rom[102882] = 12'heee;
rom[102883] = 12'heee;
rom[102884] = 12'heee;
rom[102885] = 12'heee;
rom[102886] = 12'hfff;
rom[102887] = 12'hfff;
rom[102888] = 12'hfff;
rom[102889] = 12'hfff;
rom[102890] = 12'heee;
rom[102891] = 12'heee;
rom[102892] = 12'heee;
rom[102893] = 12'heee;
rom[102894] = 12'heee;
rom[102895] = 12'heee;
rom[102896] = 12'heee;
rom[102897] = 12'heee;
rom[102898] = 12'hddd;
rom[102899] = 12'hddd;
rom[102900] = 12'hddd;
rom[102901] = 12'heee;
rom[102902] = 12'heee;
rom[102903] = 12'hfff;
rom[102904] = 12'heee;
rom[102905] = 12'heee;
rom[102906] = 12'heee;
rom[102907] = 12'hddd;
rom[102908] = 12'heee;
rom[102909] = 12'heee;
rom[102910] = 12'hfff;
rom[102911] = 12'hfff;
rom[102912] = 12'hfff;
rom[102913] = 12'hfff;
rom[102914] = 12'hfff;
rom[102915] = 12'hfff;
rom[102916] = 12'hfff;
rom[102917] = 12'hfff;
rom[102918] = 12'hfff;
rom[102919] = 12'hfff;
rom[102920] = 12'hfff;
rom[102921] = 12'hfff;
rom[102922] = 12'hfff;
rom[102923] = 12'hfff;
rom[102924] = 12'hfff;
rom[102925] = 12'hfff;
rom[102926] = 12'hfff;
rom[102927] = 12'hfff;
rom[102928] = 12'hfff;
rom[102929] = 12'hfff;
rom[102930] = 12'hfff;
rom[102931] = 12'hfff;
rom[102932] = 12'hfff;
rom[102933] = 12'hfff;
rom[102934] = 12'hfff;
rom[102935] = 12'hfff;
rom[102936] = 12'hfff;
rom[102937] = 12'hfff;
rom[102938] = 12'hfff;
rom[102939] = 12'hfff;
rom[102940] = 12'hfff;
rom[102941] = 12'hfff;
rom[102942] = 12'hfff;
rom[102943] = 12'hfff;
rom[102944] = 12'hfff;
rom[102945] = 12'hfff;
rom[102946] = 12'hfff;
rom[102947] = 12'hfff;
rom[102948] = 12'hfff;
rom[102949] = 12'hfff;
rom[102950] = 12'hfff;
rom[102951] = 12'hfff;
rom[102952] = 12'hfff;
rom[102953] = 12'hfff;
rom[102954] = 12'hfff;
rom[102955] = 12'hfff;
rom[102956] = 12'hfff;
rom[102957] = 12'hfff;
rom[102958] = 12'hfff;
rom[102959] = 12'hfff;
rom[102960] = 12'hfff;
rom[102961] = 12'hfff;
rom[102962] = 12'hfff;
rom[102963] = 12'hfff;
rom[102964] = 12'hfff;
rom[102965] = 12'hfff;
rom[102966] = 12'hfff;
rom[102967] = 12'hfff;
rom[102968] = 12'hfff;
rom[102969] = 12'hfff;
rom[102970] = 12'hfff;
rom[102971] = 12'hfff;
rom[102972] = 12'hfff;
rom[102973] = 12'hfff;
rom[102974] = 12'hfff;
rom[102975] = 12'hfff;
rom[102976] = 12'hfff;
rom[102977] = 12'hfff;
rom[102978] = 12'hfff;
rom[102979] = 12'hfff;
rom[102980] = 12'hfff;
rom[102981] = 12'hfff;
rom[102982] = 12'hfff;
rom[102983] = 12'hfff;
rom[102984] = 12'hfff;
rom[102985] = 12'hfff;
rom[102986] = 12'hfff;
rom[102987] = 12'hfff;
rom[102988] = 12'hfff;
rom[102989] = 12'hfff;
rom[102990] = 12'hfff;
rom[102991] = 12'hfff;
rom[102992] = 12'heee;
rom[102993] = 12'heee;
rom[102994] = 12'heee;
rom[102995] = 12'heee;
rom[102996] = 12'heee;
rom[102997] = 12'heee;
rom[102998] = 12'heee;
rom[102999] = 12'heee;
rom[103000] = 12'heee;
rom[103001] = 12'heee;
rom[103002] = 12'heee;
rom[103003] = 12'heee;
rom[103004] = 12'heee;
rom[103005] = 12'heee;
rom[103006] = 12'heee;
rom[103007] = 12'heee;
rom[103008] = 12'hfff;
rom[103009] = 12'hfff;
rom[103010] = 12'heee;
rom[103011] = 12'heee;
rom[103012] = 12'heee;
rom[103013] = 12'heee;
rom[103014] = 12'hfff;
rom[103015] = 12'hfff;
rom[103016] = 12'hfff;
rom[103017] = 12'hfff;
rom[103018] = 12'hfff;
rom[103019] = 12'hfff;
rom[103020] = 12'hfff;
rom[103021] = 12'hfff;
rom[103022] = 12'hfff;
rom[103023] = 12'hfff;
rom[103024] = 12'hfff;
rom[103025] = 12'hfff;
rom[103026] = 12'hfff;
rom[103027] = 12'hfff;
rom[103028] = 12'hfff;
rom[103029] = 12'hfff;
rom[103030] = 12'hfff;
rom[103031] = 12'hfff;
rom[103032] = 12'hfff;
rom[103033] = 12'hfff;
rom[103034] = 12'hfff;
rom[103035] = 12'hfff;
rom[103036] = 12'hfff;
rom[103037] = 12'hfff;
rom[103038] = 12'hfff;
rom[103039] = 12'hfff;
rom[103040] = 12'hfff;
rom[103041] = 12'hfff;
rom[103042] = 12'hfff;
rom[103043] = 12'hfff;
rom[103044] = 12'hfff;
rom[103045] = 12'hfff;
rom[103046] = 12'heee;
rom[103047] = 12'heee;
rom[103048] = 12'heee;
rom[103049] = 12'heee;
rom[103050] = 12'heee;
rom[103051] = 12'heee;
rom[103052] = 12'heee;
rom[103053] = 12'heee;
rom[103054] = 12'heee;
rom[103055] = 12'hddd;
rom[103056] = 12'hddd;
rom[103057] = 12'hddd;
rom[103058] = 12'hddd;
rom[103059] = 12'hddd;
rom[103060] = 12'hddd;
rom[103061] = 12'heee;
rom[103062] = 12'heee;
rom[103063] = 12'heee;
rom[103064] = 12'hfff;
rom[103065] = 12'heee;
rom[103066] = 12'hfff;
rom[103067] = 12'hfff;
rom[103068] = 12'hfff;
rom[103069] = 12'hfff;
rom[103070] = 12'hfff;
rom[103071] = 12'hfff;
rom[103072] = 12'heee;
rom[103073] = 12'heee;
rom[103074] = 12'hddd;
rom[103075] = 12'hccc;
rom[103076] = 12'hddd;
rom[103077] = 12'hccc;
rom[103078] = 12'haaa;
rom[103079] = 12'hbbb;
rom[103080] = 12'haaa;
rom[103081] = 12'h999;
rom[103082] = 12'h888;
rom[103083] = 12'h888;
rom[103084] = 12'h888;
rom[103085] = 12'h999;
rom[103086] = 12'haaa;
rom[103087] = 12'hbbb;
rom[103088] = 12'hddd;
rom[103089] = 12'heee;
rom[103090] = 12'heee;
rom[103091] = 12'heee;
rom[103092] = 12'hddd;
rom[103093] = 12'hddd;
rom[103094] = 12'hbbb;
rom[103095] = 12'haaa;
rom[103096] = 12'h999;
rom[103097] = 12'h777;
rom[103098] = 12'h555;
rom[103099] = 12'h444;
rom[103100] = 12'h333;
rom[103101] = 12'h333;
rom[103102] = 12'h333;
rom[103103] = 12'h222;
rom[103104] = 12'h222;
rom[103105] = 12'h222;
rom[103106] = 12'h222;
rom[103107] = 12'h222;
rom[103108] = 12'h222;
rom[103109] = 12'h222;
rom[103110] = 12'h222;
rom[103111] = 12'h222;
rom[103112] = 12'h333;
rom[103113] = 12'h333;
rom[103114] = 12'h333;
rom[103115] = 12'h444;
rom[103116] = 12'h666;
rom[103117] = 12'h888;
rom[103118] = 12'haaa;
rom[103119] = 12'hbbb;
rom[103120] = 12'haaa;
rom[103121] = 12'h888;
rom[103122] = 12'h777;
rom[103123] = 12'h666;
rom[103124] = 12'h555;
rom[103125] = 12'h444;
rom[103126] = 12'h333;
rom[103127] = 12'h222;
rom[103128] = 12'h222;
rom[103129] = 12'h222;
rom[103130] = 12'h222;
rom[103131] = 12'h222;
rom[103132] = 12'h111;
rom[103133] = 12'h111;
rom[103134] = 12'h222;
rom[103135] = 12'h222;
rom[103136] = 12'h222;
rom[103137] = 12'h222;
rom[103138] = 12'h222;
rom[103139] = 12'h333;
rom[103140] = 12'h555;
rom[103141] = 12'h888;
rom[103142] = 12'hbbb;
rom[103143] = 12'hddd;
rom[103144] = 12'hfff;
rom[103145] = 12'heee;
rom[103146] = 12'hbbb;
rom[103147] = 12'h999;
rom[103148] = 12'h666;
rom[103149] = 12'h555;
rom[103150] = 12'h444;
rom[103151] = 12'h333;
rom[103152] = 12'h222;
rom[103153] = 12'h222;
rom[103154] = 12'h111;
rom[103155] = 12'h111;
rom[103156] = 12'h111;
rom[103157] = 12'h111;
rom[103158] = 12'h111;
rom[103159] = 12'h111;
rom[103160] = 12'h111;
rom[103161] = 12'h111;
rom[103162] = 12'h111;
rom[103163] = 12'h111;
rom[103164] = 12'h  0;
rom[103165] = 12'h  0;
rom[103166] = 12'h  0;
rom[103167] = 12'h  0;
rom[103168] = 12'h  0;
rom[103169] = 12'h  0;
rom[103170] = 12'h  0;
rom[103171] = 12'h  0;
rom[103172] = 12'h  0;
rom[103173] = 12'h  0;
rom[103174] = 12'h  0;
rom[103175] = 12'h  0;
rom[103176] = 12'h  0;
rom[103177] = 12'h  0;
rom[103178] = 12'h  0;
rom[103179] = 12'h  0;
rom[103180] = 12'h  0;
rom[103181] = 12'h  0;
rom[103182] = 12'h  0;
rom[103183] = 12'h  0;
rom[103184] = 12'h  0;
rom[103185] = 12'h  0;
rom[103186] = 12'h  0;
rom[103187] = 12'h  0;
rom[103188] = 12'h  0;
rom[103189] = 12'h  0;
rom[103190] = 12'h111;
rom[103191] = 12'h111;
rom[103192] = 12'h111;
rom[103193] = 12'h111;
rom[103194] = 12'h222;
rom[103195] = 12'h111;
rom[103196] = 12'h111;
rom[103197] = 12'h111;
rom[103198] = 12'h  0;
rom[103199] = 12'h  0;
rom[103200] = 12'hfff;
rom[103201] = 12'hfff;
rom[103202] = 12'hfff;
rom[103203] = 12'hfff;
rom[103204] = 12'hfff;
rom[103205] = 12'hfff;
rom[103206] = 12'hfff;
rom[103207] = 12'hfff;
rom[103208] = 12'hfff;
rom[103209] = 12'hfff;
rom[103210] = 12'hfff;
rom[103211] = 12'hfff;
rom[103212] = 12'hfff;
rom[103213] = 12'hfff;
rom[103214] = 12'hfff;
rom[103215] = 12'hfff;
rom[103216] = 12'hfff;
rom[103217] = 12'hfff;
rom[103218] = 12'hfff;
rom[103219] = 12'hfff;
rom[103220] = 12'hfff;
rom[103221] = 12'hfff;
rom[103222] = 12'hfff;
rom[103223] = 12'hfff;
rom[103224] = 12'hfff;
rom[103225] = 12'hfff;
rom[103226] = 12'hfff;
rom[103227] = 12'hfff;
rom[103228] = 12'hfff;
rom[103229] = 12'hfff;
rom[103230] = 12'hfff;
rom[103231] = 12'hfff;
rom[103232] = 12'hfff;
rom[103233] = 12'hfff;
rom[103234] = 12'hfff;
rom[103235] = 12'hfff;
rom[103236] = 12'hfff;
rom[103237] = 12'hfff;
rom[103238] = 12'hfff;
rom[103239] = 12'hfff;
rom[103240] = 12'hfff;
rom[103241] = 12'hfff;
rom[103242] = 12'hfff;
rom[103243] = 12'hfff;
rom[103244] = 12'hfff;
rom[103245] = 12'hfff;
rom[103246] = 12'hfff;
rom[103247] = 12'hfff;
rom[103248] = 12'hfff;
rom[103249] = 12'hfff;
rom[103250] = 12'hfff;
rom[103251] = 12'hfff;
rom[103252] = 12'hfff;
rom[103253] = 12'hfff;
rom[103254] = 12'hfff;
rom[103255] = 12'hfff;
rom[103256] = 12'hfff;
rom[103257] = 12'hfff;
rom[103258] = 12'hfff;
rom[103259] = 12'hfff;
rom[103260] = 12'hfff;
rom[103261] = 12'heee;
rom[103262] = 12'heee;
rom[103263] = 12'heee;
rom[103264] = 12'heee;
rom[103265] = 12'heee;
rom[103266] = 12'heee;
rom[103267] = 12'heee;
rom[103268] = 12'hfff;
rom[103269] = 12'hfff;
rom[103270] = 12'hfff;
rom[103271] = 12'hfff;
rom[103272] = 12'hfff;
rom[103273] = 12'hfff;
rom[103274] = 12'heee;
rom[103275] = 12'heee;
rom[103276] = 12'heee;
rom[103277] = 12'heee;
rom[103278] = 12'heee;
rom[103279] = 12'heee;
rom[103280] = 12'heee;
rom[103281] = 12'heee;
rom[103282] = 12'heee;
rom[103283] = 12'heee;
rom[103284] = 12'hfff;
rom[103285] = 12'hfff;
rom[103286] = 12'hfff;
rom[103287] = 12'hfff;
rom[103288] = 12'hfff;
rom[103289] = 12'heee;
rom[103290] = 12'heee;
rom[103291] = 12'heee;
rom[103292] = 12'heee;
rom[103293] = 12'heee;
rom[103294] = 12'hddd;
rom[103295] = 12'hddd;
rom[103296] = 12'heee;
rom[103297] = 12'hddd;
rom[103298] = 12'hddd;
rom[103299] = 12'hddd;
rom[103300] = 12'heee;
rom[103301] = 12'heee;
rom[103302] = 12'heee;
rom[103303] = 12'heee;
rom[103304] = 12'heee;
rom[103305] = 12'hddd;
rom[103306] = 12'hddd;
rom[103307] = 12'hddd;
rom[103308] = 12'heee;
rom[103309] = 12'heee;
rom[103310] = 12'hfff;
rom[103311] = 12'hfff;
rom[103312] = 12'hfff;
rom[103313] = 12'heee;
rom[103314] = 12'heee;
rom[103315] = 12'heee;
rom[103316] = 12'hfff;
rom[103317] = 12'hfff;
rom[103318] = 12'hfff;
rom[103319] = 12'hfff;
rom[103320] = 12'hfff;
rom[103321] = 12'hfff;
rom[103322] = 12'hfff;
rom[103323] = 12'hfff;
rom[103324] = 12'hfff;
rom[103325] = 12'hfff;
rom[103326] = 12'hfff;
rom[103327] = 12'hfff;
rom[103328] = 12'hfff;
rom[103329] = 12'hfff;
rom[103330] = 12'hfff;
rom[103331] = 12'hfff;
rom[103332] = 12'hfff;
rom[103333] = 12'hfff;
rom[103334] = 12'hfff;
rom[103335] = 12'hfff;
rom[103336] = 12'hfff;
rom[103337] = 12'hfff;
rom[103338] = 12'hfff;
rom[103339] = 12'hfff;
rom[103340] = 12'hfff;
rom[103341] = 12'hfff;
rom[103342] = 12'hfff;
rom[103343] = 12'hfff;
rom[103344] = 12'hfff;
rom[103345] = 12'hfff;
rom[103346] = 12'hfff;
rom[103347] = 12'hfff;
rom[103348] = 12'hfff;
rom[103349] = 12'hfff;
rom[103350] = 12'hfff;
rom[103351] = 12'hfff;
rom[103352] = 12'hfff;
rom[103353] = 12'hfff;
rom[103354] = 12'hfff;
rom[103355] = 12'hfff;
rom[103356] = 12'hfff;
rom[103357] = 12'hfff;
rom[103358] = 12'hfff;
rom[103359] = 12'hfff;
rom[103360] = 12'hfff;
rom[103361] = 12'hfff;
rom[103362] = 12'hfff;
rom[103363] = 12'hfff;
rom[103364] = 12'hfff;
rom[103365] = 12'hfff;
rom[103366] = 12'hfff;
rom[103367] = 12'hfff;
rom[103368] = 12'hfff;
rom[103369] = 12'hfff;
rom[103370] = 12'hfff;
rom[103371] = 12'hfff;
rom[103372] = 12'hfff;
rom[103373] = 12'hfff;
rom[103374] = 12'hfff;
rom[103375] = 12'hfff;
rom[103376] = 12'hfff;
rom[103377] = 12'hfff;
rom[103378] = 12'hfff;
rom[103379] = 12'hfff;
rom[103380] = 12'hfff;
rom[103381] = 12'hfff;
rom[103382] = 12'hfff;
rom[103383] = 12'hfff;
rom[103384] = 12'hfff;
rom[103385] = 12'hfff;
rom[103386] = 12'hfff;
rom[103387] = 12'hfff;
rom[103388] = 12'hfff;
rom[103389] = 12'hfff;
rom[103390] = 12'hfff;
rom[103391] = 12'hfff;
rom[103392] = 12'hfff;
rom[103393] = 12'hfff;
rom[103394] = 12'heee;
rom[103395] = 12'heee;
rom[103396] = 12'hfff;
rom[103397] = 12'hfff;
rom[103398] = 12'hfff;
rom[103399] = 12'hfff;
rom[103400] = 12'hfff;
rom[103401] = 12'hfff;
rom[103402] = 12'hfff;
rom[103403] = 12'hfff;
rom[103404] = 12'hfff;
rom[103405] = 12'hfff;
rom[103406] = 12'hfff;
rom[103407] = 12'hfff;
rom[103408] = 12'hfff;
rom[103409] = 12'hfff;
rom[103410] = 12'hfff;
rom[103411] = 12'hfff;
rom[103412] = 12'hfff;
rom[103413] = 12'hfff;
rom[103414] = 12'hfff;
rom[103415] = 12'hfff;
rom[103416] = 12'hfff;
rom[103417] = 12'hfff;
rom[103418] = 12'hfff;
rom[103419] = 12'hfff;
rom[103420] = 12'hfff;
rom[103421] = 12'hfff;
rom[103422] = 12'hfff;
rom[103423] = 12'hfff;
rom[103424] = 12'hfff;
rom[103425] = 12'hfff;
rom[103426] = 12'hfff;
rom[103427] = 12'hfff;
rom[103428] = 12'hfff;
rom[103429] = 12'hfff;
rom[103430] = 12'hfff;
rom[103431] = 12'hfff;
rom[103432] = 12'hfff;
rom[103433] = 12'hfff;
rom[103434] = 12'hfff;
rom[103435] = 12'hfff;
rom[103436] = 12'hfff;
rom[103437] = 12'hfff;
rom[103438] = 12'hfff;
rom[103439] = 12'hfff;
rom[103440] = 12'hfff;
rom[103441] = 12'hfff;
rom[103442] = 12'hfff;
rom[103443] = 12'hfff;
rom[103444] = 12'hfff;
rom[103445] = 12'hfff;
rom[103446] = 12'hfff;
rom[103447] = 12'hfff;
rom[103448] = 12'hfff;
rom[103449] = 12'hfff;
rom[103450] = 12'hfff;
rom[103451] = 12'hfff;
rom[103452] = 12'hfff;
rom[103453] = 12'hfff;
rom[103454] = 12'heee;
rom[103455] = 12'heee;
rom[103456] = 12'heee;
rom[103457] = 12'heee;
rom[103458] = 12'heee;
rom[103459] = 12'heee;
rom[103460] = 12'heee;
rom[103461] = 12'heee;
rom[103462] = 12'hfff;
rom[103463] = 12'hfff;
rom[103464] = 12'hfff;
rom[103465] = 12'hfff;
rom[103466] = 12'hfff;
rom[103467] = 12'hfff;
rom[103468] = 12'hfff;
rom[103469] = 12'hfff;
rom[103470] = 12'hfff;
rom[103471] = 12'hfff;
rom[103472] = 12'hddd;
rom[103473] = 12'hddd;
rom[103474] = 12'hbbb;
rom[103475] = 12'hbbb;
rom[103476] = 12'hddd;
rom[103477] = 12'hccc;
rom[103478] = 12'hbbb;
rom[103479] = 12'hbbb;
rom[103480] = 12'hbbb;
rom[103481] = 12'haaa;
rom[103482] = 12'h888;
rom[103483] = 12'h777;
rom[103484] = 12'h777;
rom[103485] = 12'h777;
rom[103486] = 12'h888;
rom[103487] = 12'h999;
rom[103488] = 12'hccc;
rom[103489] = 12'heee;
rom[103490] = 12'hfff;
rom[103491] = 12'heee;
rom[103492] = 12'heee;
rom[103493] = 12'heee;
rom[103494] = 12'hddd;
rom[103495] = 12'hbbb;
rom[103496] = 12'haaa;
rom[103497] = 12'h999;
rom[103498] = 12'h777;
rom[103499] = 12'h555;
rom[103500] = 12'h333;
rom[103501] = 12'h333;
rom[103502] = 12'h222;
rom[103503] = 12'h222;
rom[103504] = 12'h222;
rom[103505] = 12'h222;
rom[103506] = 12'h222;
rom[103507] = 12'h222;
rom[103508] = 12'h222;
rom[103509] = 12'h222;
rom[103510] = 12'h222;
rom[103511] = 12'h222;
rom[103512] = 12'h333;
rom[103513] = 12'h333;
rom[103514] = 12'h333;
rom[103515] = 12'h222;
rom[103516] = 12'h222;
rom[103517] = 12'h444;
rom[103518] = 12'h777;
rom[103519] = 12'haaa;
rom[103520] = 12'hbbb;
rom[103521] = 12'haaa;
rom[103522] = 12'h888;
rom[103523] = 12'h666;
rom[103524] = 12'h555;
rom[103525] = 12'h444;
rom[103526] = 12'h333;
rom[103527] = 12'h333;
rom[103528] = 12'h222;
rom[103529] = 12'h222;
rom[103530] = 12'h222;
rom[103531] = 12'h111;
rom[103532] = 12'h111;
rom[103533] = 12'h111;
rom[103534] = 12'h111;
rom[103535] = 12'h222;
rom[103536] = 12'h222;
rom[103537] = 12'h111;
rom[103538] = 12'h111;
rom[103539] = 12'h111;
rom[103540] = 12'h222;
rom[103541] = 12'h444;
rom[103542] = 12'h777;
rom[103543] = 12'haaa;
rom[103544] = 12'heee;
rom[103545] = 12'hfff;
rom[103546] = 12'hfff;
rom[103547] = 12'hddd;
rom[103548] = 12'haaa;
rom[103549] = 12'h777;
rom[103550] = 12'h555;
rom[103551] = 12'h333;
rom[103552] = 12'h222;
rom[103553] = 12'h222;
rom[103554] = 12'h222;
rom[103555] = 12'h222;
rom[103556] = 12'h111;
rom[103557] = 12'h111;
rom[103558] = 12'h111;
rom[103559] = 12'h222;
rom[103560] = 12'h111;
rom[103561] = 12'h111;
rom[103562] = 12'h111;
rom[103563] = 12'h111;
rom[103564] = 12'h  0;
rom[103565] = 12'h  0;
rom[103566] = 12'h  0;
rom[103567] = 12'h  0;
rom[103568] = 12'h  0;
rom[103569] = 12'h  0;
rom[103570] = 12'h  0;
rom[103571] = 12'h  0;
rom[103572] = 12'h  0;
rom[103573] = 12'h  0;
rom[103574] = 12'h  0;
rom[103575] = 12'h  0;
rom[103576] = 12'h  0;
rom[103577] = 12'h  0;
rom[103578] = 12'h  0;
rom[103579] = 12'h  0;
rom[103580] = 12'h  0;
rom[103581] = 12'h  0;
rom[103582] = 12'h  0;
rom[103583] = 12'h  0;
rom[103584] = 12'h  0;
rom[103585] = 12'h  0;
rom[103586] = 12'h  0;
rom[103587] = 12'h  0;
rom[103588] = 12'h  0;
rom[103589] = 12'h  0;
rom[103590] = 12'h  0;
rom[103591] = 12'h111;
rom[103592] = 12'h111;
rom[103593] = 12'h111;
rom[103594] = 12'h222;
rom[103595] = 12'h222;
rom[103596] = 12'h111;
rom[103597] = 12'h111;
rom[103598] = 12'h  0;
rom[103599] = 12'h  0;
rom[103600] = 12'hfff;
rom[103601] = 12'hfff;
rom[103602] = 12'hfff;
rom[103603] = 12'hfff;
rom[103604] = 12'hfff;
rom[103605] = 12'hfff;
rom[103606] = 12'hfff;
rom[103607] = 12'hfff;
rom[103608] = 12'hfff;
rom[103609] = 12'hfff;
rom[103610] = 12'hfff;
rom[103611] = 12'hfff;
rom[103612] = 12'hfff;
rom[103613] = 12'hfff;
rom[103614] = 12'hfff;
rom[103615] = 12'hfff;
rom[103616] = 12'hfff;
rom[103617] = 12'hfff;
rom[103618] = 12'hfff;
rom[103619] = 12'hfff;
rom[103620] = 12'hfff;
rom[103621] = 12'hfff;
rom[103622] = 12'hfff;
rom[103623] = 12'hfff;
rom[103624] = 12'hfff;
rom[103625] = 12'hfff;
rom[103626] = 12'hfff;
rom[103627] = 12'hfff;
rom[103628] = 12'hfff;
rom[103629] = 12'hfff;
rom[103630] = 12'hfff;
rom[103631] = 12'hfff;
rom[103632] = 12'hfff;
rom[103633] = 12'hfff;
rom[103634] = 12'hfff;
rom[103635] = 12'hfff;
rom[103636] = 12'hfff;
rom[103637] = 12'hfff;
rom[103638] = 12'hfff;
rom[103639] = 12'hfff;
rom[103640] = 12'hfff;
rom[103641] = 12'hfff;
rom[103642] = 12'hfff;
rom[103643] = 12'hfff;
rom[103644] = 12'hfff;
rom[103645] = 12'hfff;
rom[103646] = 12'hfff;
rom[103647] = 12'hfff;
rom[103648] = 12'hfff;
rom[103649] = 12'hfff;
rom[103650] = 12'hfff;
rom[103651] = 12'hfff;
rom[103652] = 12'hfff;
rom[103653] = 12'hfff;
rom[103654] = 12'hfff;
rom[103655] = 12'hfff;
rom[103656] = 12'hfff;
rom[103657] = 12'hfff;
rom[103658] = 12'hfff;
rom[103659] = 12'hfff;
rom[103660] = 12'heee;
rom[103661] = 12'heee;
rom[103662] = 12'heee;
rom[103663] = 12'heee;
rom[103664] = 12'heee;
rom[103665] = 12'heee;
rom[103666] = 12'heee;
rom[103667] = 12'hfff;
rom[103668] = 12'hfff;
rom[103669] = 12'hfff;
rom[103670] = 12'hfff;
rom[103671] = 12'hfff;
rom[103672] = 12'heee;
rom[103673] = 12'heee;
rom[103674] = 12'heee;
rom[103675] = 12'heee;
rom[103676] = 12'heee;
rom[103677] = 12'heee;
rom[103678] = 12'heee;
rom[103679] = 12'heee;
rom[103680] = 12'heee;
rom[103681] = 12'heee;
rom[103682] = 12'heee;
rom[103683] = 12'heee;
rom[103684] = 12'hfff;
rom[103685] = 12'hfff;
rom[103686] = 12'hfff;
rom[103687] = 12'hfff;
rom[103688] = 12'heee;
rom[103689] = 12'heee;
rom[103690] = 12'heee;
rom[103691] = 12'heee;
rom[103692] = 12'hddd;
rom[103693] = 12'hddd;
rom[103694] = 12'hddd;
rom[103695] = 12'hddd;
rom[103696] = 12'hddd;
rom[103697] = 12'hddd;
rom[103698] = 12'hddd;
rom[103699] = 12'heee;
rom[103700] = 12'heee;
rom[103701] = 12'hfff;
rom[103702] = 12'heee;
rom[103703] = 12'hddd;
rom[103704] = 12'hddd;
rom[103705] = 12'hddd;
rom[103706] = 12'hddd;
rom[103707] = 12'heee;
rom[103708] = 12'heee;
rom[103709] = 12'hfff;
rom[103710] = 12'hfff;
rom[103711] = 12'hfff;
rom[103712] = 12'heee;
rom[103713] = 12'heee;
rom[103714] = 12'hddd;
rom[103715] = 12'heee;
rom[103716] = 12'hfff;
rom[103717] = 12'hfff;
rom[103718] = 12'hfff;
rom[103719] = 12'hfff;
rom[103720] = 12'hfff;
rom[103721] = 12'hfff;
rom[103722] = 12'hfff;
rom[103723] = 12'hfff;
rom[103724] = 12'hfff;
rom[103725] = 12'hfff;
rom[103726] = 12'hfff;
rom[103727] = 12'hfff;
rom[103728] = 12'hfff;
rom[103729] = 12'hfff;
rom[103730] = 12'hfff;
rom[103731] = 12'hfff;
rom[103732] = 12'hfff;
rom[103733] = 12'hfff;
rom[103734] = 12'hfff;
rom[103735] = 12'hfff;
rom[103736] = 12'hfff;
rom[103737] = 12'hfff;
rom[103738] = 12'hfff;
rom[103739] = 12'hfff;
rom[103740] = 12'hfff;
rom[103741] = 12'hfff;
rom[103742] = 12'hfff;
rom[103743] = 12'hfff;
rom[103744] = 12'hfff;
rom[103745] = 12'hfff;
rom[103746] = 12'hfff;
rom[103747] = 12'hfff;
rom[103748] = 12'hfff;
rom[103749] = 12'hfff;
rom[103750] = 12'hfff;
rom[103751] = 12'hfff;
rom[103752] = 12'hfff;
rom[103753] = 12'hfff;
rom[103754] = 12'hfff;
rom[103755] = 12'hfff;
rom[103756] = 12'hfff;
rom[103757] = 12'hfff;
rom[103758] = 12'hfff;
rom[103759] = 12'hfff;
rom[103760] = 12'hfff;
rom[103761] = 12'hfff;
rom[103762] = 12'hfff;
rom[103763] = 12'hfff;
rom[103764] = 12'hfff;
rom[103765] = 12'hfff;
rom[103766] = 12'hfff;
rom[103767] = 12'hfff;
rom[103768] = 12'hfff;
rom[103769] = 12'hfff;
rom[103770] = 12'hfff;
rom[103771] = 12'hfff;
rom[103772] = 12'hfff;
rom[103773] = 12'hfff;
rom[103774] = 12'hfff;
rom[103775] = 12'hfff;
rom[103776] = 12'hfff;
rom[103777] = 12'hfff;
rom[103778] = 12'hfff;
rom[103779] = 12'hfff;
rom[103780] = 12'hfff;
rom[103781] = 12'hfff;
rom[103782] = 12'hfff;
rom[103783] = 12'hfff;
rom[103784] = 12'hfff;
rom[103785] = 12'hfff;
rom[103786] = 12'hfff;
rom[103787] = 12'hfff;
rom[103788] = 12'hfff;
rom[103789] = 12'hfff;
rom[103790] = 12'hfff;
rom[103791] = 12'hfff;
rom[103792] = 12'hfff;
rom[103793] = 12'hfff;
rom[103794] = 12'hfff;
rom[103795] = 12'hfff;
rom[103796] = 12'hfff;
rom[103797] = 12'hfff;
rom[103798] = 12'hfff;
rom[103799] = 12'hfff;
rom[103800] = 12'heee;
rom[103801] = 12'heee;
rom[103802] = 12'heee;
rom[103803] = 12'heee;
rom[103804] = 12'heee;
rom[103805] = 12'heee;
rom[103806] = 12'heee;
rom[103807] = 12'heee;
rom[103808] = 12'heee;
rom[103809] = 12'heee;
rom[103810] = 12'heee;
rom[103811] = 12'heee;
rom[103812] = 12'heee;
rom[103813] = 12'heee;
rom[103814] = 12'heee;
rom[103815] = 12'heee;
rom[103816] = 12'heee;
rom[103817] = 12'hfff;
rom[103818] = 12'hfff;
rom[103819] = 12'hfff;
rom[103820] = 12'hfff;
rom[103821] = 12'hfff;
rom[103822] = 12'hfff;
rom[103823] = 12'hfff;
rom[103824] = 12'hfff;
rom[103825] = 12'hfff;
rom[103826] = 12'hfff;
rom[103827] = 12'hfff;
rom[103828] = 12'hfff;
rom[103829] = 12'hfff;
rom[103830] = 12'hfff;
rom[103831] = 12'hfff;
rom[103832] = 12'hfff;
rom[103833] = 12'hfff;
rom[103834] = 12'hfff;
rom[103835] = 12'hfff;
rom[103836] = 12'hfff;
rom[103837] = 12'hfff;
rom[103838] = 12'hfff;
rom[103839] = 12'hfff;
rom[103840] = 12'hfff;
rom[103841] = 12'hfff;
rom[103842] = 12'hfff;
rom[103843] = 12'hfff;
rom[103844] = 12'hfff;
rom[103845] = 12'hfff;
rom[103846] = 12'hfff;
rom[103847] = 12'hfff;
rom[103848] = 12'hfff;
rom[103849] = 12'hfff;
rom[103850] = 12'hfff;
rom[103851] = 12'hfff;
rom[103852] = 12'hfff;
rom[103853] = 12'hfff;
rom[103854] = 12'hfff;
rom[103855] = 12'heee;
rom[103856] = 12'hfff;
rom[103857] = 12'hfff;
rom[103858] = 12'hfff;
rom[103859] = 12'heee;
rom[103860] = 12'hfff;
rom[103861] = 12'hfff;
rom[103862] = 12'hfff;
rom[103863] = 12'hfff;
rom[103864] = 12'hfff;
rom[103865] = 12'hfff;
rom[103866] = 12'hfff;
rom[103867] = 12'hfff;
rom[103868] = 12'hfff;
rom[103869] = 12'heee;
rom[103870] = 12'heee;
rom[103871] = 12'heee;
rom[103872] = 12'hddd;
rom[103873] = 12'hccc;
rom[103874] = 12'hbbb;
rom[103875] = 12'hbbb;
rom[103876] = 12'hddd;
rom[103877] = 12'hddd;
rom[103878] = 12'hccc;
rom[103879] = 12'hccc;
rom[103880] = 12'hccc;
rom[103881] = 12'haaa;
rom[103882] = 12'h888;
rom[103883] = 12'h777;
rom[103884] = 12'h777;
rom[103885] = 12'h777;
rom[103886] = 12'h777;
rom[103887] = 12'h888;
rom[103888] = 12'h999;
rom[103889] = 12'hccc;
rom[103890] = 12'heee;
rom[103891] = 12'hfff;
rom[103892] = 12'heee;
rom[103893] = 12'hddd;
rom[103894] = 12'hddd;
rom[103895] = 12'hddd;
rom[103896] = 12'hbbb;
rom[103897] = 12'haaa;
rom[103898] = 12'h888;
rom[103899] = 12'h666;
rom[103900] = 12'h444;
rom[103901] = 12'h333;
rom[103902] = 12'h333;
rom[103903] = 12'h333;
rom[103904] = 12'h333;
rom[103905] = 12'h222;
rom[103906] = 12'h222;
rom[103907] = 12'h222;
rom[103908] = 12'h333;
rom[103909] = 12'h333;
rom[103910] = 12'h222;
rom[103911] = 12'h222;
rom[103912] = 12'h222;
rom[103913] = 12'h222;
rom[103914] = 12'h333;
rom[103915] = 12'h222;
rom[103916] = 12'h111;
rom[103917] = 12'h222;
rom[103918] = 12'h444;
rom[103919] = 12'h666;
rom[103920] = 12'h999;
rom[103921] = 12'haaa;
rom[103922] = 12'h999;
rom[103923] = 12'h888;
rom[103924] = 12'h666;
rom[103925] = 12'h555;
rom[103926] = 12'h444;
rom[103927] = 12'h222;
rom[103928] = 12'h222;
rom[103929] = 12'h222;
rom[103930] = 12'h111;
rom[103931] = 12'h111;
rom[103932] = 12'h111;
rom[103933] = 12'h111;
rom[103934] = 12'h111;
rom[103935] = 12'h111;
rom[103936] = 12'h111;
rom[103937] = 12'h111;
rom[103938] = 12'h111;
rom[103939] = 12'h111;
rom[103940] = 12'h111;
rom[103941] = 12'h222;
rom[103942] = 12'h444;
rom[103943] = 12'h555;
rom[103944] = 12'h999;
rom[103945] = 12'hccc;
rom[103946] = 12'hfff;
rom[103947] = 12'hfff;
rom[103948] = 12'hddd;
rom[103949] = 12'haaa;
rom[103950] = 12'h777;
rom[103951] = 12'h555;
rom[103952] = 12'h444;
rom[103953] = 12'h333;
rom[103954] = 12'h333;
rom[103955] = 12'h222;
rom[103956] = 12'h222;
rom[103957] = 12'h111;
rom[103958] = 12'h111;
rom[103959] = 12'h111;
rom[103960] = 12'h111;
rom[103961] = 12'h111;
rom[103962] = 12'h111;
rom[103963] = 12'h  0;
rom[103964] = 12'h  0;
rom[103965] = 12'h  0;
rom[103966] = 12'h  0;
rom[103967] = 12'h  0;
rom[103968] = 12'h  0;
rom[103969] = 12'h  0;
rom[103970] = 12'h  0;
rom[103971] = 12'h  0;
rom[103972] = 12'h  0;
rom[103973] = 12'h  0;
rom[103974] = 12'h  0;
rom[103975] = 12'h  0;
rom[103976] = 12'h  0;
rom[103977] = 12'h  0;
rom[103978] = 12'h  0;
rom[103979] = 12'h  0;
rom[103980] = 12'h  0;
rom[103981] = 12'h  0;
rom[103982] = 12'h  0;
rom[103983] = 12'h  0;
rom[103984] = 12'h  0;
rom[103985] = 12'h  0;
rom[103986] = 12'h  0;
rom[103987] = 12'h  0;
rom[103988] = 12'h  0;
rom[103989] = 12'h  0;
rom[103990] = 12'h  0;
rom[103991] = 12'h  0;
rom[103992] = 12'h  0;
rom[103993] = 12'h111;
rom[103994] = 12'h111;
rom[103995] = 12'h222;
rom[103996] = 12'h111;
rom[103997] = 12'h111;
rom[103998] = 12'h  0;
rom[103999] = 12'h  0;
rom[104000] = 12'hfff;
rom[104001] = 12'hfff;
rom[104002] = 12'hfff;
rom[104003] = 12'hfff;
rom[104004] = 12'hfff;
rom[104005] = 12'hfff;
rom[104006] = 12'hfff;
rom[104007] = 12'hfff;
rom[104008] = 12'hfff;
rom[104009] = 12'hfff;
rom[104010] = 12'hfff;
rom[104011] = 12'hfff;
rom[104012] = 12'hfff;
rom[104013] = 12'hfff;
rom[104014] = 12'hfff;
rom[104015] = 12'hfff;
rom[104016] = 12'hfff;
rom[104017] = 12'hfff;
rom[104018] = 12'hfff;
rom[104019] = 12'hfff;
rom[104020] = 12'hfff;
rom[104021] = 12'hfff;
rom[104022] = 12'hfff;
rom[104023] = 12'hfff;
rom[104024] = 12'hfff;
rom[104025] = 12'hfff;
rom[104026] = 12'hfff;
rom[104027] = 12'hfff;
rom[104028] = 12'hfff;
rom[104029] = 12'hfff;
rom[104030] = 12'hfff;
rom[104031] = 12'hfff;
rom[104032] = 12'hfff;
rom[104033] = 12'hfff;
rom[104034] = 12'hfff;
rom[104035] = 12'hfff;
rom[104036] = 12'hfff;
rom[104037] = 12'hfff;
rom[104038] = 12'hfff;
rom[104039] = 12'hfff;
rom[104040] = 12'hfff;
rom[104041] = 12'hfff;
rom[104042] = 12'hfff;
rom[104043] = 12'hfff;
rom[104044] = 12'hfff;
rom[104045] = 12'hfff;
rom[104046] = 12'hfff;
rom[104047] = 12'hfff;
rom[104048] = 12'hfff;
rom[104049] = 12'hfff;
rom[104050] = 12'hfff;
rom[104051] = 12'hfff;
rom[104052] = 12'hfff;
rom[104053] = 12'hfff;
rom[104054] = 12'hfff;
rom[104055] = 12'hfff;
rom[104056] = 12'hfff;
rom[104057] = 12'hfff;
rom[104058] = 12'hfff;
rom[104059] = 12'heee;
rom[104060] = 12'heee;
rom[104061] = 12'heee;
rom[104062] = 12'heee;
rom[104063] = 12'heee;
rom[104064] = 12'heee;
rom[104065] = 12'heee;
rom[104066] = 12'heee;
rom[104067] = 12'hfff;
rom[104068] = 12'hfff;
rom[104069] = 12'hfff;
rom[104070] = 12'hfff;
rom[104071] = 12'hfff;
rom[104072] = 12'heee;
rom[104073] = 12'heee;
rom[104074] = 12'heee;
rom[104075] = 12'heee;
rom[104076] = 12'heee;
rom[104077] = 12'heee;
rom[104078] = 12'heee;
rom[104079] = 12'heee;
rom[104080] = 12'heee;
rom[104081] = 12'heee;
rom[104082] = 12'heee;
rom[104083] = 12'hfff;
rom[104084] = 12'hfff;
rom[104085] = 12'hfff;
rom[104086] = 12'hfff;
rom[104087] = 12'heee;
rom[104088] = 12'heee;
rom[104089] = 12'heee;
rom[104090] = 12'hddd;
rom[104091] = 12'hddd;
rom[104092] = 12'hddd;
rom[104093] = 12'hddd;
rom[104094] = 12'hddd;
rom[104095] = 12'hddd;
rom[104096] = 12'hddd;
rom[104097] = 12'hddd;
rom[104098] = 12'hddd;
rom[104099] = 12'heee;
rom[104100] = 12'hfff;
rom[104101] = 12'heee;
rom[104102] = 12'heee;
rom[104103] = 12'hddd;
rom[104104] = 12'hddd;
rom[104105] = 12'hddd;
rom[104106] = 12'heee;
rom[104107] = 12'heee;
rom[104108] = 12'heee;
rom[104109] = 12'heee;
rom[104110] = 12'heee;
rom[104111] = 12'heee;
rom[104112] = 12'heee;
rom[104113] = 12'heee;
rom[104114] = 12'heee;
rom[104115] = 12'heee;
rom[104116] = 12'heee;
rom[104117] = 12'hfff;
rom[104118] = 12'hfff;
rom[104119] = 12'hfff;
rom[104120] = 12'hfff;
rom[104121] = 12'hfff;
rom[104122] = 12'hfff;
rom[104123] = 12'heee;
rom[104124] = 12'heee;
rom[104125] = 12'heee;
rom[104126] = 12'heee;
rom[104127] = 12'heee;
rom[104128] = 12'hfff;
rom[104129] = 12'hfff;
rom[104130] = 12'hfff;
rom[104131] = 12'hfff;
rom[104132] = 12'hfff;
rom[104133] = 12'hfff;
rom[104134] = 12'hfff;
rom[104135] = 12'hfff;
rom[104136] = 12'hfff;
rom[104137] = 12'hfff;
rom[104138] = 12'hfff;
rom[104139] = 12'hfff;
rom[104140] = 12'hfff;
rom[104141] = 12'hfff;
rom[104142] = 12'hfff;
rom[104143] = 12'hfff;
rom[104144] = 12'hfff;
rom[104145] = 12'hfff;
rom[104146] = 12'hfff;
rom[104147] = 12'hfff;
rom[104148] = 12'hfff;
rom[104149] = 12'hfff;
rom[104150] = 12'hfff;
rom[104151] = 12'hfff;
rom[104152] = 12'hfff;
rom[104153] = 12'hfff;
rom[104154] = 12'hfff;
rom[104155] = 12'hfff;
rom[104156] = 12'hfff;
rom[104157] = 12'hfff;
rom[104158] = 12'hfff;
rom[104159] = 12'hfff;
rom[104160] = 12'hfff;
rom[104161] = 12'hfff;
rom[104162] = 12'hfff;
rom[104163] = 12'hfff;
rom[104164] = 12'hfff;
rom[104165] = 12'hfff;
rom[104166] = 12'hfff;
rom[104167] = 12'hfff;
rom[104168] = 12'hfff;
rom[104169] = 12'hfff;
rom[104170] = 12'heee;
rom[104171] = 12'heee;
rom[104172] = 12'heee;
rom[104173] = 12'heee;
rom[104174] = 12'heee;
rom[104175] = 12'heee;
rom[104176] = 12'heee;
rom[104177] = 12'heee;
rom[104178] = 12'heee;
rom[104179] = 12'heee;
rom[104180] = 12'heee;
rom[104181] = 12'heee;
rom[104182] = 12'heee;
rom[104183] = 12'heee;
rom[104184] = 12'heee;
rom[104185] = 12'heee;
rom[104186] = 12'heee;
rom[104187] = 12'heee;
rom[104188] = 12'heee;
rom[104189] = 12'heee;
rom[104190] = 12'heee;
rom[104191] = 12'heee;
rom[104192] = 12'heee;
rom[104193] = 12'heee;
rom[104194] = 12'heee;
rom[104195] = 12'heee;
rom[104196] = 12'heee;
rom[104197] = 12'heee;
rom[104198] = 12'heee;
rom[104199] = 12'heee;
rom[104200] = 12'hddd;
rom[104201] = 12'hddd;
rom[104202] = 12'hddd;
rom[104203] = 12'hddd;
rom[104204] = 12'hddd;
rom[104205] = 12'hddd;
rom[104206] = 12'hddd;
rom[104207] = 12'hddd;
rom[104208] = 12'hddd;
rom[104209] = 12'hddd;
rom[104210] = 12'hddd;
rom[104211] = 12'hddd;
rom[104212] = 12'hddd;
rom[104213] = 12'hddd;
rom[104214] = 12'hddd;
rom[104215] = 12'hddd;
rom[104216] = 12'heee;
rom[104217] = 12'heee;
rom[104218] = 12'heee;
rom[104219] = 12'heee;
rom[104220] = 12'hfff;
rom[104221] = 12'hfff;
rom[104222] = 12'hfff;
rom[104223] = 12'hfff;
rom[104224] = 12'hfff;
rom[104225] = 12'hfff;
rom[104226] = 12'hfff;
rom[104227] = 12'hfff;
rom[104228] = 12'hfff;
rom[104229] = 12'hfff;
rom[104230] = 12'hfff;
rom[104231] = 12'hfff;
rom[104232] = 12'hfff;
rom[104233] = 12'hfff;
rom[104234] = 12'hfff;
rom[104235] = 12'hfff;
rom[104236] = 12'hfff;
rom[104237] = 12'hfff;
rom[104238] = 12'hfff;
rom[104239] = 12'hfff;
rom[104240] = 12'hfff;
rom[104241] = 12'hfff;
rom[104242] = 12'hfff;
rom[104243] = 12'hfff;
rom[104244] = 12'hfff;
rom[104245] = 12'hfff;
rom[104246] = 12'hfff;
rom[104247] = 12'hfff;
rom[104248] = 12'hfff;
rom[104249] = 12'hfff;
rom[104250] = 12'hfff;
rom[104251] = 12'hfff;
rom[104252] = 12'hfff;
rom[104253] = 12'hfff;
rom[104254] = 12'hfff;
rom[104255] = 12'hfff;
rom[104256] = 12'hfff;
rom[104257] = 12'hfff;
rom[104258] = 12'hfff;
rom[104259] = 12'hfff;
rom[104260] = 12'hfff;
rom[104261] = 12'hfff;
rom[104262] = 12'hfff;
rom[104263] = 12'hfff;
rom[104264] = 12'hfff;
rom[104265] = 12'hfff;
rom[104266] = 12'hfff;
rom[104267] = 12'hfff;
rom[104268] = 12'heee;
rom[104269] = 12'heee;
rom[104270] = 12'hddd;
rom[104271] = 12'hddd;
rom[104272] = 12'hccc;
rom[104273] = 12'hbbb;
rom[104274] = 12'haaa;
rom[104275] = 12'hbbb;
rom[104276] = 12'hccc;
rom[104277] = 12'hccc;
rom[104278] = 12'hddd;
rom[104279] = 12'hddd;
rom[104280] = 12'hccc;
rom[104281] = 12'haaa;
rom[104282] = 12'h888;
rom[104283] = 12'h888;
rom[104284] = 12'h777;
rom[104285] = 12'h777;
rom[104286] = 12'h666;
rom[104287] = 12'h666;
rom[104288] = 12'h777;
rom[104289] = 12'h999;
rom[104290] = 12'hccc;
rom[104291] = 12'heee;
rom[104292] = 12'heee;
rom[104293] = 12'heee;
rom[104294] = 12'heee;
rom[104295] = 12'heee;
rom[104296] = 12'hccc;
rom[104297] = 12'hbbb;
rom[104298] = 12'haaa;
rom[104299] = 12'h777;
rom[104300] = 12'h555;
rom[104301] = 12'h333;
rom[104302] = 12'h333;
rom[104303] = 12'h222;
rom[104304] = 12'h333;
rom[104305] = 12'h222;
rom[104306] = 12'h222;
rom[104307] = 12'h222;
rom[104308] = 12'h222;
rom[104309] = 12'h333;
rom[104310] = 12'h333;
rom[104311] = 12'h222;
rom[104312] = 12'h111;
rom[104313] = 12'h222;
rom[104314] = 12'h222;
rom[104315] = 12'h222;
rom[104316] = 12'h222;
rom[104317] = 12'h222;
rom[104318] = 12'h333;
rom[104319] = 12'h333;
rom[104320] = 12'h666;
rom[104321] = 12'h888;
rom[104322] = 12'h999;
rom[104323] = 12'h999;
rom[104324] = 12'h777;
rom[104325] = 12'h666;
rom[104326] = 12'h444;
rom[104327] = 12'h333;
rom[104328] = 12'h222;
rom[104329] = 12'h222;
rom[104330] = 12'h111;
rom[104331] = 12'h111;
rom[104332] = 12'h111;
rom[104333] = 12'h111;
rom[104334] = 12'h111;
rom[104335] = 12'h  0;
rom[104336] = 12'h111;
rom[104337] = 12'h111;
rom[104338] = 12'h111;
rom[104339] = 12'h111;
rom[104340] = 12'h111;
rom[104341] = 12'h111;
rom[104342] = 12'h222;
rom[104343] = 12'h222;
rom[104344] = 12'h444;
rom[104345] = 12'h888;
rom[104346] = 12'hccc;
rom[104347] = 12'heee;
rom[104348] = 12'hfff;
rom[104349] = 12'heee;
rom[104350] = 12'hbbb;
rom[104351] = 12'h888;
rom[104352] = 12'h555;
rom[104353] = 12'h444;
rom[104354] = 12'h333;
rom[104355] = 12'h222;
rom[104356] = 12'h222;
rom[104357] = 12'h222;
rom[104358] = 12'h111;
rom[104359] = 12'h111;
rom[104360] = 12'h111;
rom[104361] = 12'h111;
rom[104362] = 12'h111;
rom[104363] = 12'h111;
rom[104364] = 12'h  0;
rom[104365] = 12'h  0;
rom[104366] = 12'h  0;
rom[104367] = 12'h  0;
rom[104368] = 12'h  0;
rom[104369] = 12'h  0;
rom[104370] = 12'h  0;
rom[104371] = 12'h  0;
rom[104372] = 12'h  0;
rom[104373] = 12'h  0;
rom[104374] = 12'h  0;
rom[104375] = 12'h  0;
rom[104376] = 12'h  0;
rom[104377] = 12'h  0;
rom[104378] = 12'h  0;
rom[104379] = 12'h  0;
rom[104380] = 12'h  0;
rom[104381] = 12'h  0;
rom[104382] = 12'h  0;
rom[104383] = 12'h  0;
rom[104384] = 12'h  0;
rom[104385] = 12'h  0;
rom[104386] = 12'h  0;
rom[104387] = 12'h  0;
rom[104388] = 12'h  0;
rom[104389] = 12'h  0;
rom[104390] = 12'h  0;
rom[104391] = 12'h  0;
rom[104392] = 12'h  0;
rom[104393] = 12'h111;
rom[104394] = 12'h111;
rom[104395] = 12'h111;
rom[104396] = 12'h111;
rom[104397] = 12'h111;
rom[104398] = 12'h111;
rom[104399] = 12'h  0;
rom[104400] = 12'hfff;
rom[104401] = 12'hfff;
rom[104402] = 12'hfff;
rom[104403] = 12'hfff;
rom[104404] = 12'hfff;
rom[104405] = 12'hfff;
rom[104406] = 12'hfff;
rom[104407] = 12'hfff;
rom[104408] = 12'hfff;
rom[104409] = 12'hfff;
rom[104410] = 12'hfff;
rom[104411] = 12'hfff;
rom[104412] = 12'hfff;
rom[104413] = 12'hfff;
rom[104414] = 12'hfff;
rom[104415] = 12'hfff;
rom[104416] = 12'hfff;
rom[104417] = 12'hfff;
rom[104418] = 12'hfff;
rom[104419] = 12'hfff;
rom[104420] = 12'hfff;
rom[104421] = 12'hfff;
rom[104422] = 12'hfff;
rom[104423] = 12'hfff;
rom[104424] = 12'hfff;
rom[104425] = 12'hfff;
rom[104426] = 12'hfff;
rom[104427] = 12'hfff;
rom[104428] = 12'hfff;
rom[104429] = 12'hfff;
rom[104430] = 12'hfff;
rom[104431] = 12'hfff;
rom[104432] = 12'hfff;
rom[104433] = 12'hfff;
rom[104434] = 12'hfff;
rom[104435] = 12'hfff;
rom[104436] = 12'hfff;
rom[104437] = 12'hfff;
rom[104438] = 12'hfff;
rom[104439] = 12'hfff;
rom[104440] = 12'hfff;
rom[104441] = 12'hfff;
rom[104442] = 12'hfff;
rom[104443] = 12'hfff;
rom[104444] = 12'hfff;
rom[104445] = 12'hfff;
rom[104446] = 12'hfff;
rom[104447] = 12'hfff;
rom[104448] = 12'hfff;
rom[104449] = 12'hfff;
rom[104450] = 12'hfff;
rom[104451] = 12'hfff;
rom[104452] = 12'hfff;
rom[104453] = 12'hfff;
rom[104454] = 12'hfff;
rom[104455] = 12'hfff;
rom[104456] = 12'hfff;
rom[104457] = 12'hfff;
rom[104458] = 12'hfff;
rom[104459] = 12'heee;
rom[104460] = 12'heee;
rom[104461] = 12'heee;
rom[104462] = 12'heee;
rom[104463] = 12'heee;
rom[104464] = 12'heee;
rom[104465] = 12'heee;
rom[104466] = 12'heee;
rom[104467] = 12'hfff;
rom[104468] = 12'hfff;
rom[104469] = 12'hfff;
rom[104470] = 12'heee;
rom[104471] = 12'heee;
rom[104472] = 12'heee;
rom[104473] = 12'heee;
rom[104474] = 12'heee;
rom[104475] = 12'heee;
rom[104476] = 12'heee;
rom[104477] = 12'heee;
rom[104478] = 12'heee;
rom[104479] = 12'heee;
rom[104480] = 12'heee;
rom[104481] = 12'heee;
rom[104482] = 12'hfff;
rom[104483] = 12'hfff;
rom[104484] = 12'hfff;
rom[104485] = 12'heee;
rom[104486] = 12'heee;
rom[104487] = 12'heee;
rom[104488] = 12'heee;
rom[104489] = 12'hddd;
rom[104490] = 12'hddd;
rom[104491] = 12'hddd;
rom[104492] = 12'hddd;
rom[104493] = 12'hddd;
rom[104494] = 12'hddd;
rom[104495] = 12'hddd;
rom[104496] = 12'hddd;
rom[104497] = 12'hddd;
rom[104498] = 12'heee;
rom[104499] = 12'heee;
rom[104500] = 12'heee;
rom[104501] = 12'heee;
rom[104502] = 12'hddd;
rom[104503] = 12'hddd;
rom[104504] = 12'hddd;
rom[104505] = 12'hddd;
rom[104506] = 12'heee;
rom[104507] = 12'heee;
rom[104508] = 12'heee;
rom[104509] = 12'heee;
rom[104510] = 12'heee;
rom[104511] = 12'hddd;
rom[104512] = 12'heee;
rom[104513] = 12'heee;
rom[104514] = 12'heee;
rom[104515] = 12'heee;
rom[104516] = 12'heee;
rom[104517] = 12'heee;
rom[104518] = 12'hfff;
rom[104519] = 12'hfff;
rom[104520] = 12'hfff;
rom[104521] = 12'heee;
rom[104522] = 12'heee;
rom[104523] = 12'heee;
rom[104524] = 12'heee;
rom[104525] = 12'heee;
rom[104526] = 12'heee;
rom[104527] = 12'heee;
rom[104528] = 12'heee;
rom[104529] = 12'heee;
rom[104530] = 12'heee;
rom[104531] = 12'heee;
rom[104532] = 12'hfff;
rom[104533] = 12'hfff;
rom[104534] = 12'hfff;
rom[104535] = 12'hfff;
rom[104536] = 12'hfff;
rom[104537] = 12'hfff;
rom[104538] = 12'hfff;
rom[104539] = 12'hfff;
rom[104540] = 12'hfff;
rom[104541] = 12'hfff;
rom[104542] = 12'hfff;
rom[104543] = 12'hfff;
rom[104544] = 12'hfff;
rom[104545] = 12'hfff;
rom[104546] = 12'hfff;
rom[104547] = 12'hfff;
rom[104548] = 12'hfff;
rom[104549] = 12'hfff;
rom[104550] = 12'hfff;
rom[104551] = 12'hfff;
rom[104552] = 12'hfff;
rom[104553] = 12'hfff;
rom[104554] = 12'hfff;
rom[104555] = 12'hfff;
rom[104556] = 12'hfff;
rom[104557] = 12'hfff;
rom[104558] = 12'hfff;
rom[104559] = 12'hfff;
rom[104560] = 12'hfff;
rom[104561] = 12'hfff;
rom[104562] = 12'hfff;
rom[104563] = 12'hfff;
rom[104564] = 12'heee;
rom[104565] = 12'heee;
rom[104566] = 12'heee;
rom[104567] = 12'heee;
rom[104568] = 12'heee;
rom[104569] = 12'heee;
rom[104570] = 12'heee;
rom[104571] = 12'heee;
rom[104572] = 12'heee;
rom[104573] = 12'heee;
rom[104574] = 12'heee;
rom[104575] = 12'heee;
rom[104576] = 12'heee;
rom[104577] = 12'heee;
rom[104578] = 12'heee;
rom[104579] = 12'heee;
rom[104580] = 12'heee;
rom[104581] = 12'heee;
rom[104582] = 12'heee;
rom[104583] = 12'heee;
rom[104584] = 12'heee;
rom[104585] = 12'heee;
rom[104586] = 12'heee;
rom[104587] = 12'heee;
rom[104588] = 12'heee;
rom[104589] = 12'heee;
rom[104590] = 12'heee;
rom[104591] = 12'heee;
rom[104592] = 12'heee;
rom[104593] = 12'heee;
rom[104594] = 12'hddd;
rom[104595] = 12'hddd;
rom[104596] = 12'hddd;
rom[104597] = 12'hddd;
rom[104598] = 12'hddd;
rom[104599] = 12'hddd;
rom[104600] = 12'hccc;
rom[104601] = 12'hccc;
rom[104602] = 12'hccc;
rom[104603] = 12'hccc;
rom[104604] = 12'hccc;
rom[104605] = 12'hccc;
rom[104606] = 12'hccc;
rom[104607] = 12'hccc;
rom[104608] = 12'hccc;
rom[104609] = 12'hccc;
rom[104610] = 12'hccc;
rom[104611] = 12'hccc;
rom[104612] = 12'hccc;
rom[104613] = 12'hccc;
rom[104614] = 12'hccc;
rom[104615] = 12'hddd;
rom[104616] = 12'hddd;
rom[104617] = 12'hddd;
rom[104618] = 12'hddd;
rom[104619] = 12'heee;
rom[104620] = 12'heee;
rom[104621] = 12'heee;
rom[104622] = 12'hfff;
rom[104623] = 12'hfff;
rom[104624] = 12'hfff;
rom[104625] = 12'hfff;
rom[104626] = 12'hfff;
rom[104627] = 12'hfff;
rom[104628] = 12'hfff;
rom[104629] = 12'hfff;
rom[104630] = 12'hfff;
rom[104631] = 12'hfff;
rom[104632] = 12'hfff;
rom[104633] = 12'hfff;
rom[104634] = 12'hfff;
rom[104635] = 12'hfff;
rom[104636] = 12'hfff;
rom[104637] = 12'hfff;
rom[104638] = 12'hfff;
rom[104639] = 12'hfff;
rom[104640] = 12'hfff;
rom[104641] = 12'hfff;
rom[104642] = 12'hfff;
rom[104643] = 12'hfff;
rom[104644] = 12'hfff;
rom[104645] = 12'hfff;
rom[104646] = 12'hfff;
rom[104647] = 12'hfff;
rom[104648] = 12'hfff;
rom[104649] = 12'hfff;
rom[104650] = 12'hfff;
rom[104651] = 12'hfff;
rom[104652] = 12'hfff;
rom[104653] = 12'hfff;
rom[104654] = 12'hfff;
rom[104655] = 12'hfff;
rom[104656] = 12'hfff;
rom[104657] = 12'hfff;
rom[104658] = 12'hfff;
rom[104659] = 12'hfff;
rom[104660] = 12'hfff;
rom[104661] = 12'hfff;
rom[104662] = 12'hfff;
rom[104663] = 12'hfff;
rom[104664] = 12'hfff;
rom[104665] = 12'hfff;
rom[104666] = 12'hfff;
rom[104667] = 12'heee;
rom[104668] = 12'hddd;
rom[104669] = 12'hddd;
rom[104670] = 12'hddd;
rom[104671] = 12'hccc;
rom[104672] = 12'hbbb;
rom[104673] = 12'haaa;
rom[104674] = 12'haaa;
rom[104675] = 12'haaa;
rom[104676] = 12'haaa;
rom[104677] = 12'hbbb;
rom[104678] = 12'hddd;
rom[104679] = 12'hddd;
rom[104680] = 12'hccc;
rom[104681] = 12'hbbb;
rom[104682] = 12'h999;
rom[104683] = 12'h888;
rom[104684] = 12'h777;
rom[104685] = 12'h666;
rom[104686] = 12'h666;
rom[104687] = 12'h555;
rom[104688] = 12'h666;
rom[104689] = 12'h666;
rom[104690] = 12'h888;
rom[104691] = 12'hbbb;
rom[104692] = 12'heee;
rom[104693] = 12'hfff;
rom[104694] = 12'heee;
rom[104695] = 12'hddd;
rom[104696] = 12'hddd;
rom[104697] = 12'hddd;
rom[104698] = 12'hbbb;
rom[104699] = 12'h999;
rom[104700] = 12'h666;
rom[104701] = 12'h444;
rom[104702] = 12'h333;
rom[104703] = 12'h222;
rom[104704] = 12'h333;
rom[104705] = 12'h222;
rom[104706] = 12'h222;
rom[104707] = 12'h222;
rom[104708] = 12'h222;
rom[104709] = 12'h222;
rom[104710] = 12'h222;
rom[104711] = 12'h222;
rom[104712] = 12'h222;
rom[104713] = 12'h222;
rom[104714] = 12'h222;
rom[104715] = 12'h222;
rom[104716] = 12'h222;
rom[104717] = 12'h222;
rom[104718] = 12'h222;
rom[104719] = 12'h222;
rom[104720] = 12'h333;
rom[104721] = 12'h666;
rom[104722] = 12'h888;
rom[104723] = 12'h888;
rom[104724] = 12'h888;
rom[104725] = 12'h777;
rom[104726] = 12'h666;
rom[104727] = 12'h444;
rom[104728] = 12'h222;
rom[104729] = 12'h222;
rom[104730] = 12'h222;
rom[104731] = 12'h111;
rom[104732] = 12'h111;
rom[104733] = 12'h111;
rom[104734] = 12'h111;
rom[104735] = 12'h  0;
rom[104736] = 12'h111;
rom[104737] = 12'h111;
rom[104738] = 12'h111;
rom[104739] = 12'h111;
rom[104740] = 12'h111;
rom[104741] = 12'h111;
rom[104742] = 12'h111;
rom[104743] = 12'h111;
rom[104744] = 12'h333;
rom[104745] = 12'h444;
rom[104746] = 12'h777;
rom[104747] = 12'haaa;
rom[104748] = 12'heee;
rom[104749] = 12'hfff;
rom[104750] = 12'hfff;
rom[104751] = 12'hccc;
rom[104752] = 12'h777;
rom[104753] = 12'h666;
rom[104754] = 12'h444;
rom[104755] = 12'h333;
rom[104756] = 12'h333;
rom[104757] = 12'h333;
rom[104758] = 12'h222;
rom[104759] = 12'h111;
rom[104760] = 12'h111;
rom[104761] = 12'h111;
rom[104762] = 12'h111;
rom[104763] = 12'h111;
rom[104764] = 12'h  0;
rom[104765] = 12'h  0;
rom[104766] = 12'h  0;
rom[104767] = 12'h  0;
rom[104768] = 12'h  0;
rom[104769] = 12'h  0;
rom[104770] = 12'h  0;
rom[104771] = 12'h  0;
rom[104772] = 12'h  0;
rom[104773] = 12'h  0;
rom[104774] = 12'h  0;
rom[104775] = 12'h  0;
rom[104776] = 12'h  0;
rom[104777] = 12'h  0;
rom[104778] = 12'h  0;
rom[104779] = 12'h  0;
rom[104780] = 12'h  0;
rom[104781] = 12'h  0;
rom[104782] = 12'h  0;
rom[104783] = 12'h  0;
rom[104784] = 12'h  0;
rom[104785] = 12'h  0;
rom[104786] = 12'h  0;
rom[104787] = 12'h  0;
rom[104788] = 12'h  0;
rom[104789] = 12'h  0;
rom[104790] = 12'h  0;
rom[104791] = 12'h  0;
rom[104792] = 12'h  0;
rom[104793] = 12'h  0;
rom[104794] = 12'h111;
rom[104795] = 12'h111;
rom[104796] = 12'h111;
rom[104797] = 12'h111;
rom[104798] = 12'h111;
rom[104799] = 12'h111;
rom[104800] = 12'hfff;
rom[104801] = 12'hfff;
rom[104802] = 12'hfff;
rom[104803] = 12'hfff;
rom[104804] = 12'hfff;
rom[104805] = 12'hfff;
rom[104806] = 12'hfff;
rom[104807] = 12'hfff;
rom[104808] = 12'hfff;
rom[104809] = 12'hfff;
rom[104810] = 12'hfff;
rom[104811] = 12'hfff;
rom[104812] = 12'hfff;
rom[104813] = 12'hfff;
rom[104814] = 12'hfff;
rom[104815] = 12'hfff;
rom[104816] = 12'hfff;
rom[104817] = 12'hfff;
rom[104818] = 12'hfff;
rom[104819] = 12'hfff;
rom[104820] = 12'hfff;
rom[104821] = 12'hfff;
rom[104822] = 12'hfff;
rom[104823] = 12'hfff;
rom[104824] = 12'hfff;
rom[104825] = 12'hfff;
rom[104826] = 12'hfff;
rom[104827] = 12'hfff;
rom[104828] = 12'hfff;
rom[104829] = 12'hfff;
rom[104830] = 12'hfff;
rom[104831] = 12'hfff;
rom[104832] = 12'hfff;
rom[104833] = 12'hfff;
rom[104834] = 12'hfff;
rom[104835] = 12'hfff;
rom[104836] = 12'hfff;
rom[104837] = 12'hfff;
rom[104838] = 12'hfff;
rom[104839] = 12'hfff;
rom[104840] = 12'hfff;
rom[104841] = 12'hfff;
rom[104842] = 12'hfff;
rom[104843] = 12'hfff;
rom[104844] = 12'hfff;
rom[104845] = 12'hfff;
rom[104846] = 12'hfff;
rom[104847] = 12'hfff;
rom[104848] = 12'hfff;
rom[104849] = 12'hfff;
rom[104850] = 12'hfff;
rom[104851] = 12'hfff;
rom[104852] = 12'hfff;
rom[104853] = 12'hfff;
rom[104854] = 12'hfff;
rom[104855] = 12'hfff;
rom[104856] = 12'hfff;
rom[104857] = 12'hfff;
rom[104858] = 12'hfff;
rom[104859] = 12'hfff;
rom[104860] = 12'heee;
rom[104861] = 12'heee;
rom[104862] = 12'heee;
rom[104863] = 12'heee;
rom[104864] = 12'heee;
rom[104865] = 12'heee;
rom[104866] = 12'heee;
rom[104867] = 12'hfff;
rom[104868] = 12'heee;
rom[104869] = 12'heee;
rom[104870] = 12'heee;
rom[104871] = 12'heee;
rom[104872] = 12'heee;
rom[104873] = 12'heee;
rom[104874] = 12'heee;
rom[104875] = 12'heee;
rom[104876] = 12'heee;
rom[104877] = 12'heee;
rom[104878] = 12'heee;
rom[104879] = 12'heee;
rom[104880] = 12'hfff;
rom[104881] = 12'hfff;
rom[104882] = 12'hfff;
rom[104883] = 12'hfff;
rom[104884] = 12'heee;
rom[104885] = 12'heee;
rom[104886] = 12'heee;
rom[104887] = 12'hddd;
rom[104888] = 12'hddd;
rom[104889] = 12'hddd;
rom[104890] = 12'hddd;
rom[104891] = 12'hddd;
rom[104892] = 12'hddd;
rom[104893] = 12'hddd;
rom[104894] = 12'hddd;
rom[104895] = 12'hddd;
rom[104896] = 12'hddd;
rom[104897] = 12'heee;
rom[104898] = 12'heee;
rom[104899] = 12'heee;
rom[104900] = 12'hddd;
rom[104901] = 12'hddd;
rom[104902] = 12'hddd;
rom[104903] = 12'hddd;
rom[104904] = 12'heee;
rom[104905] = 12'heee;
rom[104906] = 12'heee;
rom[104907] = 12'heee;
rom[104908] = 12'heee;
rom[104909] = 12'heee;
rom[104910] = 12'hddd;
rom[104911] = 12'hddd;
rom[104912] = 12'hddd;
rom[104913] = 12'hddd;
rom[104914] = 12'heee;
rom[104915] = 12'heee;
rom[104916] = 12'hfff;
rom[104917] = 12'hfff;
rom[104918] = 12'heee;
rom[104919] = 12'heee;
rom[104920] = 12'heee;
rom[104921] = 12'heee;
rom[104922] = 12'hddd;
rom[104923] = 12'hddd;
rom[104924] = 12'hddd;
rom[104925] = 12'hddd;
rom[104926] = 12'hddd;
rom[104927] = 12'hddd;
rom[104928] = 12'hddd;
rom[104929] = 12'hddd;
rom[104930] = 12'hddd;
rom[104931] = 12'hddd;
rom[104932] = 12'heee;
rom[104933] = 12'heee;
rom[104934] = 12'hfff;
rom[104935] = 12'hfff;
rom[104936] = 12'hfff;
rom[104937] = 12'hfff;
rom[104938] = 12'hfff;
rom[104939] = 12'hfff;
rom[104940] = 12'hfff;
rom[104941] = 12'hfff;
rom[104942] = 12'hfff;
rom[104943] = 12'hfff;
rom[104944] = 12'hfff;
rom[104945] = 12'hfff;
rom[104946] = 12'hfff;
rom[104947] = 12'hfff;
rom[104948] = 12'hfff;
rom[104949] = 12'hfff;
rom[104950] = 12'hfff;
rom[104951] = 12'hfff;
rom[104952] = 12'hfff;
rom[104953] = 12'hfff;
rom[104954] = 12'hfff;
rom[104955] = 12'hfff;
rom[104956] = 12'hfff;
rom[104957] = 12'hfff;
rom[104958] = 12'hfff;
rom[104959] = 12'hfff;
rom[104960] = 12'hfff;
rom[104961] = 12'hfff;
rom[104962] = 12'hfff;
rom[104963] = 12'hfff;
rom[104964] = 12'heee;
rom[104965] = 12'heee;
rom[104966] = 12'heee;
rom[104967] = 12'heee;
rom[104968] = 12'heee;
rom[104969] = 12'heee;
rom[104970] = 12'heee;
rom[104971] = 12'heee;
rom[104972] = 12'heee;
rom[104973] = 12'heee;
rom[104974] = 12'heee;
rom[104975] = 12'heee;
rom[104976] = 12'heee;
rom[104977] = 12'heee;
rom[104978] = 12'heee;
rom[104979] = 12'heee;
rom[104980] = 12'heee;
rom[104981] = 12'heee;
rom[104982] = 12'heee;
rom[104983] = 12'hddd;
rom[104984] = 12'heee;
rom[104985] = 12'hddd;
rom[104986] = 12'hddd;
rom[104987] = 12'hddd;
rom[104988] = 12'hddd;
rom[104989] = 12'hddd;
rom[104990] = 12'hddd;
rom[104991] = 12'hddd;
rom[104992] = 12'hddd;
rom[104993] = 12'hddd;
rom[104994] = 12'hddd;
rom[104995] = 12'hccc;
rom[104996] = 12'hccc;
rom[104997] = 12'hccc;
rom[104998] = 12'hccc;
rom[104999] = 12'hccc;
rom[105000] = 12'hccc;
rom[105001] = 12'hccc;
rom[105002] = 12'hccc;
rom[105003] = 12'hccc;
rom[105004] = 12'hbbb;
rom[105005] = 12'hbbb;
rom[105006] = 12'hbbb;
rom[105007] = 12'hbbb;
rom[105008] = 12'hbbb;
rom[105009] = 12'hbbb;
rom[105010] = 12'hbbb;
rom[105011] = 12'hbbb;
rom[105012] = 12'hbbb;
rom[105013] = 12'hccc;
rom[105014] = 12'hccc;
rom[105015] = 12'hccc;
rom[105016] = 12'hccc;
rom[105017] = 12'hccc;
rom[105018] = 12'hddd;
rom[105019] = 12'hddd;
rom[105020] = 12'hddd;
rom[105021] = 12'heee;
rom[105022] = 12'heee;
rom[105023] = 12'heee;
rom[105024] = 12'heee;
rom[105025] = 12'hfff;
rom[105026] = 12'hfff;
rom[105027] = 12'hfff;
rom[105028] = 12'hfff;
rom[105029] = 12'hfff;
rom[105030] = 12'hfff;
rom[105031] = 12'hfff;
rom[105032] = 12'hfff;
rom[105033] = 12'hfff;
rom[105034] = 12'hfff;
rom[105035] = 12'hfff;
rom[105036] = 12'hfff;
rom[105037] = 12'hfff;
rom[105038] = 12'hfff;
rom[105039] = 12'hfff;
rom[105040] = 12'hfff;
rom[105041] = 12'hfff;
rom[105042] = 12'hfff;
rom[105043] = 12'hfff;
rom[105044] = 12'hfff;
rom[105045] = 12'hfff;
rom[105046] = 12'hfff;
rom[105047] = 12'hfff;
rom[105048] = 12'hfff;
rom[105049] = 12'hfff;
rom[105050] = 12'hfff;
rom[105051] = 12'hfff;
rom[105052] = 12'hfff;
rom[105053] = 12'hfff;
rom[105054] = 12'hfff;
rom[105055] = 12'hfff;
rom[105056] = 12'hfff;
rom[105057] = 12'hfff;
rom[105058] = 12'hfff;
rom[105059] = 12'hfff;
rom[105060] = 12'hfff;
rom[105061] = 12'hfff;
rom[105062] = 12'hfff;
rom[105063] = 12'hfff;
rom[105064] = 12'hfff;
rom[105065] = 12'heee;
rom[105066] = 12'hddd;
rom[105067] = 12'hccc;
rom[105068] = 12'hccc;
rom[105069] = 12'hddd;
rom[105070] = 12'hddd;
rom[105071] = 12'hccc;
rom[105072] = 12'haaa;
rom[105073] = 12'h999;
rom[105074] = 12'h888;
rom[105075] = 12'h999;
rom[105076] = 12'h888;
rom[105077] = 12'haaa;
rom[105078] = 12'hccc;
rom[105079] = 12'hddd;
rom[105080] = 12'hddd;
rom[105081] = 12'hccc;
rom[105082] = 12'hbbb;
rom[105083] = 12'h888;
rom[105084] = 12'h777;
rom[105085] = 12'h666;
rom[105086] = 12'h666;
rom[105087] = 12'h666;
rom[105088] = 12'h666;
rom[105089] = 12'h555;
rom[105090] = 12'h555;
rom[105091] = 12'h888;
rom[105092] = 12'hbbb;
rom[105093] = 12'heee;
rom[105094] = 12'heee;
rom[105095] = 12'hddd;
rom[105096] = 12'hddd;
rom[105097] = 12'hddd;
rom[105098] = 12'hddd;
rom[105099] = 12'hbbb;
rom[105100] = 12'h999;
rom[105101] = 12'h666;
rom[105102] = 12'h444;
rom[105103] = 12'h222;
rom[105104] = 12'h222;
rom[105105] = 12'h222;
rom[105106] = 12'h222;
rom[105107] = 12'h222;
rom[105108] = 12'h222;
rom[105109] = 12'h222;
rom[105110] = 12'h222;
rom[105111] = 12'h222;
rom[105112] = 12'h222;
rom[105113] = 12'h222;
rom[105114] = 12'h222;
rom[105115] = 12'h222;
rom[105116] = 12'h222;
rom[105117] = 12'h222;
rom[105118] = 12'h222;
rom[105119] = 12'h111;
rom[105120] = 12'h222;
rom[105121] = 12'h333;
rom[105122] = 12'h555;
rom[105123] = 12'h666;
rom[105124] = 12'h777;
rom[105125] = 12'h777;
rom[105126] = 12'h666;
rom[105127] = 12'h555;
rom[105128] = 12'h333;
rom[105129] = 12'h333;
rom[105130] = 12'h222;
rom[105131] = 12'h111;
rom[105132] = 12'h111;
rom[105133] = 12'h111;
rom[105134] = 12'h111;
rom[105135] = 12'h111;
rom[105136] = 12'h111;
rom[105137] = 12'h111;
rom[105138] = 12'h111;
rom[105139] = 12'h111;
rom[105140] = 12'h111;
rom[105141] = 12'h111;
rom[105142] = 12'h111;
rom[105143] = 12'h111;
rom[105144] = 12'h222;
rom[105145] = 12'h222;
rom[105146] = 12'h333;
rom[105147] = 12'h666;
rom[105148] = 12'haaa;
rom[105149] = 12'heee;
rom[105150] = 12'hfff;
rom[105151] = 12'heee;
rom[105152] = 12'hbbb;
rom[105153] = 12'h999;
rom[105154] = 12'h666;
rom[105155] = 12'h444;
rom[105156] = 12'h333;
rom[105157] = 12'h333;
rom[105158] = 12'h222;
rom[105159] = 12'h222;
rom[105160] = 12'h111;
rom[105161] = 12'h111;
rom[105162] = 12'h111;
rom[105163] = 12'h111;
rom[105164] = 12'h  0;
rom[105165] = 12'h  0;
rom[105166] = 12'h  0;
rom[105167] = 12'h  0;
rom[105168] = 12'h  0;
rom[105169] = 12'h  0;
rom[105170] = 12'h  0;
rom[105171] = 12'h  0;
rom[105172] = 12'h  0;
rom[105173] = 12'h  0;
rom[105174] = 12'h  0;
rom[105175] = 12'h  0;
rom[105176] = 12'h  0;
rom[105177] = 12'h  0;
rom[105178] = 12'h  0;
rom[105179] = 12'h  0;
rom[105180] = 12'h  0;
rom[105181] = 12'h  0;
rom[105182] = 12'h  0;
rom[105183] = 12'h  0;
rom[105184] = 12'h  0;
rom[105185] = 12'h  0;
rom[105186] = 12'h  0;
rom[105187] = 12'h  0;
rom[105188] = 12'h  0;
rom[105189] = 12'h  0;
rom[105190] = 12'h  0;
rom[105191] = 12'h  0;
rom[105192] = 12'h  0;
rom[105193] = 12'h  0;
rom[105194] = 12'h  0;
rom[105195] = 12'h111;
rom[105196] = 12'h111;
rom[105197] = 12'h111;
rom[105198] = 12'h111;
rom[105199] = 12'h111;
rom[105200] = 12'hfff;
rom[105201] = 12'hfff;
rom[105202] = 12'hfff;
rom[105203] = 12'hfff;
rom[105204] = 12'hfff;
rom[105205] = 12'hfff;
rom[105206] = 12'hfff;
rom[105207] = 12'hfff;
rom[105208] = 12'hfff;
rom[105209] = 12'hfff;
rom[105210] = 12'hfff;
rom[105211] = 12'hfff;
rom[105212] = 12'hfff;
rom[105213] = 12'hfff;
rom[105214] = 12'hfff;
rom[105215] = 12'hfff;
rom[105216] = 12'hfff;
rom[105217] = 12'hfff;
rom[105218] = 12'hfff;
rom[105219] = 12'hfff;
rom[105220] = 12'hfff;
rom[105221] = 12'hfff;
rom[105222] = 12'hfff;
rom[105223] = 12'hfff;
rom[105224] = 12'hfff;
rom[105225] = 12'hfff;
rom[105226] = 12'hfff;
rom[105227] = 12'hfff;
rom[105228] = 12'hfff;
rom[105229] = 12'hfff;
rom[105230] = 12'hfff;
rom[105231] = 12'hfff;
rom[105232] = 12'hfff;
rom[105233] = 12'hfff;
rom[105234] = 12'hfff;
rom[105235] = 12'hfff;
rom[105236] = 12'hfff;
rom[105237] = 12'hfff;
rom[105238] = 12'hfff;
rom[105239] = 12'hfff;
rom[105240] = 12'hfff;
rom[105241] = 12'hfff;
rom[105242] = 12'hfff;
rom[105243] = 12'hfff;
rom[105244] = 12'hfff;
rom[105245] = 12'hfff;
rom[105246] = 12'hfff;
rom[105247] = 12'hfff;
rom[105248] = 12'hfff;
rom[105249] = 12'hfff;
rom[105250] = 12'hfff;
rom[105251] = 12'hfff;
rom[105252] = 12'hfff;
rom[105253] = 12'hfff;
rom[105254] = 12'hfff;
rom[105255] = 12'hfff;
rom[105256] = 12'hfff;
rom[105257] = 12'hfff;
rom[105258] = 12'hfff;
rom[105259] = 12'hfff;
rom[105260] = 12'heee;
rom[105261] = 12'heee;
rom[105262] = 12'heee;
rom[105263] = 12'heee;
rom[105264] = 12'hfff;
rom[105265] = 12'hfff;
rom[105266] = 12'heee;
rom[105267] = 12'heee;
rom[105268] = 12'heee;
rom[105269] = 12'heee;
rom[105270] = 12'heee;
rom[105271] = 12'heee;
rom[105272] = 12'heee;
rom[105273] = 12'heee;
rom[105274] = 12'heee;
rom[105275] = 12'heee;
rom[105276] = 12'heee;
rom[105277] = 12'heee;
rom[105278] = 12'heee;
rom[105279] = 12'heee;
rom[105280] = 12'hfff;
rom[105281] = 12'hfff;
rom[105282] = 12'hfff;
rom[105283] = 12'hfff;
rom[105284] = 12'heee;
rom[105285] = 12'heee;
rom[105286] = 12'hddd;
rom[105287] = 12'hddd;
rom[105288] = 12'hddd;
rom[105289] = 12'hddd;
rom[105290] = 12'hddd;
rom[105291] = 12'hddd;
rom[105292] = 12'hddd;
rom[105293] = 12'hddd;
rom[105294] = 12'hddd;
rom[105295] = 12'hddd;
rom[105296] = 12'heee;
rom[105297] = 12'heee;
rom[105298] = 12'heee;
rom[105299] = 12'hddd;
rom[105300] = 12'hccc;
rom[105301] = 12'hccc;
rom[105302] = 12'hccc;
rom[105303] = 12'hddd;
rom[105304] = 12'heee;
rom[105305] = 12'heee;
rom[105306] = 12'heee;
rom[105307] = 12'heee;
rom[105308] = 12'heee;
rom[105309] = 12'hddd;
rom[105310] = 12'hddd;
rom[105311] = 12'hddd;
rom[105312] = 12'hddd;
rom[105313] = 12'hddd;
rom[105314] = 12'heee;
rom[105315] = 12'heee;
rom[105316] = 12'hfff;
rom[105317] = 12'hfff;
rom[105318] = 12'heee;
rom[105319] = 12'heee;
rom[105320] = 12'hddd;
rom[105321] = 12'hddd;
rom[105322] = 12'hddd;
rom[105323] = 12'hccc;
rom[105324] = 12'hccc;
rom[105325] = 12'hccc;
rom[105326] = 12'hccc;
rom[105327] = 12'hccc;
rom[105328] = 12'hccc;
rom[105329] = 12'hccc;
rom[105330] = 12'hccc;
rom[105331] = 12'hddd;
rom[105332] = 12'hddd;
rom[105333] = 12'heee;
rom[105334] = 12'heee;
rom[105335] = 12'hfff;
rom[105336] = 12'heee;
rom[105337] = 12'hfff;
rom[105338] = 12'hfff;
rom[105339] = 12'hfff;
rom[105340] = 12'hfff;
rom[105341] = 12'hfff;
rom[105342] = 12'hfff;
rom[105343] = 12'hfff;
rom[105344] = 12'hfff;
rom[105345] = 12'hfff;
rom[105346] = 12'hfff;
rom[105347] = 12'hfff;
rom[105348] = 12'hfff;
rom[105349] = 12'hfff;
rom[105350] = 12'hfff;
rom[105351] = 12'hfff;
rom[105352] = 12'hfff;
rom[105353] = 12'hfff;
rom[105354] = 12'hfff;
rom[105355] = 12'hfff;
rom[105356] = 12'hfff;
rom[105357] = 12'hfff;
rom[105358] = 12'hfff;
rom[105359] = 12'hfff;
rom[105360] = 12'hfff;
rom[105361] = 12'hfff;
rom[105362] = 12'hfff;
rom[105363] = 12'hfff;
rom[105364] = 12'heee;
rom[105365] = 12'heee;
rom[105366] = 12'heee;
rom[105367] = 12'heee;
rom[105368] = 12'heee;
rom[105369] = 12'heee;
rom[105370] = 12'heee;
rom[105371] = 12'heee;
rom[105372] = 12'heee;
rom[105373] = 12'heee;
rom[105374] = 12'heee;
rom[105375] = 12'heee;
rom[105376] = 12'heee;
rom[105377] = 12'heee;
rom[105378] = 12'heee;
rom[105379] = 12'heee;
rom[105380] = 12'heee;
rom[105381] = 12'heee;
rom[105382] = 12'heee;
rom[105383] = 12'heee;
rom[105384] = 12'hddd;
rom[105385] = 12'hddd;
rom[105386] = 12'hddd;
rom[105387] = 12'hddd;
rom[105388] = 12'hddd;
rom[105389] = 12'hddd;
rom[105390] = 12'hccc;
rom[105391] = 12'hccc;
rom[105392] = 12'hccc;
rom[105393] = 12'hccc;
rom[105394] = 12'hccc;
rom[105395] = 12'hccc;
rom[105396] = 12'hccc;
rom[105397] = 12'hccc;
rom[105398] = 12'hbbb;
rom[105399] = 12'hbbb;
rom[105400] = 12'hbbb;
rom[105401] = 12'hbbb;
rom[105402] = 12'hbbb;
rom[105403] = 12'hbbb;
rom[105404] = 12'hbbb;
rom[105405] = 12'hbbb;
rom[105406] = 12'hbbb;
rom[105407] = 12'hbbb;
rom[105408] = 12'hbbb;
rom[105409] = 12'hbbb;
rom[105410] = 12'hbbb;
rom[105411] = 12'hbbb;
rom[105412] = 12'hbbb;
rom[105413] = 12'hbbb;
rom[105414] = 12'hbbb;
rom[105415] = 12'hbbb;
rom[105416] = 12'hccc;
rom[105417] = 12'hccc;
rom[105418] = 12'hccc;
rom[105419] = 12'hccc;
rom[105420] = 12'hddd;
rom[105421] = 12'hddd;
rom[105422] = 12'hddd;
rom[105423] = 12'hddd;
rom[105424] = 12'heee;
rom[105425] = 12'heee;
rom[105426] = 12'heee;
rom[105427] = 12'hfff;
rom[105428] = 12'hfff;
rom[105429] = 12'hfff;
rom[105430] = 12'hfff;
rom[105431] = 12'hfff;
rom[105432] = 12'hfff;
rom[105433] = 12'hfff;
rom[105434] = 12'hfff;
rom[105435] = 12'hfff;
rom[105436] = 12'hfff;
rom[105437] = 12'hfff;
rom[105438] = 12'hfff;
rom[105439] = 12'hfff;
rom[105440] = 12'hfff;
rom[105441] = 12'hfff;
rom[105442] = 12'hfff;
rom[105443] = 12'hfff;
rom[105444] = 12'hfff;
rom[105445] = 12'hfff;
rom[105446] = 12'hfff;
rom[105447] = 12'hfff;
rom[105448] = 12'hfff;
rom[105449] = 12'hfff;
rom[105450] = 12'hfff;
rom[105451] = 12'hfff;
rom[105452] = 12'hfff;
rom[105453] = 12'hfff;
rom[105454] = 12'hfff;
rom[105455] = 12'hfff;
rom[105456] = 12'hfff;
rom[105457] = 12'hfff;
rom[105458] = 12'hfff;
rom[105459] = 12'hfff;
rom[105460] = 12'hfff;
rom[105461] = 12'hfff;
rom[105462] = 12'heee;
rom[105463] = 12'heee;
rom[105464] = 12'heee;
rom[105465] = 12'hddd;
rom[105466] = 12'hccc;
rom[105467] = 12'hbbb;
rom[105468] = 12'hbbb;
rom[105469] = 12'hddd;
rom[105470] = 12'hddd;
rom[105471] = 12'hddd;
rom[105472] = 12'haaa;
rom[105473] = 12'h888;
rom[105474] = 12'h777;
rom[105475] = 12'h777;
rom[105476] = 12'h666;
rom[105477] = 12'h888;
rom[105478] = 12'hbbb;
rom[105479] = 12'hddd;
rom[105480] = 12'hddd;
rom[105481] = 12'heee;
rom[105482] = 12'hccc;
rom[105483] = 12'h999;
rom[105484] = 12'h666;
rom[105485] = 12'h666;
rom[105486] = 12'h666;
rom[105487] = 12'h666;
rom[105488] = 12'h555;
rom[105489] = 12'h555;
rom[105490] = 12'h444;
rom[105491] = 12'h555;
rom[105492] = 12'h888;
rom[105493] = 12'hccc;
rom[105494] = 12'heee;
rom[105495] = 12'heee;
rom[105496] = 12'hddd;
rom[105497] = 12'hddd;
rom[105498] = 12'hddd;
rom[105499] = 12'hccc;
rom[105500] = 12'haaa;
rom[105501] = 12'h777;
rom[105502] = 12'h555;
rom[105503] = 12'h333;
rom[105504] = 12'h222;
rom[105505] = 12'h222;
rom[105506] = 12'h222;
rom[105507] = 12'h222;
rom[105508] = 12'h222;
rom[105509] = 12'h222;
rom[105510] = 12'h222;
rom[105511] = 12'h222;
rom[105512] = 12'h222;
rom[105513] = 12'h222;
rom[105514] = 12'h222;
rom[105515] = 12'h222;
rom[105516] = 12'h222;
rom[105517] = 12'h111;
rom[105518] = 12'h111;
rom[105519] = 12'h222;
rom[105520] = 12'h111;
rom[105521] = 12'h222;
rom[105522] = 12'h333;
rom[105523] = 12'h555;
rom[105524] = 12'h777;
rom[105525] = 12'h777;
rom[105526] = 12'h666;
rom[105527] = 12'h555;
rom[105528] = 12'h444;
rom[105529] = 12'h333;
rom[105530] = 12'h222;
rom[105531] = 12'h111;
rom[105532] = 12'h111;
rom[105533] = 12'h111;
rom[105534] = 12'h111;
rom[105535] = 12'h111;
rom[105536] = 12'h111;
rom[105537] = 12'h111;
rom[105538] = 12'h111;
rom[105539] = 12'h111;
rom[105540] = 12'h111;
rom[105541] = 12'h111;
rom[105542] = 12'h111;
rom[105543] = 12'h222;
rom[105544] = 12'h111;
rom[105545] = 12'h222;
rom[105546] = 12'h222;
rom[105547] = 12'h333;
rom[105548] = 12'h666;
rom[105549] = 12'haaa;
rom[105550] = 12'hddd;
rom[105551] = 12'hfff;
rom[105552] = 12'heee;
rom[105553] = 12'hccc;
rom[105554] = 12'h888;
rom[105555] = 12'h555;
rom[105556] = 12'h333;
rom[105557] = 12'h333;
rom[105558] = 12'h222;
rom[105559] = 12'h222;
rom[105560] = 12'h111;
rom[105561] = 12'h111;
rom[105562] = 12'h111;
rom[105563] = 12'h111;
rom[105564] = 12'h111;
rom[105565] = 12'h  0;
rom[105566] = 12'h  0;
rom[105567] = 12'h  0;
rom[105568] = 12'h  0;
rom[105569] = 12'h  0;
rom[105570] = 12'h  0;
rom[105571] = 12'h  0;
rom[105572] = 12'h  0;
rom[105573] = 12'h  0;
rom[105574] = 12'h  0;
rom[105575] = 12'h  0;
rom[105576] = 12'h  0;
rom[105577] = 12'h  0;
rom[105578] = 12'h  0;
rom[105579] = 12'h  0;
rom[105580] = 12'h  0;
rom[105581] = 12'h  0;
rom[105582] = 12'h  0;
rom[105583] = 12'h  0;
rom[105584] = 12'h  0;
rom[105585] = 12'h  0;
rom[105586] = 12'h  0;
rom[105587] = 12'h  0;
rom[105588] = 12'h  0;
rom[105589] = 12'h  0;
rom[105590] = 12'h  0;
rom[105591] = 12'h  0;
rom[105592] = 12'h  0;
rom[105593] = 12'h  0;
rom[105594] = 12'h  0;
rom[105595] = 12'h  0;
rom[105596] = 12'h111;
rom[105597] = 12'h111;
rom[105598] = 12'h111;
rom[105599] = 12'h111;
rom[105600] = 12'hfff;
rom[105601] = 12'hfff;
rom[105602] = 12'hfff;
rom[105603] = 12'hfff;
rom[105604] = 12'hfff;
rom[105605] = 12'hfff;
rom[105606] = 12'hfff;
rom[105607] = 12'hfff;
rom[105608] = 12'hfff;
rom[105609] = 12'hfff;
rom[105610] = 12'hfff;
rom[105611] = 12'hfff;
rom[105612] = 12'hfff;
rom[105613] = 12'hfff;
rom[105614] = 12'hfff;
rom[105615] = 12'hfff;
rom[105616] = 12'hfff;
rom[105617] = 12'hfff;
rom[105618] = 12'hfff;
rom[105619] = 12'hfff;
rom[105620] = 12'hfff;
rom[105621] = 12'hfff;
rom[105622] = 12'hfff;
rom[105623] = 12'hfff;
rom[105624] = 12'hfff;
rom[105625] = 12'hfff;
rom[105626] = 12'hfff;
rom[105627] = 12'hfff;
rom[105628] = 12'hfff;
rom[105629] = 12'hfff;
rom[105630] = 12'hfff;
rom[105631] = 12'hfff;
rom[105632] = 12'hfff;
rom[105633] = 12'hfff;
rom[105634] = 12'hfff;
rom[105635] = 12'hfff;
rom[105636] = 12'hfff;
rom[105637] = 12'hfff;
rom[105638] = 12'hfff;
rom[105639] = 12'hfff;
rom[105640] = 12'hfff;
rom[105641] = 12'hfff;
rom[105642] = 12'hfff;
rom[105643] = 12'hfff;
rom[105644] = 12'hfff;
rom[105645] = 12'hfff;
rom[105646] = 12'hfff;
rom[105647] = 12'hfff;
rom[105648] = 12'hfff;
rom[105649] = 12'hfff;
rom[105650] = 12'hfff;
rom[105651] = 12'hfff;
rom[105652] = 12'hfff;
rom[105653] = 12'hfff;
rom[105654] = 12'hfff;
rom[105655] = 12'heee;
rom[105656] = 12'heee;
rom[105657] = 12'heee;
rom[105658] = 12'heee;
rom[105659] = 12'hfff;
rom[105660] = 12'hfff;
rom[105661] = 12'hfff;
rom[105662] = 12'heee;
rom[105663] = 12'heee;
rom[105664] = 12'hfff;
rom[105665] = 12'hfff;
rom[105666] = 12'hfff;
rom[105667] = 12'hfff;
rom[105668] = 12'heee;
rom[105669] = 12'heee;
rom[105670] = 12'heee;
rom[105671] = 12'heee;
rom[105672] = 12'heee;
rom[105673] = 12'heee;
rom[105674] = 12'heee;
rom[105675] = 12'heee;
rom[105676] = 12'heee;
rom[105677] = 12'heee;
rom[105678] = 12'heee;
rom[105679] = 12'heee;
rom[105680] = 12'hfff;
rom[105681] = 12'hfff;
rom[105682] = 12'heee;
rom[105683] = 12'heee;
rom[105684] = 12'heee;
rom[105685] = 12'hddd;
rom[105686] = 12'hddd;
rom[105687] = 12'hddd;
rom[105688] = 12'hccc;
rom[105689] = 12'hddd;
rom[105690] = 12'hddd;
rom[105691] = 12'hddd;
rom[105692] = 12'hddd;
rom[105693] = 12'hddd;
rom[105694] = 12'hddd;
rom[105695] = 12'hddd;
rom[105696] = 12'hfff;
rom[105697] = 12'heee;
rom[105698] = 12'hddd;
rom[105699] = 12'hccc;
rom[105700] = 12'hccc;
rom[105701] = 12'hccc;
rom[105702] = 12'hddd;
rom[105703] = 12'heee;
rom[105704] = 12'heee;
rom[105705] = 12'heee;
rom[105706] = 12'hddd;
rom[105707] = 12'hddd;
rom[105708] = 12'hddd;
rom[105709] = 12'hccc;
rom[105710] = 12'hccc;
rom[105711] = 12'hccc;
rom[105712] = 12'hddd;
rom[105713] = 12'hddd;
rom[105714] = 12'heee;
rom[105715] = 12'hfff;
rom[105716] = 12'hfff;
rom[105717] = 12'hfff;
rom[105718] = 12'heee;
rom[105719] = 12'hddd;
rom[105720] = 12'hddd;
rom[105721] = 12'hccc;
rom[105722] = 12'hbbb;
rom[105723] = 12'hbbb;
rom[105724] = 12'hccc;
rom[105725] = 12'hccc;
rom[105726] = 12'hccc;
rom[105727] = 12'hccc;
rom[105728] = 12'hbbb;
rom[105729] = 12'hccc;
rom[105730] = 12'hccc;
rom[105731] = 12'hccc;
rom[105732] = 12'hddd;
rom[105733] = 12'heee;
rom[105734] = 12'heee;
rom[105735] = 12'heee;
rom[105736] = 12'heee;
rom[105737] = 12'heee;
rom[105738] = 12'heee;
rom[105739] = 12'heee;
rom[105740] = 12'hfff;
rom[105741] = 12'hfff;
rom[105742] = 12'hfff;
rom[105743] = 12'hfff;
rom[105744] = 12'hfff;
rom[105745] = 12'hfff;
rom[105746] = 12'hfff;
rom[105747] = 12'hfff;
rom[105748] = 12'hfff;
rom[105749] = 12'hfff;
rom[105750] = 12'hfff;
rom[105751] = 12'hfff;
rom[105752] = 12'hfff;
rom[105753] = 12'hfff;
rom[105754] = 12'hfff;
rom[105755] = 12'hfff;
rom[105756] = 12'hfff;
rom[105757] = 12'hfff;
rom[105758] = 12'hfff;
rom[105759] = 12'hfff;
rom[105760] = 12'hfff;
rom[105761] = 12'hfff;
rom[105762] = 12'hfff;
rom[105763] = 12'hfff;
rom[105764] = 12'hfff;
rom[105765] = 12'heee;
rom[105766] = 12'heee;
rom[105767] = 12'heee;
rom[105768] = 12'heee;
rom[105769] = 12'heee;
rom[105770] = 12'heee;
rom[105771] = 12'heee;
rom[105772] = 12'heee;
rom[105773] = 12'heee;
rom[105774] = 12'heee;
rom[105775] = 12'heee;
rom[105776] = 12'heee;
rom[105777] = 12'heee;
rom[105778] = 12'heee;
rom[105779] = 12'heee;
rom[105780] = 12'hddd;
rom[105781] = 12'hddd;
rom[105782] = 12'hddd;
rom[105783] = 12'hddd;
rom[105784] = 12'hddd;
rom[105785] = 12'hddd;
rom[105786] = 12'hddd;
rom[105787] = 12'hddd;
rom[105788] = 12'hccc;
rom[105789] = 12'hccc;
rom[105790] = 12'hccc;
rom[105791] = 12'hccc;
rom[105792] = 12'hccc;
rom[105793] = 12'hccc;
rom[105794] = 12'hccc;
rom[105795] = 12'hccc;
rom[105796] = 12'hccc;
rom[105797] = 12'hbbb;
rom[105798] = 12'hbbb;
rom[105799] = 12'hbbb;
rom[105800] = 12'hbbb;
rom[105801] = 12'hbbb;
rom[105802] = 12'hbbb;
rom[105803] = 12'hbbb;
rom[105804] = 12'hbbb;
rom[105805] = 12'hbbb;
rom[105806] = 12'hbbb;
rom[105807] = 12'hbbb;
rom[105808] = 12'hbbb;
rom[105809] = 12'hbbb;
rom[105810] = 12'hbbb;
rom[105811] = 12'hbbb;
rom[105812] = 12'hbbb;
rom[105813] = 12'hbbb;
rom[105814] = 12'hbbb;
rom[105815] = 12'hbbb;
rom[105816] = 12'hbbb;
rom[105817] = 12'hbbb;
rom[105818] = 12'hccc;
rom[105819] = 12'hccc;
rom[105820] = 12'hccc;
rom[105821] = 12'hddd;
rom[105822] = 12'hddd;
rom[105823] = 12'hddd;
rom[105824] = 12'heee;
rom[105825] = 12'heee;
rom[105826] = 12'heee;
rom[105827] = 12'hfff;
rom[105828] = 12'hfff;
rom[105829] = 12'hfff;
rom[105830] = 12'hfff;
rom[105831] = 12'hfff;
rom[105832] = 12'hfff;
rom[105833] = 12'hfff;
rom[105834] = 12'hfff;
rom[105835] = 12'hfff;
rom[105836] = 12'hfff;
rom[105837] = 12'hfff;
rom[105838] = 12'hfff;
rom[105839] = 12'hfff;
rom[105840] = 12'hfff;
rom[105841] = 12'hfff;
rom[105842] = 12'hfff;
rom[105843] = 12'hfff;
rom[105844] = 12'hfff;
rom[105845] = 12'hfff;
rom[105846] = 12'hfff;
rom[105847] = 12'hfff;
rom[105848] = 12'hfff;
rom[105849] = 12'hfff;
rom[105850] = 12'hfff;
rom[105851] = 12'hfff;
rom[105852] = 12'hfff;
rom[105853] = 12'hfff;
rom[105854] = 12'hfff;
rom[105855] = 12'hfff;
rom[105856] = 12'hfff;
rom[105857] = 12'hfff;
rom[105858] = 12'heee;
rom[105859] = 12'heee;
rom[105860] = 12'heee;
rom[105861] = 12'hddd;
rom[105862] = 12'hddd;
rom[105863] = 12'heee;
rom[105864] = 12'hddd;
rom[105865] = 12'hddd;
rom[105866] = 12'hbbb;
rom[105867] = 12'h999;
rom[105868] = 12'haaa;
rom[105869] = 12'hccc;
rom[105870] = 12'heee;
rom[105871] = 12'hddd;
rom[105872] = 12'haaa;
rom[105873] = 12'h777;
rom[105874] = 12'h555;
rom[105875] = 12'h555;
rom[105876] = 12'h555;
rom[105877] = 12'h666;
rom[105878] = 12'h888;
rom[105879] = 12'hbbb;
rom[105880] = 12'heee;
rom[105881] = 12'heee;
rom[105882] = 12'hddd;
rom[105883] = 12'haaa;
rom[105884] = 12'h777;
rom[105885] = 12'h666;
rom[105886] = 12'h666;
rom[105887] = 12'h666;
rom[105888] = 12'h555;
rom[105889] = 12'h555;
rom[105890] = 12'h555;
rom[105891] = 12'h444;
rom[105892] = 12'h555;
rom[105893] = 12'h888;
rom[105894] = 12'hbbb;
rom[105895] = 12'hfff;
rom[105896] = 12'hddd;
rom[105897] = 12'hddd;
rom[105898] = 12'hccc;
rom[105899] = 12'hddd;
rom[105900] = 12'hccc;
rom[105901] = 12'haaa;
rom[105902] = 12'h777;
rom[105903] = 12'h444;
rom[105904] = 12'h333;
rom[105905] = 12'h333;
rom[105906] = 12'h333;
rom[105907] = 12'h222;
rom[105908] = 12'h222;
rom[105909] = 12'h333;
rom[105910] = 12'h222;
rom[105911] = 12'h222;
rom[105912] = 12'h222;
rom[105913] = 12'h222;
rom[105914] = 12'h222;
rom[105915] = 12'h222;
rom[105916] = 12'h222;
rom[105917] = 12'h111;
rom[105918] = 12'h111;
rom[105919] = 12'h111;
rom[105920] = 12'h111;
rom[105921] = 12'h111;
rom[105922] = 12'h222;
rom[105923] = 12'h333;
rom[105924] = 12'h555;
rom[105925] = 12'h666;
rom[105926] = 12'h666;
rom[105927] = 12'h555;
rom[105928] = 12'h444;
rom[105929] = 12'h444;
rom[105930] = 12'h222;
rom[105931] = 12'h222;
rom[105932] = 12'h111;
rom[105933] = 12'h111;
rom[105934] = 12'h111;
rom[105935] = 12'h111;
rom[105936] = 12'h111;
rom[105937] = 12'h111;
rom[105938] = 12'h111;
rom[105939] = 12'h111;
rom[105940] = 12'h111;
rom[105941] = 12'h111;
rom[105942] = 12'h111;
rom[105943] = 12'h111;
rom[105944] = 12'h111;
rom[105945] = 12'h111;
rom[105946] = 12'h222;
rom[105947] = 12'h222;
rom[105948] = 12'h333;
rom[105949] = 12'h444;
rom[105950] = 12'h888;
rom[105951] = 12'hbbb;
rom[105952] = 12'hfff;
rom[105953] = 12'heee;
rom[105954] = 12'hccc;
rom[105955] = 12'h999;
rom[105956] = 12'h666;
rom[105957] = 12'h444;
rom[105958] = 12'h333;
rom[105959] = 12'h222;
rom[105960] = 12'h222;
rom[105961] = 12'h222;
rom[105962] = 12'h111;
rom[105963] = 12'h111;
rom[105964] = 12'h111;
rom[105965] = 12'h111;
rom[105966] = 12'h111;
rom[105967] = 12'h  0;
rom[105968] = 12'h  0;
rom[105969] = 12'h  0;
rom[105970] = 12'h  0;
rom[105971] = 12'h  0;
rom[105972] = 12'h  0;
rom[105973] = 12'h  0;
rom[105974] = 12'h  0;
rom[105975] = 12'h  0;
rom[105976] = 12'h  0;
rom[105977] = 12'h  0;
rom[105978] = 12'h  0;
rom[105979] = 12'h  0;
rom[105980] = 12'h  0;
rom[105981] = 12'h  0;
rom[105982] = 12'h  0;
rom[105983] = 12'h  0;
rom[105984] = 12'h  0;
rom[105985] = 12'h  0;
rom[105986] = 12'h  0;
rom[105987] = 12'h  0;
rom[105988] = 12'h  0;
rom[105989] = 12'h  0;
rom[105990] = 12'h  0;
rom[105991] = 12'h  0;
rom[105992] = 12'h  0;
rom[105993] = 12'h  0;
rom[105994] = 12'h  0;
rom[105995] = 12'h  0;
rom[105996] = 12'h111;
rom[105997] = 12'h111;
rom[105998] = 12'h111;
rom[105999] = 12'h111;
rom[106000] = 12'hfff;
rom[106001] = 12'hfff;
rom[106002] = 12'hfff;
rom[106003] = 12'hfff;
rom[106004] = 12'hfff;
rom[106005] = 12'hfff;
rom[106006] = 12'hfff;
rom[106007] = 12'hfff;
rom[106008] = 12'hfff;
rom[106009] = 12'hfff;
rom[106010] = 12'hfff;
rom[106011] = 12'hfff;
rom[106012] = 12'hfff;
rom[106013] = 12'hfff;
rom[106014] = 12'hfff;
rom[106015] = 12'hfff;
rom[106016] = 12'hfff;
rom[106017] = 12'hfff;
rom[106018] = 12'hfff;
rom[106019] = 12'hfff;
rom[106020] = 12'hfff;
rom[106021] = 12'hfff;
rom[106022] = 12'hfff;
rom[106023] = 12'hfff;
rom[106024] = 12'hfff;
rom[106025] = 12'hfff;
rom[106026] = 12'hfff;
rom[106027] = 12'hfff;
rom[106028] = 12'hfff;
rom[106029] = 12'hfff;
rom[106030] = 12'hfff;
rom[106031] = 12'hfff;
rom[106032] = 12'hfff;
rom[106033] = 12'hfff;
rom[106034] = 12'hfff;
rom[106035] = 12'hfff;
rom[106036] = 12'hfff;
rom[106037] = 12'hfff;
rom[106038] = 12'hfff;
rom[106039] = 12'hfff;
rom[106040] = 12'hfff;
rom[106041] = 12'hfff;
rom[106042] = 12'hfff;
rom[106043] = 12'hfff;
rom[106044] = 12'hfff;
rom[106045] = 12'hfff;
rom[106046] = 12'hfff;
rom[106047] = 12'hfff;
rom[106048] = 12'hfff;
rom[106049] = 12'hfff;
rom[106050] = 12'hfff;
rom[106051] = 12'hfff;
rom[106052] = 12'hfff;
rom[106053] = 12'hfff;
rom[106054] = 12'hfff;
rom[106055] = 12'heee;
rom[106056] = 12'heee;
rom[106057] = 12'heee;
rom[106058] = 12'heee;
rom[106059] = 12'hfff;
rom[106060] = 12'hfff;
rom[106061] = 12'heee;
rom[106062] = 12'heee;
rom[106063] = 12'heee;
rom[106064] = 12'heee;
rom[106065] = 12'heee;
rom[106066] = 12'heee;
rom[106067] = 12'heee;
rom[106068] = 12'heee;
rom[106069] = 12'heee;
rom[106070] = 12'heee;
rom[106071] = 12'heee;
rom[106072] = 12'heee;
rom[106073] = 12'heee;
rom[106074] = 12'heee;
rom[106075] = 12'heee;
rom[106076] = 12'heee;
rom[106077] = 12'heee;
rom[106078] = 12'heee;
rom[106079] = 12'hfff;
rom[106080] = 12'hfff;
rom[106081] = 12'hfff;
rom[106082] = 12'heee;
rom[106083] = 12'heee;
rom[106084] = 12'hddd;
rom[106085] = 12'hddd;
rom[106086] = 12'hddd;
rom[106087] = 12'hddd;
rom[106088] = 12'hccc;
rom[106089] = 12'hddd;
rom[106090] = 12'hddd;
rom[106091] = 12'hddd;
rom[106092] = 12'hddd;
rom[106093] = 12'hddd;
rom[106094] = 12'hddd;
rom[106095] = 12'heee;
rom[106096] = 12'hfff;
rom[106097] = 12'hddd;
rom[106098] = 12'hccc;
rom[106099] = 12'hccc;
rom[106100] = 12'hccc;
rom[106101] = 12'hddd;
rom[106102] = 12'heee;
rom[106103] = 12'heee;
rom[106104] = 12'heee;
rom[106105] = 12'hddd;
rom[106106] = 12'hccc;
rom[106107] = 12'hccc;
rom[106108] = 12'hccc;
rom[106109] = 12'hccc;
rom[106110] = 12'hccc;
rom[106111] = 12'hccc;
rom[106112] = 12'hddd;
rom[106113] = 12'heee;
rom[106114] = 12'hfff;
rom[106115] = 12'hfff;
rom[106116] = 12'hfff;
rom[106117] = 12'heee;
rom[106118] = 12'hddd;
rom[106119] = 12'hddd;
rom[106120] = 12'hccc;
rom[106121] = 12'hbbb;
rom[106122] = 12'hbbb;
rom[106123] = 12'hbbb;
rom[106124] = 12'hbbb;
rom[106125] = 12'hbbb;
rom[106126] = 12'hbbb;
rom[106127] = 12'hbbb;
rom[106128] = 12'hbbb;
rom[106129] = 12'hccc;
rom[106130] = 12'hccc;
rom[106131] = 12'hddd;
rom[106132] = 12'hddd;
rom[106133] = 12'heee;
rom[106134] = 12'heee;
rom[106135] = 12'hddd;
rom[106136] = 12'hddd;
rom[106137] = 12'hddd;
rom[106138] = 12'hddd;
rom[106139] = 12'hddd;
rom[106140] = 12'heee;
rom[106141] = 12'heee;
rom[106142] = 12'hfff;
rom[106143] = 12'hfff;
rom[106144] = 12'hfff;
rom[106145] = 12'hfff;
rom[106146] = 12'hfff;
rom[106147] = 12'hfff;
rom[106148] = 12'hfff;
rom[106149] = 12'hfff;
rom[106150] = 12'hfff;
rom[106151] = 12'hfff;
rom[106152] = 12'hfff;
rom[106153] = 12'hfff;
rom[106154] = 12'hfff;
rom[106155] = 12'hfff;
rom[106156] = 12'hfff;
rom[106157] = 12'hfff;
rom[106158] = 12'hfff;
rom[106159] = 12'hfff;
rom[106160] = 12'hfff;
rom[106161] = 12'hfff;
rom[106162] = 12'hfff;
rom[106163] = 12'hfff;
rom[106164] = 12'hfff;
rom[106165] = 12'heee;
rom[106166] = 12'heee;
rom[106167] = 12'heee;
rom[106168] = 12'heee;
rom[106169] = 12'heee;
rom[106170] = 12'heee;
rom[106171] = 12'heee;
rom[106172] = 12'heee;
rom[106173] = 12'heee;
rom[106174] = 12'heee;
rom[106175] = 12'heee;
rom[106176] = 12'hddd;
rom[106177] = 12'hddd;
rom[106178] = 12'hddd;
rom[106179] = 12'hddd;
rom[106180] = 12'hddd;
rom[106181] = 12'hddd;
rom[106182] = 12'hddd;
rom[106183] = 12'hddd;
rom[106184] = 12'hddd;
rom[106185] = 12'hddd;
rom[106186] = 12'hccc;
rom[106187] = 12'hccc;
rom[106188] = 12'hccc;
rom[106189] = 12'hccc;
rom[106190] = 12'hccc;
rom[106191] = 12'hccc;
rom[106192] = 12'hccc;
rom[106193] = 12'hccc;
rom[106194] = 12'hccc;
rom[106195] = 12'hccc;
rom[106196] = 12'hccc;
rom[106197] = 12'hbbb;
rom[106198] = 12'hbbb;
rom[106199] = 12'hbbb;
rom[106200] = 12'hbbb;
rom[106201] = 12'hbbb;
rom[106202] = 12'hbbb;
rom[106203] = 12'hbbb;
rom[106204] = 12'hbbb;
rom[106205] = 12'hbbb;
rom[106206] = 12'hbbb;
rom[106207] = 12'hbbb;
rom[106208] = 12'hbbb;
rom[106209] = 12'hbbb;
rom[106210] = 12'hbbb;
rom[106211] = 12'hbbb;
rom[106212] = 12'hbbb;
rom[106213] = 12'hbbb;
rom[106214] = 12'hbbb;
rom[106215] = 12'hbbb;
rom[106216] = 12'hbbb;
rom[106217] = 12'hbbb;
rom[106218] = 12'hccc;
rom[106219] = 12'hccc;
rom[106220] = 12'hccc;
rom[106221] = 12'hddd;
rom[106222] = 12'hddd;
rom[106223] = 12'hddd;
rom[106224] = 12'hddd;
rom[106225] = 12'heee;
rom[106226] = 12'heee;
rom[106227] = 12'heee;
rom[106228] = 12'hfff;
rom[106229] = 12'hfff;
rom[106230] = 12'hfff;
rom[106231] = 12'hfff;
rom[106232] = 12'hfff;
rom[106233] = 12'hfff;
rom[106234] = 12'hfff;
rom[106235] = 12'hfff;
rom[106236] = 12'hfff;
rom[106237] = 12'hfff;
rom[106238] = 12'hfff;
rom[106239] = 12'hfff;
rom[106240] = 12'hfff;
rom[106241] = 12'hfff;
rom[106242] = 12'hfff;
rom[106243] = 12'hfff;
rom[106244] = 12'hfff;
rom[106245] = 12'hfff;
rom[106246] = 12'hfff;
rom[106247] = 12'hfff;
rom[106248] = 12'hfff;
rom[106249] = 12'hfff;
rom[106250] = 12'hfff;
rom[106251] = 12'hfff;
rom[106252] = 12'hfff;
rom[106253] = 12'hfff;
rom[106254] = 12'hfff;
rom[106255] = 12'hfff;
rom[106256] = 12'hfff;
rom[106257] = 12'heee;
rom[106258] = 12'hddd;
rom[106259] = 12'hddd;
rom[106260] = 12'hddd;
rom[106261] = 12'hddd;
rom[106262] = 12'hddd;
rom[106263] = 12'heee;
rom[106264] = 12'heee;
rom[106265] = 12'hddd;
rom[106266] = 12'hbbb;
rom[106267] = 12'h999;
rom[106268] = 12'h999;
rom[106269] = 12'hccc;
rom[106270] = 12'heee;
rom[106271] = 12'hddd;
rom[106272] = 12'haaa;
rom[106273] = 12'h777;
rom[106274] = 12'h555;
rom[106275] = 12'h555;
rom[106276] = 12'h444;
rom[106277] = 12'h444;
rom[106278] = 12'h666;
rom[106279] = 12'h888;
rom[106280] = 12'hccc;
rom[106281] = 12'hddd;
rom[106282] = 12'heee;
rom[106283] = 12'hccc;
rom[106284] = 12'h999;
rom[106285] = 12'h666;
rom[106286] = 12'h555;
rom[106287] = 12'h555;
rom[106288] = 12'h555;
rom[106289] = 12'h555;
rom[106290] = 12'h555;
rom[106291] = 12'h444;
rom[106292] = 12'h444;
rom[106293] = 12'h666;
rom[106294] = 12'h999;
rom[106295] = 12'hccc;
rom[106296] = 12'hddd;
rom[106297] = 12'hddd;
rom[106298] = 12'hccc;
rom[106299] = 12'hddd;
rom[106300] = 12'heee;
rom[106301] = 12'hccc;
rom[106302] = 12'h999;
rom[106303] = 12'h666;
rom[106304] = 12'h444;
rom[106305] = 12'h333;
rom[106306] = 12'h333;
rom[106307] = 12'h222;
rom[106308] = 12'h222;
rom[106309] = 12'h222;
rom[106310] = 12'h222;
rom[106311] = 12'h222;
rom[106312] = 12'h222;
rom[106313] = 12'h222;
rom[106314] = 12'h222;
rom[106315] = 12'h111;
rom[106316] = 12'h111;
rom[106317] = 12'h111;
rom[106318] = 12'h111;
rom[106319] = 12'h111;
rom[106320] = 12'h111;
rom[106321] = 12'h111;
rom[106322] = 12'h111;
rom[106323] = 12'h222;
rom[106324] = 12'h444;
rom[106325] = 12'h555;
rom[106326] = 12'h555;
rom[106327] = 12'h555;
rom[106328] = 12'h555;
rom[106329] = 12'h444;
rom[106330] = 12'h333;
rom[106331] = 12'h222;
rom[106332] = 12'h111;
rom[106333] = 12'h111;
rom[106334] = 12'h111;
rom[106335] = 12'h111;
rom[106336] = 12'h111;
rom[106337] = 12'h111;
rom[106338] = 12'h111;
rom[106339] = 12'h111;
rom[106340] = 12'h111;
rom[106341] = 12'h111;
rom[106342] = 12'h111;
rom[106343] = 12'h111;
rom[106344] = 12'h111;
rom[106345] = 12'h111;
rom[106346] = 12'h111;
rom[106347] = 12'h222;
rom[106348] = 12'h222;
rom[106349] = 12'h333;
rom[106350] = 12'h555;
rom[106351] = 12'h888;
rom[106352] = 12'hddd;
rom[106353] = 12'hddd;
rom[106354] = 12'hddd;
rom[106355] = 12'hbbb;
rom[106356] = 12'h888;
rom[106357] = 12'h666;
rom[106358] = 12'h444;
rom[106359] = 12'h333;
rom[106360] = 12'h222;
rom[106361] = 12'h222;
rom[106362] = 12'h222;
rom[106363] = 12'h111;
rom[106364] = 12'h111;
rom[106365] = 12'h111;
rom[106366] = 12'h111;
rom[106367] = 12'h111;
rom[106368] = 12'h  0;
rom[106369] = 12'h  0;
rom[106370] = 12'h  0;
rom[106371] = 12'h  0;
rom[106372] = 12'h  0;
rom[106373] = 12'h  0;
rom[106374] = 12'h  0;
rom[106375] = 12'h  0;
rom[106376] = 12'h  0;
rom[106377] = 12'h  0;
rom[106378] = 12'h  0;
rom[106379] = 12'h  0;
rom[106380] = 12'h  0;
rom[106381] = 12'h  0;
rom[106382] = 12'h  0;
rom[106383] = 12'h  0;
rom[106384] = 12'h  0;
rom[106385] = 12'h  0;
rom[106386] = 12'h  0;
rom[106387] = 12'h  0;
rom[106388] = 12'h  0;
rom[106389] = 12'h  0;
rom[106390] = 12'h  0;
rom[106391] = 12'h  0;
rom[106392] = 12'h  0;
rom[106393] = 12'h  0;
rom[106394] = 12'h  0;
rom[106395] = 12'h  0;
rom[106396] = 12'h  0;
rom[106397] = 12'h111;
rom[106398] = 12'h111;
rom[106399] = 12'h111;
rom[106400] = 12'hfff;
rom[106401] = 12'hfff;
rom[106402] = 12'hfff;
rom[106403] = 12'hfff;
rom[106404] = 12'hfff;
rom[106405] = 12'hfff;
rom[106406] = 12'hfff;
rom[106407] = 12'hfff;
rom[106408] = 12'hfff;
rom[106409] = 12'hfff;
rom[106410] = 12'hfff;
rom[106411] = 12'hfff;
rom[106412] = 12'hfff;
rom[106413] = 12'hfff;
rom[106414] = 12'hfff;
rom[106415] = 12'hfff;
rom[106416] = 12'hfff;
rom[106417] = 12'hfff;
rom[106418] = 12'hfff;
rom[106419] = 12'hfff;
rom[106420] = 12'hfff;
rom[106421] = 12'hfff;
rom[106422] = 12'hfff;
rom[106423] = 12'hfff;
rom[106424] = 12'hfff;
rom[106425] = 12'hfff;
rom[106426] = 12'hfff;
rom[106427] = 12'hfff;
rom[106428] = 12'hfff;
rom[106429] = 12'hfff;
rom[106430] = 12'hfff;
rom[106431] = 12'hfff;
rom[106432] = 12'hfff;
rom[106433] = 12'hfff;
rom[106434] = 12'hfff;
rom[106435] = 12'hfff;
rom[106436] = 12'hfff;
rom[106437] = 12'hfff;
rom[106438] = 12'hfff;
rom[106439] = 12'hfff;
rom[106440] = 12'hfff;
rom[106441] = 12'hfff;
rom[106442] = 12'hfff;
rom[106443] = 12'hfff;
rom[106444] = 12'hfff;
rom[106445] = 12'hfff;
rom[106446] = 12'hfff;
rom[106447] = 12'hfff;
rom[106448] = 12'hfff;
rom[106449] = 12'hfff;
rom[106450] = 12'hfff;
rom[106451] = 12'hfff;
rom[106452] = 12'hfff;
rom[106453] = 12'hfff;
rom[106454] = 12'hfff;
rom[106455] = 12'heee;
rom[106456] = 12'heee;
rom[106457] = 12'heee;
rom[106458] = 12'heee;
rom[106459] = 12'heee;
rom[106460] = 12'heee;
rom[106461] = 12'heee;
rom[106462] = 12'heee;
rom[106463] = 12'heee;
rom[106464] = 12'heee;
rom[106465] = 12'heee;
rom[106466] = 12'heee;
rom[106467] = 12'heee;
rom[106468] = 12'heee;
rom[106469] = 12'heee;
rom[106470] = 12'heee;
rom[106471] = 12'heee;
rom[106472] = 12'heee;
rom[106473] = 12'heee;
rom[106474] = 12'heee;
rom[106475] = 12'heee;
rom[106476] = 12'heee;
rom[106477] = 12'heee;
rom[106478] = 12'heee;
rom[106479] = 12'hfff;
rom[106480] = 12'hfff;
rom[106481] = 12'heee;
rom[106482] = 12'heee;
rom[106483] = 12'hddd;
rom[106484] = 12'hddd;
rom[106485] = 12'hddd;
rom[106486] = 12'hddd;
rom[106487] = 12'hddd;
rom[106488] = 12'hccc;
rom[106489] = 12'hccc;
rom[106490] = 12'hccc;
rom[106491] = 12'hddd;
rom[106492] = 12'hddd;
rom[106493] = 12'hddd;
rom[106494] = 12'heee;
rom[106495] = 12'hfff;
rom[106496] = 12'heee;
rom[106497] = 12'hddd;
rom[106498] = 12'hbbb;
rom[106499] = 12'hbbb;
rom[106500] = 12'hddd;
rom[106501] = 12'heee;
rom[106502] = 12'heee;
rom[106503] = 12'heee;
rom[106504] = 12'hddd;
rom[106505] = 12'hccc;
rom[106506] = 12'hccc;
rom[106507] = 12'hccc;
rom[106508] = 12'hccc;
rom[106509] = 12'hccc;
rom[106510] = 12'hbbb;
rom[106511] = 12'hbbb;
rom[106512] = 12'hddd;
rom[106513] = 12'hfff;
rom[106514] = 12'hfff;
rom[106515] = 12'hfff;
rom[106516] = 12'heee;
rom[106517] = 12'hddd;
rom[106518] = 12'hccc;
rom[106519] = 12'hccc;
rom[106520] = 12'hbbb;
rom[106521] = 12'haaa;
rom[106522] = 12'haaa;
rom[106523] = 12'haaa;
rom[106524] = 12'haaa;
rom[106525] = 12'haaa;
rom[106526] = 12'haaa;
rom[106527] = 12'haaa;
rom[106528] = 12'hbbb;
rom[106529] = 12'hbbb;
rom[106530] = 12'hccc;
rom[106531] = 12'hddd;
rom[106532] = 12'heee;
rom[106533] = 12'heee;
rom[106534] = 12'hddd;
rom[106535] = 12'hddd;
rom[106536] = 12'hddd;
rom[106537] = 12'hddd;
rom[106538] = 12'hccc;
rom[106539] = 12'hccc;
rom[106540] = 12'hddd;
rom[106541] = 12'hddd;
rom[106542] = 12'heee;
rom[106543] = 12'heee;
rom[106544] = 12'hfff;
rom[106545] = 12'hfff;
rom[106546] = 12'hfff;
rom[106547] = 12'hfff;
rom[106548] = 12'hfff;
rom[106549] = 12'hfff;
rom[106550] = 12'hfff;
rom[106551] = 12'hfff;
rom[106552] = 12'hfff;
rom[106553] = 12'hfff;
rom[106554] = 12'hfff;
rom[106555] = 12'hfff;
rom[106556] = 12'hfff;
rom[106557] = 12'hfff;
rom[106558] = 12'hfff;
rom[106559] = 12'hfff;
rom[106560] = 12'hfff;
rom[106561] = 12'hfff;
rom[106562] = 12'hfff;
rom[106563] = 12'hfff;
rom[106564] = 12'hfff;
rom[106565] = 12'hfff;
rom[106566] = 12'heee;
rom[106567] = 12'heee;
rom[106568] = 12'heee;
rom[106569] = 12'heee;
rom[106570] = 12'heee;
rom[106571] = 12'heee;
rom[106572] = 12'heee;
rom[106573] = 12'heee;
rom[106574] = 12'heee;
rom[106575] = 12'heee;
rom[106576] = 12'hddd;
rom[106577] = 12'hddd;
rom[106578] = 12'hddd;
rom[106579] = 12'hddd;
rom[106580] = 12'hddd;
rom[106581] = 12'hddd;
rom[106582] = 12'hddd;
rom[106583] = 12'hddd;
rom[106584] = 12'hddd;
rom[106585] = 12'hccc;
rom[106586] = 12'hccc;
rom[106587] = 12'hccc;
rom[106588] = 12'hccc;
rom[106589] = 12'hccc;
rom[106590] = 12'hccc;
rom[106591] = 12'hccc;
rom[106592] = 12'hccc;
rom[106593] = 12'hccc;
rom[106594] = 12'hccc;
rom[106595] = 12'hccc;
rom[106596] = 12'hccc;
rom[106597] = 12'hbbb;
rom[106598] = 12'hbbb;
rom[106599] = 12'hbbb;
rom[106600] = 12'hbbb;
rom[106601] = 12'hbbb;
rom[106602] = 12'hbbb;
rom[106603] = 12'hbbb;
rom[106604] = 12'hbbb;
rom[106605] = 12'hbbb;
rom[106606] = 12'hbbb;
rom[106607] = 12'hbbb;
rom[106608] = 12'hbbb;
rom[106609] = 12'hbbb;
rom[106610] = 12'hbbb;
rom[106611] = 12'hbbb;
rom[106612] = 12'hbbb;
rom[106613] = 12'hbbb;
rom[106614] = 12'hbbb;
rom[106615] = 12'hbbb;
rom[106616] = 12'hbbb;
rom[106617] = 12'hccc;
rom[106618] = 12'hccc;
rom[106619] = 12'hccc;
rom[106620] = 12'hddd;
rom[106621] = 12'hddd;
rom[106622] = 12'hddd;
rom[106623] = 12'heee;
rom[106624] = 12'heee;
rom[106625] = 12'heee;
rom[106626] = 12'heee;
rom[106627] = 12'hfff;
rom[106628] = 12'hfff;
rom[106629] = 12'hfff;
rom[106630] = 12'hfff;
rom[106631] = 12'hfff;
rom[106632] = 12'hfff;
rom[106633] = 12'hfff;
rom[106634] = 12'hfff;
rom[106635] = 12'hfff;
rom[106636] = 12'hfff;
rom[106637] = 12'hfff;
rom[106638] = 12'hfff;
rom[106639] = 12'hfff;
rom[106640] = 12'hfff;
rom[106641] = 12'hfff;
rom[106642] = 12'hfff;
rom[106643] = 12'hfff;
rom[106644] = 12'hfff;
rom[106645] = 12'hfff;
rom[106646] = 12'hfff;
rom[106647] = 12'hfff;
rom[106648] = 12'hfff;
rom[106649] = 12'hfff;
rom[106650] = 12'hfff;
rom[106651] = 12'hfff;
rom[106652] = 12'hfff;
rom[106653] = 12'hfff;
rom[106654] = 12'heee;
rom[106655] = 12'heee;
rom[106656] = 12'hddd;
rom[106657] = 12'hccc;
rom[106658] = 12'hccc;
rom[106659] = 12'hccc;
rom[106660] = 12'hccc;
rom[106661] = 12'hddd;
rom[106662] = 12'hddd;
rom[106663] = 12'heee;
rom[106664] = 12'heee;
rom[106665] = 12'hddd;
rom[106666] = 12'hbbb;
rom[106667] = 12'h999;
rom[106668] = 12'h999;
rom[106669] = 12'hbbb;
rom[106670] = 12'hddd;
rom[106671] = 12'heee;
rom[106672] = 12'hbbb;
rom[106673] = 12'h777;
rom[106674] = 12'h555;
rom[106675] = 12'h444;
rom[106676] = 12'h444;
rom[106677] = 12'h333;
rom[106678] = 12'h333;
rom[106679] = 12'h555;
rom[106680] = 12'h999;
rom[106681] = 12'hccc;
rom[106682] = 12'hfff;
rom[106683] = 12'heee;
rom[106684] = 12'haaa;
rom[106685] = 12'h777;
rom[106686] = 12'h555;
rom[106687] = 12'h555;
rom[106688] = 12'h555;
rom[106689] = 12'h555;
rom[106690] = 12'h555;
rom[106691] = 12'h444;
rom[106692] = 12'h333;
rom[106693] = 12'h444;
rom[106694] = 12'h666;
rom[106695] = 12'h888;
rom[106696] = 12'hccc;
rom[106697] = 12'hddd;
rom[106698] = 12'hddd;
rom[106699] = 12'hccc;
rom[106700] = 12'hddd;
rom[106701] = 12'heee;
rom[106702] = 12'hccc;
rom[106703] = 12'h999;
rom[106704] = 12'h555;
rom[106705] = 12'h444;
rom[106706] = 12'h333;
rom[106707] = 12'h333;
rom[106708] = 12'h222;
rom[106709] = 12'h222;
rom[106710] = 12'h222;
rom[106711] = 12'h222;
rom[106712] = 12'h222;
rom[106713] = 12'h111;
rom[106714] = 12'h111;
rom[106715] = 12'h111;
rom[106716] = 12'h111;
rom[106717] = 12'h111;
rom[106718] = 12'h111;
rom[106719] = 12'h111;
rom[106720] = 12'h  0;
rom[106721] = 12'h111;
rom[106722] = 12'h111;
rom[106723] = 12'h222;
rom[106724] = 12'h222;
rom[106725] = 12'h444;
rom[106726] = 12'h555;
rom[106727] = 12'h555;
rom[106728] = 12'h555;
rom[106729] = 12'h444;
rom[106730] = 12'h333;
rom[106731] = 12'h222;
rom[106732] = 12'h111;
rom[106733] = 12'h111;
rom[106734] = 12'h111;
rom[106735] = 12'h111;
rom[106736] = 12'h111;
rom[106737] = 12'h111;
rom[106738] = 12'h111;
rom[106739] = 12'h111;
rom[106740] = 12'h111;
rom[106741] = 12'h111;
rom[106742] = 12'h111;
rom[106743] = 12'h111;
rom[106744] = 12'h111;
rom[106745] = 12'h111;
rom[106746] = 12'h111;
rom[106747] = 12'h111;
rom[106748] = 12'h111;
rom[106749] = 12'h111;
rom[106750] = 12'h333;
rom[106751] = 12'h444;
rom[106752] = 12'h999;
rom[106753] = 12'hbbb;
rom[106754] = 12'heee;
rom[106755] = 12'heee;
rom[106756] = 12'hbbb;
rom[106757] = 12'h888;
rom[106758] = 12'h555;
rom[106759] = 12'h333;
rom[106760] = 12'h333;
rom[106761] = 12'h222;
rom[106762] = 12'h222;
rom[106763] = 12'h111;
rom[106764] = 12'h111;
rom[106765] = 12'h111;
rom[106766] = 12'h111;
rom[106767] = 12'h111;
rom[106768] = 12'h111;
rom[106769] = 12'h  0;
rom[106770] = 12'h  0;
rom[106771] = 12'h  0;
rom[106772] = 12'h  0;
rom[106773] = 12'h  0;
rom[106774] = 12'h  0;
rom[106775] = 12'h  0;
rom[106776] = 12'h  0;
rom[106777] = 12'h  0;
rom[106778] = 12'h  0;
rom[106779] = 12'h  0;
rom[106780] = 12'h  0;
rom[106781] = 12'h  0;
rom[106782] = 12'h  0;
rom[106783] = 12'h  0;
rom[106784] = 12'h  0;
rom[106785] = 12'h  0;
rom[106786] = 12'h  0;
rom[106787] = 12'h  0;
rom[106788] = 12'h  0;
rom[106789] = 12'h  0;
rom[106790] = 12'h  0;
rom[106791] = 12'h  0;
rom[106792] = 12'h  0;
rom[106793] = 12'h  0;
rom[106794] = 12'h  0;
rom[106795] = 12'h  0;
rom[106796] = 12'h  0;
rom[106797] = 12'h111;
rom[106798] = 12'h111;
rom[106799] = 12'h111;
rom[106800] = 12'hfff;
rom[106801] = 12'hfff;
rom[106802] = 12'hfff;
rom[106803] = 12'hfff;
rom[106804] = 12'hfff;
rom[106805] = 12'hfff;
rom[106806] = 12'hfff;
rom[106807] = 12'hfff;
rom[106808] = 12'hfff;
rom[106809] = 12'hfff;
rom[106810] = 12'hfff;
rom[106811] = 12'hfff;
rom[106812] = 12'hfff;
rom[106813] = 12'hfff;
rom[106814] = 12'hfff;
rom[106815] = 12'hfff;
rom[106816] = 12'hfff;
rom[106817] = 12'hfff;
rom[106818] = 12'hfff;
rom[106819] = 12'hfff;
rom[106820] = 12'hfff;
rom[106821] = 12'hfff;
rom[106822] = 12'hfff;
rom[106823] = 12'hfff;
rom[106824] = 12'hfff;
rom[106825] = 12'hfff;
rom[106826] = 12'hfff;
rom[106827] = 12'hfff;
rom[106828] = 12'hfff;
rom[106829] = 12'hfff;
rom[106830] = 12'hfff;
rom[106831] = 12'hfff;
rom[106832] = 12'hfff;
rom[106833] = 12'hfff;
rom[106834] = 12'hfff;
rom[106835] = 12'hfff;
rom[106836] = 12'hfff;
rom[106837] = 12'hfff;
rom[106838] = 12'hfff;
rom[106839] = 12'hfff;
rom[106840] = 12'hfff;
rom[106841] = 12'hfff;
rom[106842] = 12'hfff;
rom[106843] = 12'hfff;
rom[106844] = 12'hfff;
rom[106845] = 12'hfff;
rom[106846] = 12'hfff;
rom[106847] = 12'hfff;
rom[106848] = 12'hfff;
rom[106849] = 12'hfff;
rom[106850] = 12'hfff;
rom[106851] = 12'hfff;
rom[106852] = 12'hfff;
rom[106853] = 12'hfff;
rom[106854] = 12'heee;
rom[106855] = 12'heee;
rom[106856] = 12'heee;
rom[106857] = 12'heee;
rom[106858] = 12'heee;
rom[106859] = 12'heee;
rom[106860] = 12'heee;
rom[106861] = 12'heee;
rom[106862] = 12'heee;
rom[106863] = 12'heee;
rom[106864] = 12'heee;
rom[106865] = 12'heee;
rom[106866] = 12'heee;
rom[106867] = 12'heee;
rom[106868] = 12'heee;
rom[106869] = 12'heee;
rom[106870] = 12'heee;
rom[106871] = 12'heee;
rom[106872] = 12'heee;
rom[106873] = 12'heee;
rom[106874] = 12'heee;
rom[106875] = 12'heee;
rom[106876] = 12'heee;
rom[106877] = 12'heee;
rom[106878] = 12'heee;
rom[106879] = 12'hfff;
rom[106880] = 12'heee;
rom[106881] = 12'heee;
rom[106882] = 12'hddd;
rom[106883] = 12'hddd;
rom[106884] = 12'hccc;
rom[106885] = 12'hccc;
rom[106886] = 12'hccc;
rom[106887] = 12'hccc;
rom[106888] = 12'hccc;
rom[106889] = 12'hccc;
rom[106890] = 12'hccc;
rom[106891] = 12'hddd;
rom[106892] = 12'heee;
rom[106893] = 12'heee;
rom[106894] = 12'heee;
rom[106895] = 12'heee;
rom[106896] = 12'hddd;
rom[106897] = 12'hccc;
rom[106898] = 12'hccc;
rom[106899] = 12'hccc;
rom[106900] = 12'heee;
rom[106901] = 12'heee;
rom[106902] = 12'heee;
rom[106903] = 12'hddd;
rom[106904] = 12'hccc;
rom[106905] = 12'hccc;
rom[106906] = 12'hbbb;
rom[106907] = 12'hccc;
rom[106908] = 12'hccc;
rom[106909] = 12'hbbb;
rom[106910] = 12'hbbb;
rom[106911] = 12'hbbb;
rom[106912] = 12'heee;
rom[106913] = 12'hfff;
rom[106914] = 12'hfff;
rom[106915] = 12'heee;
rom[106916] = 12'hccc;
rom[106917] = 12'hbbb;
rom[106918] = 12'hbbb;
rom[106919] = 12'hbbb;
rom[106920] = 12'haaa;
rom[106921] = 12'haaa;
rom[106922] = 12'haaa;
rom[106923] = 12'haaa;
rom[106924] = 12'haaa;
rom[106925] = 12'haaa;
rom[106926] = 12'haaa;
rom[106927] = 12'haaa;
rom[106928] = 12'hbbb;
rom[106929] = 12'hbbb;
rom[106930] = 12'hccc;
rom[106931] = 12'heee;
rom[106932] = 12'heee;
rom[106933] = 12'hddd;
rom[106934] = 12'hccc;
rom[106935] = 12'hccc;
rom[106936] = 12'hccc;
rom[106937] = 12'hccc;
rom[106938] = 12'hccc;
rom[106939] = 12'hccc;
rom[106940] = 12'hccc;
rom[106941] = 12'hddd;
rom[106942] = 12'hddd;
rom[106943] = 12'heee;
rom[106944] = 12'heee;
rom[106945] = 12'heee;
rom[106946] = 12'hfff;
rom[106947] = 12'hfff;
rom[106948] = 12'hfff;
rom[106949] = 12'hfff;
rom[106950] = 12'hfff;
rom[106951] = 12'hfff;
rom[106952] = 12'hfff;
rom[106953] = 12'hfff;
rom[106954] = 12'hfff;
rom[106955] = 12'hfff;
rom[106956] = 12'hfff;
rom[106957] = 12'hfff;
rom[106958] = 12'hfff;
rom[106959] = 12'hfff;
rom[106960] = 12'hfff;
rom[106961] = 12'hfff;
rom[106962] = 12'hfff;
rom[106963] = 12'hfff;
rom[106964] = 12'hfff;
rom[106965] = 12'hfff;
rom[106966] = 12'hfff;
rom[106967] = 12'hfff;
rom[106968] = 12'heee;
rom[106969] = 12'heee;
rom[106970] = 12'heee;
rom[106971] = 12'heee;
rom[106972] = 12'heee;
rom[106973] = 12'heee;
rom[106974] = 12'heee;
rom[106975] = 12'heee;
rom[106976] = 12'hddd;
rom[106977] = 12'hddd;
rom[106978] = 12'hddd;
rom[106979] = 12'hddd;
rom[106980] = 12'hddd;
rom[106981] = 12'hddd;
rom[106982] = 12'hddd;
rom[106983] = 12'hddd;
rom[106984] = 12'hccc;
rom[106985] = 12'hccc;
rom[106986] = 12'hccc;
rom[106987] = 12'hccc;
rom[106988] = 12'hccc;
rom[106989] = 12'hccc;
rom[106990] = 12'hccc;
rom[106991] = 12'hccc;
rom[106992] = 12'hccc;
rom[106993] = 12'hccc;
rom[106994] = 12'hccc;
rom[106995] = 12'hccc;
rom[106996] = 12'hccc;
rom[106997] = 12'hccc;
rom[106998] = 12'hbbb;
rom[106999] = 12'hbbb;
rom[107000] = 12'hbbb;
rom[107001] = 12'hbbb;
rom[107002] = 12'hbbb;
rom[107003] = 12'hbbb;
rom[107004] = 12'hbbb;
rom[107005] = 12'hbbb;
rom[107006] = 12'hbbb;
rom[107007] = 12'hbbb;
rom[107008] = 12'hbbb;
rom[107009] = 12'hbbb;
rom[107010] = 12'hbbb;
rom[107011] = 12'hbbb;
rom[107012] = 12'hbbb;
rom[107013] = 12'hbbb;
rom[107014] = 12'hbbb;
rom[107015] = 12'hbbb;
rom[107016] = 12'hbbb;
rom[107017] = 12'hccc;
rom[107018] = 12'hccc;
rom[107019] = 12'hddd;
rom[107020] = 12'hddd;
rom[107021] = 12'hddd;
rom[107022] = 12'heee;
rom[107023] = 12'heee;
rom[107024] = 12'heee;
rom[107025] = 12'heee;
rom[107026] = 12'hfff;
rom[107027] = 12'hfff;
rom[107028] = 12'hfff;
rom[107029] = 12'hfff;
rom[107030] = 12'hfff;
rom[107031] = 12'hfff;
rom[107032] = 12'hfff;
rom[107033] = 12'hfff;
rom[107034] = 12'hfff;
rom[107035] = 12'hfff;
rom[107036] = 12'hfff;
rom[107037] = 12'hfff;
rom[107038] = 12'hfff;
rom[107039] = 12'hfff;
rom[107040] = 12'hfff;
rom[107041] = 12'hfff;
rom[107042] = 12'hfff;
rom[107043] = 12'hfff;
rom[107044] = 12'hfff;
rom[107045] = 12'hfff;
rom[107046] = 12'hfff;
rom[107047] = 12'hfff;
rom[107048] = 12'hfff;
rom[107049] = 12'hfff;
rom[107050] = 12'hfff;
rom[107051] = 12'hfff;
rom[107052] = 12'hfff;
rom[107053] = 12'heee;
rom[107054] = 12'hddd;
rom[107055] = 12'hccc;
rom[107056] = 12'hbbb;
rom[107057] = 12'hbbb;
rom[107058] = 12'hbbb;
rom[107059] = 12'hbbb;
rom[107060] = 12'hccc;
rom[107061] = 12'hccc;
rom[107062] = 12'hddd;
rom[107063] = 12'heee;
rom[107064] = 12'heee;
rom[107065] = 12'hddd;
rom[107066] = 12'haaa;
rom[107067] = 12'h888;
rom[107068] = 12'h888;
rom[107069] = 12'haaa;
rom[107070] = 12'hccc;
rom[107071] = 12'hfff;
rom[107072] = 12'hbbb;
rom[107073] = 12'h888;
rom[107074] = 12'h444;
rom[107075] = 12'h333;
rom[107076] = 12'h333;
rom[107077] = 12'h222;
rom[107078] = 12'h222;
rom[107079] = 12'h333;
rom[107080] = 12'h666;
rom[107081] = 12'h999;
rom[107082] = 12'hddd;
rom[107083] = 12'heee;
rom[107084] = 12'hccc;
rom[107085] = 12'h888;
rom[107086] = 12'h666;
rom[107087] = 12'h555;
rom[107088] = 12'h444;
rom[107089] = 12'h555;
rom[107090] = 12'h555;
rom[107091] = 12'h444;
rom[107092] = 12'h333;
rom[107093] = 12'h333;
rom[107094] = 12'h444;
rom[107095] = 12'h666;
rom[107096] = 12'h999;
rom[107097] = 12'hccc;
rom[107098] = 12'hddd;
rom[107099] = 12'hbbb;
rom[107100] = 12'hbbb;
rom[107101] = 12'heee;
rom[107102] = 12'heee;
rom[107103] = 12'hccc;
rom[107104] = 12'h888;
rom[107105] = 12'h555;
rom[107106] = 12'h333;
rom[107107] = 12'h333;
rom[107108] = 12'h333;
rom[107109] = 12'h222;
rom[107110] = 12'h222;
rom[107111] = 12'h222;
rom[107112] = 12'h222;
rom[107113] = 12'h111;
rom[107114] = 12'h111;
rom[107115] = 12'h111;
rom[107116] = 12'h111;
rom[107117] = 12'h111;
rom[107118] = 12'h111;
rom[107119] = 12'h111;
rom[107120] = 12'h  0;
rom[107121] = 12'h111;
rom[107122] = 12'h111;
rom[107123] = 12'h111;
rom[107124] = 12'h111;
rom[107125] = 12'h222;
rom[107126] = 12'h444;
rom[107127] = 12'h555;
rom[107128] = 12'h555;
rom[107129] = 12'h444;
rom[107130] = 12'h333;
rom[107131] = 12'h222;
rom[107132] = 12'h111;
rom[107133] = 12'h111;
rom[107134] = 12'h111;
rom[107135] = 12'h111;
rom[107136] = 12'h111;
rom[107137] = 12'h111;
rom[107138] = 12'h  0;
rom[107139] = 12'h111;
rom[107140] = 12'h111;
rom[107141] = 12'h111;
rom[107142] = 12'h  0;
rom[107143] = 12'h  0;
rom[107144] = 12'h111;
rom[107145] = 12'h111;
rom[107146] = 12'h111;
rom[107147] = 12'h111;
rom[107148] = 12'h111;
rom[107149] = 12'h111;
rom[107150] = 12'h222;
rom[107151] = 12'h333;
rom[107152] = 12'h555;
rom[107153] = 12'h888;
rom[107154] = 12'hccc;
rom[107155] = 12'heee;
rom[107156] = 12'heee;
rom[107157] = 12'hbbb;
rom[107158] = 12'h777;
rom[107159] = 12'h444;
rom[107160] = 12'h333;
rom[107161] = 12'h333;
rom[107162] = 12'h222;
rom[107163] = 12'h222;
rom[107164] = 12'h222;
rom[107165] = 12'h111;
rom[107166] = 12'h111;
rom[107167] = 12'h111;
rom[107168] = 12'h111;
rom[107169] = 12'h111;
rom[107170] = 12'h  0;
rom[107171] = 12'h  0;
rom[107172] = 12'h  0;
rom[107173] = 12'h  0;
rom[107174] = 12'h  0;
rom[107175] = 12'h  0;
rom[107176] = 12'h  0;
rom[107177] = 12'h  0;
rom[107178] = 12'h  0;
rom[107179] = 12'h  0;
rom[107180] = 12'h  0;
rom[107181] = 12'h  0;
rom[107182] = 12'h  0;
rom[107183] = 12'h  0;
rom[107184] = 12'h  0;
rom[107185] = 12'h  0;
rom[107186] = 12'h  0;
rom[107187] = 12'h  0;
rom[107188] = 12'h  0;
rom[107189] = 12'h  0;
rom[107190] = 12'h  0;
rom[107191] = 12'h  0;
rom[107192] = 12'h  0;
rom[107193] = 12'h  0;
rom[107194] = 12'h  0;
rom[107195] = 12'h  0;
rom[107196] = 12'h  0;
rom[107197] = 12'h  0;
rom[107198] = 12'h111;
rom[107199] = 12'h111;
rom[107200] = 12'hfff;
rom[107201] = 12'hfff;
rom[107202] = 12'hfff;
rom[107203] = 12'hfff;
rom[107204] = 12'hfff;
rom[107205] = 12'hfff;
rom[107206] = 12'hfff;
rom[107207] = 12'hfff;
rom[107208] = 12'hfff;
rom[107209] = 12'hfff;
rom[107210] = 12'hfff;
rom[107211] = 12'hfff;
rom[107212] = 12'hfff;
rom[107213] = 12'hfff;
rom[107214] = 12'hfff;
rom[107215] = 12'hfff;
rom[107216] = 12'hfff;
rom[107217] = 12'hfff;
rom[107218] = 12'hfff;
rom[107219] = 12'hfff;
rom[107220] = 12'hfff;
rom[107221] = 12'hfff;
rom[107222] = 12'hfff;
rom[107223] = 12'hfff;
rom[107224] = 12'hfff;
rom[107225] = 12'hfff;
rom[107226] = 12'hfff;
rom[107227] = 12'hfff;
rom[107228] = 12'hfff;
rom[107229] = 12'hfff;
rom[107230] = 12'hfff;
rom[107231] = 12'hfff;
rom[107232] = 12'hfff;
rom[107233] = 12'hfff;
rom[107234] = 12'hfff;
rom[107235] = 12'hfff;
rom[107236] = 12'hfff;
rom[107237] = 12'hfff;
rom[107238] = 12'hfff;
rom[107239] = 12'hfff;
rom[107240] = 12'hfff;
rom[107241] = 12'hfff;
rom[107242] = 12'hfff;
rom[107243] = 12'hfff;
rom[107244] = 12'hfff;
rom[107245] = 12'hfff;
rom[107246] = 12'hfff;
rom[107247] = 12'hfff;
rom[107248] = 12'hfff;
rom[107249] = 12'hfff;
rom[107250] = 12'hfff;
rom[107251] = 12'hfff;
rom[107252] = 12'hfff;
rom[107253] = 12'hfff;
rom[107254] = 12'heee;
rom[107255] = 12'heee;
rom[107256] = 12'heee;
rom[107257] = 12'heee;
rom[107258] = 12'heee;
rom[107259] = 12'heee;
rom[107260] = 12'heee;
rom[107261] = 12'heee;
rom[107262] = 12'heee;
rom[107263] = 12'heee;
rom[107264] = 12'heee;
rom[107265] = 12'heee;
rom[107266] = 12'heee;
rom[107267] = 12'heee;
rom[107268] = 12'heee;
rom[107269] = 12'heee;
rom[107270] = 12'heee;
rom[107271] = 12'heee;
rom[107272] = 12'heee;
rom[107273] = 12'heee;
rom[107274] = 12'heee;
rom[107275] = 12'heee;
rom[107276] = 12'heee;
rom[107277] = 12'heee;
rom[107278] = 12'heee;
rom[107279] = 12'heee;
rom[107280] = 12'hddd;
rom[107281] = 12'hddd;
rom[107282] = 12'hddd;
rom[107283] = 12'hccc;
rom[107284] = 12'hccc;
rom[107285] = 12'hccc;
rom[107286] = 12'hccc;
rom[107287] = 12'hccc;
rom[107288] = 12'hccc;
rom[107289] = 12'hccc;
rom[107290] = 12'hccc;
rom[107291] = 12'hddd;
rom[107292] = 12'heee;
rom[107293] = 12'hfff;
rom[107294] = 12'heee;
rom[107295] = 12'hddd;
rom[107296] = 12'hccc;
rom[107297] = 12'hccc;
rom[107298] = 12'hddd;
rom[107299] = 12'hddd;
rom[107300] = 12'heee;
rom[107301] = 12'heee;
rom[107302] = 12'hddd;
rom[107303] = 12'hccc;
rom[107304] = 12'hbbb;
rom[107305] = 12'hbbb;
rom[107306] = 12'hbbb;
rom[107307] = 12'hbbb;
rom[107308] = 12'hbbb;
rom[107309] = 12'hbbb;
rom[107310] = 12'hccc;
rom[107311] = 12'hddd;
rom[107312] = 12'hfff;
rom[107313] = 12'hfff;
rom[107314] = 12'heee;
rom[107315] = 12'hccc;
rom[107316] = 12'hbbb;
rom[107317] = 12'hbbb;
rom[107318] = 12'hbbb;
rom[107319] = 12'haaa;
rom[107320] = 12'haaa;
rom[107321] = 12'haaa;
rom[107322] = 12'h999;
rom[107323] = 12'haaa;
rom[107324] = 12'haaa;
rom[107325] = 12'haaa;
rom[107326] = 12'haaa;
rom[107327] = 12'haaa;
rom[107328] = 12'haaa;
rom[107329] = 12'hbbb;
rom[107330] = 12'hddd;
rom[107331] = 12'heee;
rom[107332] = 12'hddd;
rom[107333] = 12'hccc;
rom[107334] = 12'hccc;
rom[107335] = 12'hccc;
rom[107336] = 12'hccc;
rom[107337] = 12'hccc;
rom[107338] = 12'hccc;
rom[107339] = 12'hccc;
rom[107340] = 12'hccc;
rom[107341] = 12'hccc;
rom[107342] = 12'hccc;
rom[107343] = 12'hddd;
rom[107344] = 12'hddd;
rom[107345] = 12'hddd;
rom[107346] = 12'heee;
rom[107347] = 12'hfff;
rom[107348] = 12'hfff;
rom[107349] = 12'hfff;
rom[107350] = 12'hfff;
rom[107351] = 12'hfff;
rom[107352] = 12'hfff;
rom[107353] = 12'hfff;
rom[107354] = 12'hfff;
rom[107355] = 12'hfff;
rom[107356] = 12'hfff;
rom[107357] = 12'hfff;
rom[107358] = 12'hfff;
rom[107359] = 12'hfff;
rom[107360] = 12'hfff;
rom[107361] = 12'hfff;
rom[107362] = 12'hfff;
rom[107363] = 12'hfff;
rom[107364] = 12'hfff;
rom[107365] = 12'hfff;
rom[107366] = 12'hfff;
rom[107367] = 12'hfff;
rom[107368] = 12'heee;
rom[107369] = 12'heee;
rom[107370] = 12'heee;
rom[107371] = 12'heee;
rom[107372] = 12'heee;
rom[107373] = 12'heee;
rom[107374] = 12'heee;
rom[107375] = 12'heee;
rom[107376] = 12'heee;
rom[107377] = 12'heee;
rom[107378] = 12'hddd;
rom[107379] = 12'hddd;
rom[107380] = 12'hddd;
rom[107381] = 12'hddd;
rom[107382] = 12'hddd;
rom[107383] = 12'hddd;
rom[107384] = 12'hccc;
rom[107385] = 12'hccc;
rom[107386] = 12'hccc;
rom[107387] = 12'hccc;
rom[107388] = 12'hccc;
rom[107389] = 12'hccc;
rom[107390] = 12'hccc;
rom[107391] = 12'hccc;
rom[107392] = 12'hccc;
rom[107393] = 12'hccc;
rom[107394] = 12'hccc;
rom[107395] = 12'hccc;
rom[107396] = 12'hccc;
rom[107397] = 12'hccc;
rom[107398] = 12'hbbb;
rom[107399] = 12'hbbb;
rom[107400] = 12'hbbb;
rom[107401] = 12'hbbb;
rom[107402] = 12'hbbb;
rom[107403] = 12'hbbb;
rom[107404] = 12'hbbb;
rom[107405] = 12'hbbb;
rom[107406] = 12'hbbb;
rom[107407] = 12'hbbb;
rom[107408] = 12'hbbb;
rom[107409] = 12'hbbb;
rom[107410] = 12'hbbb;
rom[107411] = 12'hbbb;
rom[107412] = 12'hbbb;
rom[107413] = 12'hbbb;
rom[107414] = 12'hbbb;
rom[107415] = 12'hccc;
rom[107416] = 12'hccc;
rom[107417] = 12'hccc;
rom[107418] = 12'hccc;
rom[107419] = 12'hddd;
rom[107420] = 12'hddd;
rom[107421] = 12'hddd;
rom[107422] = 12'heee;
rom[107423] = 12'heee;
rom[107424] = 12'heee;
rom[107425] = 12'hfff;
rom[107426] = 12'hfff;
rom[107427] = 12'hfff;
rom[107428] = 12'hfff;
rom[107429] = 12'hfff;
rom[107430] = 12'hfff;
rom[107431] = 12'hfff;
rom[107432] = 12'hfff;
rom[107433] = 12'hfff;
rom[107434] = 12'hfff;
rom[107435] = 12'hfff;
rom[107436] = 12'hfff;
rom[107437] = 12'hfff;
rom[107438] = 12'hfff;
rom[107439] = 12'hfff;
rom[107440] = 12'hfff;
rom[107441] = 12'hfff;
rom[107442] = 12'hfff;
rom[107443] = 12'hfff;
rom[107444] = 12'hfff;
rom[107445] = 12'hfff;
rom[107446] = 12'hfff;
rom[107447] = 12'hfff;
rom[107448] = 12'heee;
rom[107449] = 12'hfff;
rom[107450] = 12'hfff;
rom[107451] = 12'hfff;
rom[107452] = 12'heee;
rom[107453] = 12'hccc;
rom[107454] = 12'hbbb;
rom[107455] = 12'haaa;
rom[107456] = 12'haaa;
rom[107457] = 12'haaa;
rom[107458] = 12'haaa;
rom[107459] = 12'haaa;
rom[107460] = 12'hbbb;
rom[107461] = 12'hccc;
rom[107462] = 12'heee;
rom[107463] = 12'heee;
rom[107464] = 12'hfff;
rom[107465] = 12'hddd;
rom[107466] = 12'haaa;
rom[107467] = 12'h888;
rom[107468] = 12'h888;
rom[107469] = 12'h999;
rom[107470] = 12'hbbb;
rom[107471] = 12'hfff;
rom[107472] = 12'hccc;
rom[107473] = 12'h888;
rom[107474] = 12'h444;
rom[107475] = 12'h333;
rom[107476] = 12'h333;
rom[107477] = 12'h222;
rom[107478] = 12'h222;
rom[107479] = 12'h222;
rom[107480] = 12'h333;
rom[107481] = 12'h666;
rom[107482] = 12'hbbb;
rom[107483] = 12'heee;
rom[107484] = 12'hddd;
rom[107485] = 12'haaa;
rom[107486] = 12'h777;
rom[107487] = 12'h555;
rom[107488] = 12'h555;
rom[107489] = 12'h444;
rom[107490] = 12'h444;
rom[107491] = 12'h333;
rom[107492] = 12'h333;
rom[107493] = 12'h333;
rom[107494] = 12'h333;
rom[107495] = 12'h444;
rom[107496] = 12'h555;
rom[107497] = 12'haaa;
rom[107498] = 12'hddd;
rom[107499] = 12'hccc;
rom[107500] = 12'hbbb;
rom[107501] = 12'hccc;
rom[107502] = 12'hddd;
rom[107503] = 12'heee;
rom[107504] = 12'hbbb;
rom[107505] = 12'h888;
rom[107506] = 12'h444;
rom[107507] = 12'h222;
rom[107508] = 12'h333;
rom[107509] = 12'h333;
rom[107510] = 12'h222;
rom[107511] = 12'h222;
rom[107512] = 12'h222;
rom[107513] = 12'h111;
rom[107514] = 12'h111;
rom[107515] = 12'h111;
rom[107516] = 12'h111;
rom[107517] = 12'h111;
rom[107518] = 12'h111;
rom[107519] = 12'h111;
rom[107520] = 12'h  0;
rom[107521] = 12'h111;
rom[107522] = 12'h111;
rom[107523] = 12'h111;
rom[107524] = 12'h111;
rom[107525] = 12'h111;
rom[107526] = 12'h333;
rom[107527] = 12'h444;
rom[107528] = 12'h444;
rom[107529] = 12'h444;
rom[107530] = 12'h333;
rom[107531] = 12'h222;
rom[107532] = 12'h222;
rom[107533] = 12'h111;
rom[107534] = 12'h111;
rom[107535] = 12'h111;
rom[107536] = 12'h111;
rom[107537] = 12'h111;
rom[107538] = 12'h111;
rom[107539] = 12'h  0;
rom[107540] = 12'h  0;
rom[107541] = 12'h  0;
rom[107542] = 12'h  0;
rom[107543] = 12'h  0;
rom[107544] = 12'h  0;
rom[107545] = 12'h  0;
rom[107546] = 12'h  0;
rom[107547] = 12'h111;
rom[107548] = 12'h111;
rom[107549] = 12'h111;
rom[107550] = 12'h111;
rom[107551] = 12'h222;
rom[107552] = 12'h222;
rom[107553] = 12'h555;
rom[107554] = 12'h888;
rom[107555] = 12'hbbb;
rom[107556] = 12'heee;
rom[107557] = 12'heee;
rom[107558] = 12'hbbb;
rom[107559] = 12'h777;
rom[107560] = 12'h444;
rom[107561] = 12'h333;
rom[107562] = 12'h222;
rom[107563] = 12'h222;
rom[107564] = 12'h222;
rom[107565] = 12'h111;
rom[107566] = 12'h111;
rom[107567] = 12'h111;
rom[107568] = 12'h111;
rom[107569] = 12'h111;
rom[107570] = 12'h  0;
rom[107571] = 12'h  0;
rom[107572] = 12'h  0;
rom[107573] = 12'h  0;
rom[107574] = 12'h  0;
rom[107575] = 12'h  0;
rom[107576] = 12'h  0;
rom[107577] = 12'h  0;
rom[107578] = 12'h  0;
rom[107579] = 12'h  0;
rom[107580] = 12'h  0;
rom[107581] = 12'h  0;
rom[107582] = 12'h  0;
rom[107583] = 12'h  0;
rom[107584] = 12'h  0;
rom[107585] = 12'h  0;
rom[107586] = 12'h  0;
rom[107587] = 12'h  0;
rom[107588] = 12'h  0;
rom[107589] = 12'h  0;
rom[107590] = 12'h  0;
rom[107591] = 12'h  0;
rom[107592] = 12'h  0;
rom[107593] = 12'h  0;
rom[107594] = 12'h  0;
rom[107595] = 12'h  0;
rom[107596] = 12'h  0;
rom[107597] = 12'h  0;
rom[107598] = 12'h  0;
rom[107599] = 12'h  0;
rom[107600] = 12'hfff;
rom[107601] = 12'hfff;
rom[107602] = 12'hfff;
rom[107603] = 12'hfff;
rom[107604] = 12'hfff;
rom[107605] = 12'hfff;
rom[107606] = 12'hfff;
rom[107607] = 12'hfff;
rom[107608] = 12'hfff;
rom[107609] = 12'hfff;
rom[107610] = 12'hfff;
rom[107611] = 12'hfff;
rom[107612] = 12'hfff;
rom[107613] = 12'hfff;
rom[107614] = 12'hfff;
rom[107615] = 12'hfff;
rom[107616] = 12'hfff;
rom[107617] = 12'hfff;
rom[107618] = 12'hfff;
rom[107619] = 12'hfff;
rom[107620] = 12'hfff;
rom[107621] = 12'hfff;
rom[107622] = 12'hfff;
rom[107623] = 12'hfff;
rom[107624] = 12'hfff;
rom[107625] = 12'hfff;
rom[107626] = 12'hfff;
rom[107627] = 12'hfff;
rom[107628] = 12'hfff;
rom[107629] = 12'hfff;
rom[107630] = 12'hfff;
rom[107631] = 12'hfff;
rom[107632] = 12'hfff;
rom[107633] = 12'hfff;
rom[107634] = 12'hfff;
rom[107635] = 12'hfff;
rom[107636] = 12'hfff;
rom[107637] = 12'hfff;
rom[107638] = 12'hfff;
rom[107639] = 12'hfff;
rom[107640] = 12'hfff;
rom[107641] = 12'hfff;
rom[107642] = 12'hfff;
rom[107643] = 12'hfff;
rom[107644] = 12'hfff;
rom[107645] = 12'hfff;
rom[107646] = 12'hfff;
rom[107647] = 12'hfff;
rom[107648] = 12'hfff;
rom[107649] = 12'hfff;
rom[107650] = 12'hfff;
rom[107651] = 12'hfff;
rom[107652] = 12'hfff;
rom[107653] = 12'hfff;
rom[107654] = 12'heee;
rom[107655] = 12'heee;
rom[107656] = 12'heee;
rom[107657] = 12'heee;
rom[107658] = 12'heee;
rom[107659] = 12'heee;
rom[107660] = 12'heee;
rom[107661] = 12'heee;
rom[107662] = 12'heee;
rom[107663] = 12'heee;
rom[107664] = 12'heee;
rom[107665] = 12'heee;
rom[107666] = 12'heee;
rom[107667] = 12'heee;
rom[107668] = 12'heee;
rom[107669] = 12'heee;
rom[107670] = 12'heee;
rom[107671] = 12'hddd;
rom[107672] = 12'hddd;
rom[107673] = 12'heee;
rom[107674] = 12'heee;
rom[107675] = 12'heee;
rom[107676] = 12'heee;
rom[107677] = 12'heee;
rom[107678] = 12'heee;
rom[107679] = 12'heee;
rom[107680] = 12'hddd;
rom[107681] = 12'hccc;
rom[107682] = 12'hccc;
rom[107683] = 12'hccc;
rom[107684] = 12'hccc;
rom[107685] = 12'hccc;
rom[107686] = 12'hccc;
rom[107687] = 12'hccc;
rom[107688] = 12'hccc;
rom[107689] = 12'hccc;
rom[107690] = 12'hccc;
rom[107691] = 12'hddd;
rom[107692] = 12'heee;
rom[107693] = 12'hfff;
rom[107694] = 12'heee;
rom[107695] = 12'hbbb;
rom[107696] = 12'hccc;
rom[107697] = 12'hccc;
rom[107698] = 12'hddd;
rom[107699] = 12'heee;
rom[107700] = 12'heee;
rom[107701] = 12'hddd;
rom[107702] = 12'hccc;
rom[107703] = 12'hbbb;
rom[107704] = 12'hbbb;
rom[107705] = 12'hbbb;
rom[107706] = 12'hbbb;
rom[107707] = 12'hbbb;
rom[107708] = 12'haaa;
rom[107709] = 12'hbbb;
rom[107710] = 12'hddd;
rom[107711] = 12'heee;
rom[107712] = 12'hfff;
rom[107713] = 12'heee;
rom[107714] = 12'hccc;
rom[107715] = 12'hbbb;
rom[107716] = 12'hbbb;
rom[107717] = 12'hbbb;
rom[107718] = 12'haaa;
rom[107719] = 12'haaa;
rom[107720] = 12'haaa;
rom[107721] = 12'h999;
rom[107722] = 12'h999;
rom[107723] = 12'h999;
rom[107724] = 12'h999;
rom[107725] = 12'h999;
rom[107726] = 12'h999;
rom[107727] = 12'haaa;
rom[107728] = 12'haaa;
rom[107729] = 12'hbbb;
rom[107730] = 12'hddd;
rom[107731] = 12'hddd;
rom[107732] = 12'hccc;
rom[107733] = 12'hbbb;
rom[107734] = 12'hbbb;
rom[107735] = 12'hccc;
rom[107736] = 12'hbbb;
rom[107737] = 12'hccc;
rom[107738] = 12'hccc;
rom[107739] = 12'hccc;
rom[107740] = 12'hccc;
rom[107741] = 12'hccc;
rom[107742] = 12'hccc;
rom[107743] = 12'hccc;
rom[107744] = 12'hccc;
rom[107745] = 12'hddd;
rom[107746] = 12'hddd;
rom[107747] = 12'heee;
rom[107748] = 12'heee;
rom[107749] = 12'hfff;
rom[107750] = 12'hfff;
rom[107751] = 12'hfff;
rom[107752] = 12'hfff;
rom[107753] = 12'hfff;
rom[107754] = 12'hfff;
rom[107755] = 12'hfff;
rom[107756] = 12'hfff;
rom[107757] = 12'hfff;
rom[107758] = 12'hfff;
rom[107759] = 12'hfff;
rom[107760] = 12'hfff;
rom[107761] = 12'hfff;
rom[107762] = 12'hfff;
rom[107763] = 12'hfff;
rom[107764] = 12'hfff;
rom[107765] = 12'hfff;
rom[107766] = 12'hfff;
rom[107767] = 12'hfff;
rom[107768] = 12'hfff;
rom[107769] = 12'hfff;
rom[107770] = 12'heee;
rom[107771] = 12'heee;
rom[107772] = 12'heee;
rom[107773] = 12'heee;
rom[107774] = 12'heee;
rom[107775] = 12'heee;
rom[107776] = 12'heee;
rom[107777] = 12'heee;
rom[107778] = 12'heee;
rom[107779] = 12'hddd;
rom[107780] = 12'hddd;
rom[107781] = 12'hddd;
rom[107782] = 12'hddd;
rom[107783] = 12'hddd;
rom[107784] = 12'hccc;
rom[107785] = 12'hccc;
rom[107786] = 12'hccc;
rom[107787] = 12'hccc;
rom[107788] = 12'hccc;
rom[107789] = 12'hccc;
rom[107790] = 12'hccc;
rom[107791] = 12'hccc;
rom[107792] = 12'hccc;
rom[107793] = 12'hccc;
rom[107794] = 12'hccc;
rom[107795] = 12'hccc;
rom[107796] = 12'hccc;
rom[107797] = 12'hccc;
rom[107798] = 12'hccc;
rom[107799] = 12'hbbb;
rom[107800] = 12'hbbb;
rom[107801] = 12'hbbb;
rom[107802] = 12'hbbb;
rom[107803] = 12'hbbb;
rom[107804] = 12'hbbb;
rom[107805] = 12'hbbb;
rom[107806] = 12'hbbb;
rom[107807] = 12'hbbb;
rom[107808] = 12'hbbb;
rom[107809] = 12'hbbb;
rom[107810] = 12'hbbb;
rom[107811] = 12'hbbb;
rom[107812] = 12'hbbb;
rom[107813] = 12'hbbb;
rom[107814] = 12'hbbb;
rom[107815] = 12'hccc;
rom[107816] = 12'hccc;
rom[107817] = 12'hccc;
rom[107818] = 12'hddd;
rom[107819] = 12'hddd;
rom[107820] = 12'heee;
rom[107821] = 12'heee;
rom[107822] = 12'heee;
rom[107823] = 12'hfff;
rom[107824] = 12'hfff;
rom[107825] = 12'hfff;
rom[107826] = 12'hfff;
rom[107827] = 12'hfff;
rom[107828] = 12'hfff;
rom[107829] = 12'hfff;
rom[107830] = 12'hfff;
rom[107831] = 12'hfff;
rom[107832] = 12'hfff;
rom[107833] = 12'hfff;
rom[107834] = 12'hfff;
rom[107835] = 12'hfff;
rom[107836] = 12'hfff;
rom[107837] = 12'hfff;
rom[107838] = 12'hfff;
rom[107839] = 12'hfff;
rom[107840] = 12'hfff;
rom[107841] = 12'hfff;
rom[107842] = 12'hfff;
rom[107843] = 12'hfff;
rom[107844] = 12'hfff;
rom[107845] = 12'hfff;
rom[107846] = 12'heee;
rom[107847] = 12'heee;
rom[107848] = 12'heee;
rom[107849] = 12'heee;
rom[107850] = 12'hfff;
rom[107851] = 12'heee;
rom[107852] = 12'hddd;
rom[107853] = 12'hbbb;
rom[107854] = 12'haaa;
rom[107855] = 12'h999;
rom[107856] = 12'h999;
rom[107857] = 12'h999;
rom[107858] = 12'haaa;
rom[107859] = 12'haaa;
rom[107860] = 12'haaa;
rom[107861] = 12'hccc;
rom[107862] = 12'hddd;
rom[107863] = 12'heee;
rom[107864] = 12'hfff;
rom[107865] = 12'hddd;
rom[107866] = 12'haaa;
rom[107867] = 12'h888;
rom[107868] = 12'h888;
rom[107869] = 12'h777;
rom[107870] = 12'haaa;
rom[107871] = 12'heee;
rom[107872] = 12'hddd;
rom[107873] = 12'h999;
rom[107874] = 12'h444;
rom[107875] = 12'h333;
rom[107876] = 12'h222;
rom[107877] = 12'h222;
rom[107878] = 12'h222;
rom[107879] = 12'h222;
rom[107880] = 12'h222;
rom[107881] = 12'h444;
rom[107882] = 12'h888;
rom[107883] = 12'hccc;
rom[107884] = 12'heee;
rom[107885] = 12'hddd;
rom[107886] = 12'h999;
rom[107887] = 12'h555;
rom[107888] = 12'h555;
rom[107889] = 12'h444;
rom[107890] = 12'h444;
rom[107891] = 12'h333;
rom[107892] = 12'h333;
rom[107893] = 12'h333;
rom[107894] = 12'h333;
rom[107895] = 12'h222;
rom[107896] = 12'h333;
rom[107897] = 12'h666;
rom[107898] = 12'haaa;
rom[107899] = 12'hddd;
rom[107900] = 12'hccc;
rom[107901] = 12'hbbb;
rom[107902] = 12'hccc;
rom[107903] = 12'heee;
rom[107904] = 12'heee;
rom[107905] = 12'hbbb;
rom[107906] = 12'h666;
rom[107907] = 12'h333;
rom[107908] = 12'h333;
rom[107909] = 12'h333;
rom[107910] = 12'h222;
rom[107911] = 12'h222;
rom[107912] = 12'h222;
rom[107913] = 12'h111;
rom[107914] = 12'h111;
rom[107915] = 12'h111;
rom[107916] = 12'h111;
rom[107917] = 12'h111;
rom[107918] = 12'h111;
rom[107919] = 12'h  0;
rom[107920] = 12'h  0;
rom[107921] = 12'h111;
rom[107922] = 12'h111;
rom[107923] = 12'h111;
rom[107924] = 12'h  0;
rom[107925] = 12'h111;
rom[107926] = 12'h111;
rom[107927] = 12'h222;
rom[107928] = 12'h444;
rom[107929] = 12'h444;
rom[107930] = 12'h444;
rom[107931] = 12'h333;
rom[107932] = 12'h222;
rom[107933] = 12'h111;
rom[107934] = 12'h111;
rom[107935] = 12'h  0;
rom[107936] = 12'h111;
rom[107937] = 12'h111;
rom[107938] = 12'h  0;
rom[107939] = 12'h  0;
rom[107940] = 12'h  0;
rom[107941] = 12'h  0;
rom[107942] = 12'h  0;
rom[107943] = 12'h  0;
rom[107944] = 12'h  0;
rom[107945] = 12'h  0;
rom[107946] = 12'h  0;
rom[107947] = 12'h  0;
rom[107948] = 12'h  0;
rom[107949] = 12'h111;
rom[107950] = 12'h111;
rom[107951] = 12'h111;
rom[107952] = 12'h222;
rom[107953] = 12'h333;
rom[107954] = 12'h555;
rom[107955] = 12'h888;
rom[107956] = 12'hccc;
rom[107957] = 12'hfff;
rom[107958] = 12'hddd;
rom[107959] = 12'hbbb;
rom[107960] = 12'h666;
rom[107961] = 12'h444;
rom[107962] = 12'h333;
rom[107963] = 12'h222;
rom[107964] = 12'h222;
rom[107965] = 12'h222;
rom[107966] = 12'h111;
rom[107967] = 12'h111;
rom[107968] = 12'h111;
rom[107969] = 12'h111;
rom[107970] = 12'h111;
rom[107971] = 12'h  0;
rom[107972] = 12'h  0;
rom[107973] = 12'h  0;
rom[107974] = 12'h  0;
rom[107975] = 12'h  0;
rom[107976] = 12'h  0;
rom[107977] = 12'h  0;
rom[107978] = 12'h  0;
rom[107979] = 12'h  0;
rom[107980] = 12'h  0;
rom[107981] = 12'h  0;
rom[107982] = 12'h  0;
rom[107983] = 12'h  0;
rom[107984] = 12'h  0;
rom[107985] = 12'h  0;
rom[107986] = 12'h  0;
rom[107987] = 12'h  0;
rom[107988] = 12'h  0;
rom[107989] = 12'h  0;
rom[107990] = 12'h  0;
rom[107991] = 12'h  0;
rom[107992] = 12'h  0;
rom[107993] = 12'h  0;
rom[107994] = 12'h  0;
rom[107995] = 12'h  0;
rom[107996] = 12'h  0;
rom[107997] = 12'h  0;
rom[107998] = 12'h  0;
rom[107999] = 12'h  0;
rom[108000] = 12'hfff;
rom[108001] = 12'hfff;
rom[108002] = 12'hfff;
rom[108003] = 12'hfff;
rom[108004] = 12'hfff;
rom[108005] = 12'hfff;
rom[108006] = 12'hfff;
rom[108007] = 12'hfff;
rom[108008] = 12'hfff;
rom[108009] = 12'hfff;
rom[108010] = 12'hfff;
rom[108011] = 12'hfff;
rom[108012] = 12'hfff;
rom[108013] = 12'hfff;
rom[108014] = 12'hfff;
rom[108015] = 12'hfff;
rom[108016] = 12'hfff;
rom[108017] = 12'hfff;
rom[108018] = 12'hfff;
rom[108019] = 12'hfff;
rom[108020] = 12'hfff;
rom[108021] = 12'hfff;
rom[108022] = 12'hfff;
rom[108023] = 12'hfff;
rom[108024] = 12'hfff;
rom[108025] = 12'hfff;
rom[108026] = 12'hfff;
rom[108027] = 12'hfff;
rom[108028] = 12'hfff;
rom[108029] = 12'hfff;
rom[108030] = 12'hfff;
rom[108031] = 12'hfff;
rom[108032] = 12'hfff;
rom[108033] = 12'hfff;
rom[108034] = 12'hfff;
rom[108035] = 12'hfff;
rom[108036] = 12'hfff;
rom[108037] = 12'hfff;
rom[108038] = 12'hfff;
rom[108039] = 12'hfff;
rom[108040] = 12'hfff;
rom[108041] = 12'hfff;
rom[108042] = 12'hfff;
rom[108043] = 12'hfff;
rom[108044] = 12'hfff;
rom[108045] = 12'hfff;
rom[108046] = 12'hfff;
rom[108047] = 12'hfff;
rom[108048] = 12'hfff;
rom[108049] = 12'hfff;
rom[108050] = 12'hfff;
rom[108051] = 12'hfff;
rom[108052] = 12'hfff;
rom[108053] = 12'heee;
rom[108054] = 12'heee;
rom[108055] = 12'heee;
rom[108056] = 12'heee;
rom[108057] = 12'heee;
rom[108058] = 12'heee;
rom[108059] = 12'heee;
rom[108060] = 12'heee;
rom[108061] = 12'heee;
rom[108062] = 12'heee;
rom[108063] = 12'heee;
rom[108064] = 12'heee;
rom[108065] = 12'heee;
rom[108066] = 12'hddd;
rom[108067] = 12'heee;
rom[108068] = 12'heee;
rom[108069] = 12'heee;
rom[108070] = 12'hddd;
rom[108071] = 12'hddd;
rom[108072] = 12'hddd;
rom[108073] = 12'hddd;
rom[108074] = 12'heee;
rom[108075] = 12'heee;
rom[108076] = 12'heee;
rom[108077] = 12'heee;
rom[108078] = 12'hddd;
rom[108079] = 12'hddd;
rom[108080] = 12'hccc;
rom[108081] = 12'hccc;
rom[108082] = 12'hccc;
rom[108083] = 12'hccc;
rom[108084] = 12'hccc;
rom[108085] = 12'hccc;
rom[108086] = 12'hccc;
rom[108087] = 12'hccc;
rom[108088] = 12'hccc;
rom[108089] = 12'hccc;
rom[108090] = 12'hddd;
rom[108091] = 12'heee;
rom[108092] = 12'heee;
rom[108093] = 12'heee;
rom[108094] = 12'hddd;
rom[108095] = 12'hccc;
rom[108096] = 12'hddd;
rom[108097] = 12'hddd;
rom[108098] = 12'heee;
rom[108099] = 12'hddd;
rom[108100] = 12'hccc;
rom[108101] = 12'hbbb;
rom[108102] = 12'hbbb;
rom[108103] = 12'hbbb;
rom[108104] = 12'hbbb;
rom[108105] = 12'hbbb;
rom[108106] = 12'hbbb;
rom[108107] = 12'haaa;
rom[108108] = 12'haaa;
rom[108109] = 12'hbbb;
rom[108110] = 12'hddd;
rom[108111] = 12'hfff;
rom[108112] = 12'heee;
rom[108113] = 12'hccc;
rom[108114] = 12'hbbb;
rom[108115] = 12'haaa;
rom[108116] = 12'haaa;
rom[108117] = 12'haaa;
rom[108118] = 12'haaa;
rom[108119] = 12'haaa;
rom[108120] = 12'h999;
rom[108121] = 12'h999;
rom[108122] = 12'h999;
rom[108123] = 12'h999;
rom[108124] = 12'h999;
rom[108125] = 12'h999;
rom[108126] = 12'h999;
rom[108127] = 12'haaa;
rom[108128] = 12'hbbb;
rom[108129] = 12'hccc;
rom[108130] = 12'hddd;
rom[108131] = 12'hccc;
rom[108132] = 12'hbbb;
rom[108133] = 12'hbbb;
rom[108134] = 12'hbbb;
rom[108135] = 12'hbbb;
rom[108136] = 12'hbbb;
rom[108137] = 12'hbbb;
rom[108138] = 12'hbbb;
rom[108139] = 12'hbbb;
rom[108140] = 12'hbbb;
rom[108141] = 12'hbbb;
rom[108142] = 12'hccc;
rom[108143] = 12'hccc;
rom[108144] = 12'hccc;
rom[108145] = 12'hccc;
rom[108146] = 12'hddd;
rom[108147] = 12'hddd;
rom[108148] = 12'heee;
rom[108149] = 12'heee;
rom[108150] = 12'hfff;
rom[108151] = 12'hfff;
rom[108152] = 12'hfff;
rom[108153] = 12'hfff;
rom[108154] = 12'hfff;
rom[108155] = 12'hfff;
rom[108156] = 12'hfff;
rom[108157] = 12'hfff;
rom[108158] = 12'hfff;
rom[108159] = 12'hfff;
rom[108160] = 12'hfff;
rom[108161] = 12'hfff;
rom[108162] = 12'hfff;
rom[108163] = 12'hfff;
rom[108164] = 12'hfff;
rom[108165] = 12'hfff;
rom[108166] = 12'hfff;
rom[108167] = 12'hfff;
rom[108168] = 12'hfff;
rom[108169] = 12'hfff;
rom[108170] = 12'hfff;
rom[108171] = 12'heee;
rom[108172] = 12'heee;
rom[108173] = 12'heee;
rom[108174] = 12'heee;
rom[108175] = 12'heee;
rom[108176] = 12'heee;
rom[108177] = 12'heee;
rom[108178] = 12'heee;
rom[108179] = 12'hddd;
rom[108180] = 12'hddd;
rom[108181] = 12'hddd;
rom[108182] = 12'hddd;
rom[108183] = 12'hddd;
rom[108184] = 12'hccc;
rom[108185] = 12'hccc;
rom[108186] = 12'hccc;
rom[108187] = 12'hccc;
rom[108188] = 12'hccc;
rom[108189] = 12'hccc;
rom[108190] = 12'hccc;
rom[108191] = 12'hccc;
rom[108192] = 12'hccc;
rom[108193] = 12'hccc;
rom[108194] = 12'hccc;
rom[108195] = 12'hccc;
rom[108196] = 12'hccc;
rom[108197] = 12'hccc;
rom[108198] = 12'hccc;
rom[108199] = 12'hccc;
rom[108200] = 12'hbbb;
rom[108201] = 12'hbbb;
rom[108202] = 12'hbbb;
rom[108203] = 12'hbbb;
rom[108204] = 12'hbbb;
rom[108205] = 12'hbbb;
rom[108206] = 12'hbbb;
rom[108207] = 12'hbbb;
rom[108208] = 12'hbbb;
rom[108209] = 12'hbbb;
rom[108210] = 12'hbbb;
rom[108211] = 12'hbbb;
rom[108212] = 12'hbbb;
rom[108213] = 12'hbbb;
rom[108214] = 12'hccc;
rom[108215] = 12'hccc;
rom[108216] = 12'hddd;
rom[108217] = 12'hddd;
rom[108218] = 12'hddd;
rom[108219] = 12'heee;
rom[108220] = 12'heee;
rom[108221] = 12'heee;
rom[108222] = 12'hfff;
rom[108223] = 12'hfff;
rom[108224] = 12'hfff;
rom[108225] = 12'hfff;
rom[108226] = 12'hfff;
rom[108227] = 12'hfff;
rom[108228] = 12'hfff;
rom[108229] = 12'hfff;
rom[108230] = 12'hfff;
rom[108231] = 12'hfff;
rom[108232] = 12'hfff;
rom[108233] = 12'hfff;
rom[108234] = 12'hfff;
rom[108235] = 12'hfff;
rom[108236] = 12'hfff;
rom[108237] = 12'hfff;
rom[108238] = 12'hfff;
rom[108239] = 12'hfff;
rom[108240] = 12'hfff;
rom[108241] = 12'hfff;
rom[108242] = 12'heee;
rom[108243] = 12'heee;
rom[108244] = 12'hddd;
rom[108245] = 12'hddd;
rom[108246] = 12'hddd;
rom[108247] = 12'hddd;
rom[108248] = 12'heee;
rom[108249] = 12'heee;
rom[108250] = 12'heee;
rom[108251] = 12'hddd;
rom[108252] = 12'hbbb;
rom[108253] = 12'h999;
rom[108254] = 12'h888;
rom[108255] = 12'h888;
rom[108256] = 12'h777;
rom[108257] = 12'h888;
rom[108258] = 12'h999;
rom[108259] = 12'h999;
rom[108260] = 12'h999;
rom[108261] = 12'hbbb;
rom[108262] = 12'hddd;
rom[108263] = 12'hfff;
rom[108264] = 12'hfff;
rom[108265] = 12'hddd;
rom[108266] = 12'haaa;
rom[108267] = 12'h888;
rom[108268] = 12'h888;
rom[108269] = 12'h666;
rom[108270] = 12'h888;
rom[108271] = 12'hccc;
rom[108272] = 12'heee;
rom[108273] = 12'haaa;
rom[108274] = 12'h555;
rom[108275] = 12'h222;
rom[108276] = 12'h222;
rom[108277] = 12'h222;
rom[108278] = 12'h222;
rom[108279] = 12'h222;
rom[108280] = 12'h111;
rom[108281] = 12'h111;
rom[108282] = 12'h444;
rom[108283] = 12'haaa;
rom[108284] = 12'heee;
rom[108285] = 12'heee;
rom[108286] = 12'hbbb;
rom[108287] = 12'h777;
rom[108288] = 12'h555;
rom[108289] = 12'h444;
rom[108290] = 12'h444;
rom[108291] = 12'h333;
rom[108292] = 12'h333;
rom[108293] = 12'h333;
rom[108294] = 12'h222;
rom[108295] = 12'h222;
rom[108296] = 12'h333;
rom[108297] = 12'h333;
rom[108298] = 12'h666;
rom[108299] = 12'hbbb;
rom[108300] = 12'hccc;
rom[108301] = 12'hbbb;
rom[108302] = 12'hbbb;
rom[108303] = 12'hddd;
rom[108304] = 12'heee;
rom[108305] = 12'hddd;
rom[108306] = 12'haaa;
rom[108307] = 12'h666;
rom[108308] = 12'h333;
rom[108309] = 12'h333;
rom[108310] = 12'h333;
rom[108311] = 12'h222;
rom[108312] = 12'h222;
rom[108313] = 12'h111;
rom[108314] = 12'h111;
rom[108315] = 12'h111;
rom[108316] = 12'h111;
rom[108317] = 12'h111;
rom[108318] = 12'h111;
rom[108319] = 12'h  0;
rom[108320] = 12'h111;
rom[108321] = 12'h111;
rom[108322] = 12'h111;
rom[108323] = 12'h111;
rom[108324] = 12'h  0;
rom[108325] = 12'h111;
rom[108326] = 12'h111;
rom[108327] = 12'h222;
rom[108328] = 12'h333;
rom[108329] = 12'h333;
rom[108330] = 12'h333;
rom[108331] = 12'h333;
rom[108332] = 12'h222;
rom[108333] = 12'h111;
rom[108334] = 12'h  0;
rom[108335] = 12'h  0;
rom[108336] = 12'h  0;
rom[108337] = 12'h  0;
rom[108338] = 12'h  0;
rom[108339] = 12'h  0;
rom[108340] = 12'h  0;
rom[108341] = 12'h  0;
rom[108342] = 12'h  0;
rom[108343] = 12'h  0;
rom[108344] = 12'h  0;
rom[108345] = 12'h  0;
rom[108346] = 12'h  0;
rom[108347] = 12'h  0;
rom[108348] = 12'h  0;
rom[108349] = 12'h111;
rom[108350] = 12'h111;
rom[108351] = 12'h111;
rom[108352] = 12'h111;
rom[108353] = 12'h222;
rom[108354] = 12'h333;
rom[108355] = 12'h555;
rom[108356] = 12'h888;
rom[108357] = 12'hccc;
rom[108358] = 12'heee;
rom[108359] = 12'heee;
rom[108360] = 12'h999;
rom[108361] = 12'h777;
rom[108362] = 12'h444;
rom[108363] = 12'h333;
rom[108364] = 12'h333;
rom[108365] = 12'h222;
rom[108366] = 12'h222;
rom[108367] = 12'h111;
rom[108368] = 12'h111;
rom[108369] = 12'h111;
rom[108370] = 12'h111;
rom[108371] = 12'h  0;
rom[108372] = 12'h  0;
rom[108373] = 12'h  0;
rom[108374] = 12'h  0;
rom[108375] = 12'h  0;
rom[108376] = 12'h  0;
rom[108377] = 12'h  0;
rom[108378] = 12'h  0;
rom[108379] = 12'h  0;
rom[108380] = 12'h  0;
rom[108381] = 12'h  0;
rom[108382] = 12'h  0;
rom[108383] = 12'h  0;
rom[108384] = 12'h  0;
rom[108385] = 12'h  0;
rom[108386] = 12'h  0;
rom[108387] = 12'h  0;
rom[108388] = 12'h  0;
rom[108389] = 12'h  0;
rom[108390] = 12'h  0;
rom[108391] = 12'h  0;
rom[108392] = 12'h  0;
rom[108393] = 12'h  0;
rom[108394] = 12'h  0;
rom[108395] = 12'h  0;
rom[108396] = 12'h  0;
rom[108397] = 12'h  0;
rom[108398] = 12'h  0;
rom[108399] = 12'h  0;
rom[108400] = 12'hfff;
rom[108401] = 12'hfff;
rom[108402] = 12'hfff;
rom[108403] = 12'hfff;
rom[108404] = 12'hfff;
rom[108405] = 12'hfff;
rom[108406] = 12'hfff;
rom[108407] = 12'hfff;
rom[108408] = 12'hfff;
rom[108409] = 12'hfff;
rom[108410] = 12'hfff;
rom[108411] = 12'hfff;
rom[108412] = 12'hfff;
rom[108413] = 12'hfff;
rom[108414] = 12'hfff;
rom[108415] = 12'hfff;
rom[108416] = 12'hfff;
rom[108417] = 12'hfff;
rom[108418] = 12'hfff;
rom[108419] = 12'hfff;
rom[108420] = 12'hfff;
rom[108421] = 12'hfff;
rom[108422] = 12'hfff;
rom[108423] = 12'hfff;
rom[108424] = 12'hfff;
rom[108425] = 12'hfff;
rom[108426] = 12'hfff;
rom[108427] = 12'hfff;
rom[108428] = 12'hfff;
rom[108429] = 12'hfff;
rom[108430] = 12'hfff;
rom[108431] = 12'hfff;
rom[108432] = 12'hfff;
rom[108433] = 12'hfff;
rom[108434] = 12'hfff;
rom[108435] = 12'hfff;
rom[108436] = 12'hfff;
rom[108437] = 12'hfff;
rom[108438] = 12'hfff;
rom[108439] = 12'hfff;
rom[108440] = 12'hfff;
rom[108441] = 12'hfff;
rom[108442] = 12'hfff;
rom[108443] = 12'hfff;
rom[108444] = 12'hfff;
rom[108445] = 12'hfff;
rom[108446] = 12'hfff;
rom[108447] = 12'hfff;
rom[108448] = 12'hfff;
rom[108449] = 12'hfff;
rom[108450] = 12'hfff;
rom[108451] = 12'hfff;
rom[108452] = 12'hfff;
rom[108453] = 12'heee;
rom[108454] = 12'heee;
rom[108455] = 12'heee;
rom[108456] = 12'heee;
rom[108457] = 12'heee;
rom[108458] = 12'heee;
rom[108459] = 12'heee;
rom[108460] = 12'heee;
rom[108461] = 12'heee;
rom[108462] = 12'heee;
rom[108463] = 12'heee;
rom[108464] = 12'heee;
rom[108465] = 12'heee;
rom[108466] = 12'hddd;
rom[108467] = 12'hddd;
rom[108468] = 12'hddd;
rom[108469] = 12'hddd;
rom[108470] = 12'hddd;
rom[108471] = 12'hddd;
rom[108472] = 12'hddd;
rom[108473] = 12'hddd;
rom[108474] = 12'heee;
rom[108475] = 12'heee;
rom[108476] = 12'heee;
rom[108477] = 12'heee;
rom[108478] = 12'hddd;
rom[108479] = 12'hddd;
rom[108480] = 12'hccc;
rom[108481] = 12'hccc;
rom[108482] = 12'hccc;
rom[108483] = 12'hccc;
rom[108484] = 12'hccc;
rom[108485] = 12'hccc;
rom[108486] = 12'hccc;
rom[108487] = 12'hccc;
rom[108488] = 12'hccc;
rom[108489] = 12'hccc;
rom[108490] = 12'heee;
rom[108491] = 12'heee;
rom[108492] = 12'heee;
rom[108493] = 12'hccc;
rom[108494] = 12'hccc;
rom[108495] = 12'hddd;
rom[108496] = 12'heee;
rom[108497] = 12'heee;
rom[108498] = 12'heee;
rom[108499] = 12'hddd;
rom[108500] = 12'hbbb;
rom[108501] = 12'hbbb;
rom[108502] = 12'hbbb;
rom[108503] = 12'hbbb;
rom[108504] = 12'haaa;
rom[108505] = 12'haaa;
rom[108506] = 12'haaa;
rom[108507] = 12'hbbb;
rom[108508] = 12'hbbb;
rom[108509] = 12'hccc;
rom[108510] = 12'hddd;
rom[108511] = 12'hfff;
rom[108512] = 12'hddd;
rom[108513] = 12'hbbb;
rom[108514] = 12'haaa;
rom[108515] = 12'haaa;
rom[108516] = 12'haaa;
rom[108517] = 12'h999;
rom[108518] = 12'h999;
rom[108519] = 12'haaa;
rom[108520] = 12'h999;
rom[108521] = 12'h999;
rom[108522] = 12'h999;
rom[108523] = 12'h999;
rom[108524] = 12'h999;
rom[108525] = 12'h999;
rom[108526] = 12'haaa;
rom[108527] = 12'haaa;
rom[108528] = 12'hbbb;
rom[108529] = 12'hccc;
rom[108530] = 12'hccc;
rom[108531] = 12'hbbb;
rom[108532] = 12'hbbb;
rom[108533] = 12'hbbb;
rom[108534] = 12'hbbb;
rom[108535] = 12'hbbb;
rom[108536] = 12'hbbb;
rom[108537] = 12'hbbb;
rom[108538] = 12'hbbb;
rom[108539] = 12'hbbb;
rom[108540] = 12'hbbb;
rom[108541] = 12'hccc;
rom[108542] = 12'hccc;
rom[108543] = 12'hccc;
rom[108544] = 12'hccc;
rom[108545] = 12'hccc;
rom[108546] = 12'hccc;
rom[108547] = 12'hddd;
rom[108548] = 12'hddd;
rom[108549] = 12'heee;
rom[108550] = 12'heee;
rom[108551] = 12'hfff;
rom[108552] = 12'hfff;
rom[108553] = 12'hfff;
rom[108554] = 12'hfff;
rom[108555] = 12'hfff;
rom[108556] = 12'hfff;
rom[108557] = 12'hfff;
rom[108558] = 12'hfff;
rom[108559] = 12'hfff;
rom[108560] = 12'hfff;
rom[108561] = 12'hfff;
rom[108562] = 12'hfff;
rom[108563] = 12'hfff;
rom[108564] = 12'hfff;
rom[108565] = 12'hfff;
rom[108566] = 12'hfff;
rom[108567] = 12'hfff;
rom[108568] = 12'hfff;
rom[108569] = 12'hfff;
rom[108570] = 12'hfff;
rom[108571] = 12'heee;
rom[108572] = 12'heee;
rom[108573] = 12'heee;
rom[108574] = 12'heee;
rom[108575] = 12'heee;
rom[108576] = 12'heee;
rom[108577] = 12'heee;
rom[108578] = 12'heee;
rom[108579] = 12'hddd;
rom[108580] = 12'hddd;
rom[108581] = 12'hddd;
rom[108582] = 12'hddd;
rom[108583] = 12'hddd;
rom[108584] = 12'hccc;
rom[108585] = 12'hccc;
rom[108586] = 12'hccc;
rom[108587] = 12'hccc;
rom[108588] = 12'hccc;
rom[108589] = 12'hccc;
rom[108590] = 12'hccc;
rom[108591] = 12'hccc;
rom[108592] = 12'hccc;
rom[108593] = 12'hccc;
rom[108594] = 12'hccc;
rom[108595] = 12'hccc;
rom[108596] = 12'hccc;
rom[108597] = 12'hccc;
rom[108598] = 12'hccc;
rom[108599] = 12'hccc;
rom[108600] = 12'hbbb;
rom[108601] = 12'hbbb;
rom[108602] = 12'hbbb;
rom[108603] = 12'hbbb;
rom[108604] = 12'hbbb;
rom[108605] = 12'hbbb;
rom[108606] = 12'hbbb;
rom[108607] = 12'hbbb;
rom[108608] = 12'hbbb;
rom[108609] = 12'hbbb;
rom[108610] = 12'hbbb;
rom[108611] = 12'hbbb;
rom[108612] = 12'hbbb;
rom[108613] = 12'hccc;
rom[108614] = 12'hccc;
rom[108615] = 12'hccc;
rom[108616] = 12'hddd;
rom[108617] = 12'hddd;
rom[108618] = 12'heee;
rom[108619] = 12'heee;
rom[108620] = 12'heee;
rom[108621] = 12'hfff;
rom[108622] = 12'hfff;
rom[108623] = 12'hfff;
rom[108624] = 12'hfff;
rom[108625] = 12'hfff;
rom[108626] = 12'hfff;
rom[108627] = 12'hfff;
rom[108628] = 12'hfff;
rom[108629] = 12'hfff;
rom[108630] = 12'hfff;
rom[108631] = 12'hfff;
rom[108632] = 12'hfff;
rom[108633] = 12'hfff;
rom[108634] = 12'hfff;
rom[108635] = 12'hfff;
rom[108636] = 12'hfff;
rom[108637] = 12'hfff;
rom[108638] = 12'hfff;
rom[108639] = 12'hfff;
rom[108640] = 12'heee;
rom[108641] = 12'hddd;
rom[108642] = 12'hccc;
rom[108643] = 12'hccc;
rom[108644] = 12'hbbb;
rom[108645] = 12'hbbb;
rom[108646] = 12'hccc;
rom[108647] = 12'hccc;
rom[108648] = 12'heee;
rom[108649] = 12'heee;
rom[108650] = 12'hddd;
rom[108651] = 12'hccc;
rom[108652] = 12'haaa;
rom[108653] = 12'h888;
rom[108654] = 12'h777;
rom[108655] = 12'h777;
rom[108656] = 12'h777;
rom[108657] = 12'h888;
rom[108658] = 12'h888;
rom[108659] = 12'h888;
rom[108660] = 12'h888;
rom[108661] = 12'haaa;
rom[108662] = 12'hddd;
rom[108663] = 12'hfff;
rom[108664] = 12'hfff;
rom[108665] = 12'hddd;
rom[108666] = 12'haaa;
rom[108667] = 12'h888;
rom[108668] = 12'h777;
rom[108669] = 12'h666;
rom[108670] = 12'h666;
rom[108671] = 12'hbbb;
rom[108672] = 12'hfff;
rom[108673] = 12'hbbb;
rom[108674] = 12'h555;
rom[108675] = 12'h333;
rom[108676] = 12'h222;
rom[108677] = 12'h222;
rom[108678] = 12'h222;
rom[108679] = 12'h222;
rom[108680] = 12'h111;
rom[108681] = 12'h  0;
rom[108682] = 12'h222;
rom[108683] = 12'h777;
rom[108684] = 12'hddd;
rom[108685] = 12'hfff;
rom[108686] = 12'hccc;
rom[108687] = 12'h999;
rom[108688] = 12'h555;
rom[108689] = 12'h555;
rom[108690] = 12'h444;
rom[108691] = 12'h333;
rom[108692] = 12'h333;
rom[108693] = 12'h222;
rom[108694] = 12'h222;
rom[108695] = 12'h222;
rom[108696] = 12'h222;
rom[108697] = 12'h222;
rom[108698] = 12'h333;
rom[108699] = 12'h777;
rom[108700] = 12'hbbb;
rom[108701] = 12'hccc;
rom[108702] = 12'hccc;
rom[108703] = 12'hbbb;
rom[108704] = 12'hddd;
rom[108705] = 12'heee;
rom[108706] = 12'hccc;
rom[108707] = 12'h888;
rom[108708] = 12'h555;
rom[108709] = 12'h333;
rom[108710] = 12'h333;
rom[108711] = 12'h222;
rom[108712] = 12'h222;
rom[108713] = 12'h222;
rom[108714] = 12'h111;
rom[108715] = 12'h111;
rom[108716] = 12'h111;
rom[108717] = 12'h111;
rom[108718] = 12'h111;
rom[108719] = 12'h111;
rom[108720] = 12'h111;
rom[108721] = 12'h111;
rom[108722] = 12'h111;
rom[108723] = 12'h111;
rom[108724] = 12'h111;
rom[108725] = 12'h111;
rom[108726] = 12'h111;
rom[108727] = 12'h111;
rom[108728] = 12'h222;
rom[108729] = 12'h222;
rom[108730] = 12'h333;
rom[108731] = 12'h333;
rom[108732] = 12'h222;
rom[108733] = 12'h111;
rom[108734] = 12'h111;
rom[108735] = 12'h  0;
rom[108736] = 12'h  0;
rom[108737] = 12'h  0;
rom[108738] = 12'h  0;
rom[108739] = 12'h  0;
rom[108740] = 12'h  0;
rom[108741] = 12'h  0;
rom[108742] = 12'h  0;
rom[108743] = 12'h  0;
rom[108744] = 12'h  0;
rom[108745] = 12'h  0;
rom[108746] = 12'h  0;
rom[108747] = 12'h  0;
rom[108748] = 12'h  0;
rom[108749] = 12'h  0;
rom[108750] = 12'h111;
rom[108751] = 12'h  0;
rom[108752] = 12'h111;
rom[108753] = 12'h222;
rom[108754] = 12'h222;
rom[108755] = 12'h333;
rom[108756] = 12'h555;
rom[108757] = 12'h999;
rom[108758] = 12'hccc;
rom[108759] = 12'heee;
rom[108760] = 12'hddd;
rom[108761] = 12'h999;
rom[108762] = 12'h555;
rom[108763] = 12'h444;
rom[108764] = 12'h333;
rom[108765] = 12'h333;
rom[108766] = 12'h222;
rom[108767] = 12'h111;
rom[108768] = 12'h111;
rom[108769] = 12'h111;
rom[108770] = 12'h111;
rom[108771] = 12'h  0;
rom[108772] = 12'h  0;
rom[108773] = 12'h  0;
rom[108774] = 12'h  0;
rom[108775] = 12'h  0;
rom[108776] = 12'h  0;
rom[108777] = 12'h  0;
rom[108778] = 12'h  0;
rom[108779] = 12'h  0;
rom[108780] = 12'h  0;
rom[108781] = 12'h  0;
rom[108782] = 12'h  0;
rom[108783] = 12'h  0;
rom[108784] = 12'h  0;
rom[108785] = 12'h  0;
rom[108786] = 12'h  0;
rom[108787] = 12'h  0;
rom[108788] = 12'h  0;
rom[108789] = 12'h  0;
rom[108790] = 12'h  0;
rom[108791] = 12'h  0;
rom[108792] = 12'h  0;
rom[108793] = 12'h  0;
rom[108794] = 12'h  0;
rom[108795] = 12'h  0;
rom[108796] = 12'h  0;
rom[108797] = 12'h  0;
rom[108798] = 12'h  0;
rom[108799] = 12'h  0;
rom[108800] = 12'hfff;
rom[108801] = 12'hfff;
rom[108802] = 12'hfff;
rom[108803] = 12'hfff;
rom[108804] = 12'hfff;
rom[108805] = 12'hfff;
rom[108806] = 12'hfff;
rom[108807] = 12'hfff;
rom[108808] = 12'hfff;
rom[108809] = 12'hfff;
rom[108810] = 12'hfff;
rom[108811] = 12'hfff;
rom[108812] = 12'hfff;
rom[108813] = 12'hfff;
rom[108814] = 12'hfff;
rom[108815] = 12'hfff;
rom[108816] = 12'hfff;
rom[108817] = 12'hfff;
rom[108818] = 12'hfff;
rom[108819] = 12'hfff;
rom[108820] = 12'hfff;
rom[108821] = 12'hfff;
rom[108822] = 12'hfff;
rom[108823] = 12'hfff;
rom[108824] = 12'hfff;
rom[108825] = 12'hfff;
rom[108826] = 12'hfff;
rom[108827] = 12'hfff;
rom[108828] = 12'hfff;
rom[108829] = 12'hfff;
rom[108830] = 12'hfff;
rom[108831] = 12'hfff;
rom[108832] = 12'hfff;
rom[108833] = 12'hfff;
rom[108834] = 12'hfff;
rom[108835] = 12'hfff;
rom[108836] = 12'hfff;
rom[108837] = 12'hfff;
rom[108838] = 12'hfff;
rom[108839] = 12'hfff;
rom[108840] = 12'hfff;
rom[108841] = 12'hfff;
rom[108842] = 12'hfff;
rom[108843] = 12'hfff;
rom[108844] = 12'hfff;
rom[108845] = 12'hfff;
rom[108846] = 12'hfff;
rom[108847] = 12'hfff;
rom[108848] = 12'hfff;
rom[108849] = 12'hfff;
rom[108850] = 12'hfff;
rom[108851] = 12'heee;
rom[108852] = 12'heee;
rom[108853] = 12'heee;
rom[108854] = 12'hfff;
rom[108855] = 12'hfff;
rom[108856] = 12'heee;
rom[108857] = 12'heee;
rom[108858] = 12'heee;
rom[108859] = 12'heee;
rom[108860] = 12'heee;
rom[108861] = 12'heee;
rom[108862] = 12'heee;
rom[108863] = 12'heee;
rom[108864] = 12'hddd;
rom[108865] = 12'hddd;
rom[108866] = 12'hddd;
rom[108867] = 12'hddd;
rom[108868] = 12'hddd;
rom[108869] = 12'hddd;
rom[108870] = 12'hddd;
rom[108871] = 12'hddd;
rom[108872] = 12'hddd;
rom[108873] = 12'heee;
rom[108874] = 12'heee;
rom[108875] = 12'hddd;
rom[108876] = 12'hddd;
rom[108877] = 12'hddd;
rom[108878] = 12'hddd;
rom[108879] = 12'hccc;
rom[108880] = 12'hccc;
rom[108881] = 12'hccc;
rom[108882] = 12'hccc;
rom[108883] = 12'hccc;
rom[108884] = 12'hccc;
rom[108885] = 12'hccc;
rom[108886] = 12'hccc;
rom[108887] = 12'hccc;
rom[108888] = 12'hccc;
rom[108889] = 12'hddd;
rom[108890] = 12'heee;
rom[108891] = 12'heee;
rom[108892] = 12'hddd;
rom[108893] = 12'hccc;
rom[108894] = 12'hccc;
rom[108895] = 12'heee;
rom[108896] = 12'hfff;
rom[108897] = 12'heee;
rom[108898] = 12'hccc;
rom[108899] = 12'hbbb;
rom[108900] = 12'hbbb;
rom[108901] = 12'hbbb;
rom[108902] = 12'hbbb;
rom[108903] = 12'hbbb;
rom[108904] = 12'haaa;
rom[108905] = 12'haaa;
rom[108906] = 12'haaa;
rom[108907] = 12'hbbb;
rom[108908] = 12'hccc;
rom[108909] = 12'hddd;
rom[108910] = 12'heee;
rom[108911] = 12'heee;
rom[108912] = 12'hbbb;
rom[108913] = 12'haaa;
rom[108914] = 12'haaa;
rom[108915] = 12'haaa;
rom[108916] = 12'h999;
rom[108917] = 12'h999;
rom[108918] = 12'h999;
rom[108919] = 12'h999;
rom[108920] = 12'h999;
rom[108921] = 12'h888;
rom[108922] = 12'h888;
rom[108923] = 12'h999;
rom[108924] = 12'h999;
rom[108925] = 12'haaa;
rom[108926] = 12'haaa;
rom[108927] = 12'haaa;
rom[108928] = 12'hbbb;
rom[108929] = 12'hccc;
rom[108930] = 12'hbbb;
rom[108931] = 12'haaa;
rom[108932] = 12'haaa;
rom[108933] = 12'hbbb;
rom[108934] = 12'hbbb;
rom[108935] = 12'haaa;
rom[108936] = 12'haaa;
rom[108937] = 12'hbbb;
rom[108938] = 12'hbbb;
rom[108939] = 12'hbbb;
rom[108940] = 12'hbbb;
rom[108941] = 12'hbbb;
rom[108942] = 12'hccc;
rom[108943] = 12'hbbb;
rom[108944] = 12'hbbb;
rom[108945] = 12'hccc;
rom[108946] = 12'hccc;
rom[108947] = 12'hccc;
rom[108948] = 12'hddd;
rom[108949] = 12'hddd;
rom[108950] = 12'hddd;
rom[108951] = 12'heee;
rom[108952] = 12'heee;
rom[108953] = 12'heee;
rom[108954] = 12'hfff;
rom[108955] = 12'hfff;
rom[108956] = 12'hfff;
rom[108957] = 12'hfff;
rom[108958] = 12'hfff;
rom[108959] = 12'hfff;
rom[108960] = 12'hfff;
rom[108961] = 12'hfff;
rom[108962] = 12'hfff;
rom[108963] = 12'hfff;
rom[108964] = 12'hfff;
rom[108965] = 12'hfff;
rom[108966] = 12'hfff;
rom[108967] = 12'hfff;
rom[108968] = 12'hfff;
rom[108969] = 12'hfff;
rom[108970] = 12'hfff;
rom[108971] = 12'hfff;
rom[108972] = 12'hfff;
rom[108973] = 12'heee;
rom[108974] = 12'heee;
rom[108975] = 12'heee;
rom[108976] = 12'heee;
rom[108977] = 12'heee;
rom[108978] = 12'heee;
rom[108979] = 12'hddd;
rom[108980] = 12'hddd;
rom[108981] = 12'hddd;
rom[108982] = 12'hddd;
rom[108983] = 12'hddd;
rom[108984] = 12'hccc;
rom[108985] = 12'hccc;
rom[108986] = 12'hccc;
rom[108987] = 12'hccc;
rom[108988] = 12'hccc;
rom[108989] = 12'hccc;
rom[108990] = 12'hccc;
rom[108991] = 12'hccc;
rom[108992] = 12'hccc;
rom[108993] = 12'hccc;
rom[108994] = 12'hccc;
rom[108995] = 12'hccc;
rom[108996] = 12'hccc;
rom[108997] = 12'hccc;
rom[108998] = 12'hccc;
rom[108999] = 12'hccc;
rom[109000] = 12'hccc;
rom[109001] = 12'hccc;
rom[109002] = 12'hccc;
rom[109003] = 12'hbbb;
rom[109004] = 12'hbbb;
rom[109005] = 12'hbbb;
rom[109006] = 12'hbbb;
rom[109007] = 12'hbbb;
rom[109008] = 12'hbbb;
rom[109009] = 12'hbbb;
rom[109010] = 12'hccc;
rom[109011] = 12'hccc;
rom[109012] = 12'hccc;
rom[109013] = 12'hccc;
rom[109014] = 12'hddd;
rom[109015] = 12'hddd;
rom[109016] = 12'heee;
rom[109017] = 12'heee;
rom[109018] = 12'heee;
rom[109019] = 12'heee;
rom[109020] = 12'hfff;
rom[109021] = 12'hfff;
rom[109022] = 12'hfff;
rom[109023] = 12'hfff;
rom[109024] = 12'hfff;
rom[109025] = 12'hfff;
rom[109026] = 12'hfff;
rom[109027] = 12'hfff;
rom[109028] = 12'hfff;
rom[109029] = 12'hfff;
rom[109030] = 12'hfff;
rom[109031] = 12'hfff;
rom[109032] = 12'hfff;
rom[109033] = 12'hfff;
rom[109034] = 12'hfff;
rom[109035] = 12'hfff;
rom[109036] = 12'hfff;
rom[109037] = 12'heee;
rom[109038] = 12'hddd;
rom[109039] = 12'hccc;
rom[109040] = 12'hbbb;
rom[109041] = 12'haaa;
rom[109042] = 12'haaa;
rom[109043] = 12'h999;
rom[109044] = 12'h999;
rom[109045] = 12'h999;
rom[109046] = 12'hbbb;
rom[109047] = 12'hddd;
rom[109048] = 12'heee;
rom[109049] = 12'heee;
rom[109050] = 12'hddd;
rom[109051] = 12'haaa;
rom[109052] = 12'h888;
rom[109053] = 12'h666;
rom[109054] = 12'h666;
rom[109055] = 12'h666;
rom[109056] = 12'h666;
rom[109057] = 12'h777;
rom[109058] = 12'h777;
rom[109059] = 12'h666;
rom[109060] = 12'h777;
rom[109061] = 12'h999;
rom[109062] = 12'hccc;
rom[109063] = 12'hfff;
rom[109064] = 12'hfff;
rom[109065] = 12'hddd;
rom[109066] = 12'haaa;
rom[109067] = 12'h888;
rom[109068] = 12'h777;
rom[109069] = 12'h555;
rom[109070] = 12'h555;
rom[109071] = 12'h888;
rom[109072] = 12'hfff;
rom[109073] = 12'hbbb;
rom[109074] = 12'h777;
rom[109075] = 12'h333;
rom[109076] = 12'h111;
rom[109077] = 12'h222;
rom[109078] = 12'h222;
rom[109079] = 12'h111;
rom[109080] = 12'h111;
rom[109081] = 12'h  0;
rom[109082] = 12'h111;
rom[109083] = 12'h444;
rom[109084] = 12'h999;
rom[109085] = 12'heee;
rom[109086] = 12'heee;
rom[109087] = 12'hbbb;
rom[109088] = 12'h666;
rom[109089] = 12'h555;
rom[109090] = 12'h333;
rom[109091] = 12'h333;
rom[109092] = 12'h333;
rom[109093] = 12'h222;
rom[109094] = 12'h222;
rom[109095] = 12'h222;
rom[109096] = 12'h222;
rom[109097] = 12'h222;
rom[109098] = 12'h222;
rom[109099] = 12'h444;
rom[109100] = 12'h777;
rom[109101] = 12'hbbb;
rom[109102] = 12'hccc;
rom[109103] = 12'hbbb;
rom[109104] = 12'haaa;
rom[109105] = 12'hddd;
rom[109106] = 12'hfff;
rom[109107] = 12'hccc;
rom[109108] = 12'h888;
rom[109109] = 12'h444;
rom[109110] = 12'h333;
rom[109111] = 12'h333;
rom[109112] = 12'h222;
rom[109113] = 12'h222;
rom[109114] = 12'h222;
rom[109115] = 12'h111;
rom[109116] = 12'h111;
rom[109117] = 12'h111;
rom[109118] = 12'h111;
rom[109119] = 12'h  0;
rom[109120] = 12'h111;
rom[109121] = 12'h111;
rom[109122] = 12'h  0;
rom[109123] = 12'h  0;
rom[109124] = 12'h111;
rom[109125] = 12'h111;
rom[109126] = 12'h111;
rom[109127] = 12'h111;
rom[109128] = 12'h111;
rom[109129] = 12'h222;
rom[109130] = 12'h222;
rom[109131] = 12'h222;
rom[109132] = 12'h222;
rom[109133] = 12'h111;
rom[109134] = 12'h111;
rom[109135] = 12'h111;
rom[109136] = 12'h  0;
rom[109137] = 12'h  0;
rom[109138] = 12'h  0;
rom[109139] = 12'h  0;
rom[109140] = 12'h  0;
rom[109141] = 12'h  0;
rom[109142] = 12'h  0;
rom[109143] = 12'h  0;
rom[109144] = 12'h  0;
rom[109145] = 12'h  0;
rom[109146] = 12'h  0;
rom[109147] = 12'h  0;
rom[109148] = 12'h  0;
rom[109149] = 12'h  0;
rom[109150] = 12'h  0;
rom[109151] = 12'h  0;
rom[109152] = 12'h111;
rom[109153] = 12'h111;
rom[109154] = 12'h111;
rom[109155] = 12'h333;
rom[109156] = 12'h333;
rom[109157] = 12'h555;
rom[109158] = 12'h999;
rom[109159] = 12'hddd;
rom[109160] = 12'heee;
rom[109161] = 12'hddd;
rom[109162] = 12'h999;
rom[109163] = 12'h555;
rom[109164] = 12'h444;
rom[109165] = 12'h333;
rom[109166] = 12'h222;
rom[109167] = 12'h222;
rom[109168] = 12'h111;
rom[109169] = 12'h111;
rom[109170] = 12'h111;
rom[109171] = 12'h111;
rom[109172] = 12'h111;
rom[109173] = 12'h  0;
rom[109174] = 12'h  0;
rom[109175] = 12'h  0;
rom[109176] = 12'h  0;
rom[109177] = 12'h  0;
rom[109178] = 12'h  0;
rom[109179] = 12'h  0;
rom[109180] = 12'h  0;
rom[109181] = 12'h  0;
rom[109182] = 12'h  0;
rom[109183] = 12'h  0;
rom[109184] = 12'h  0;
rom[109185] = 12'h  0;
rom[109186] = 12'h  0;
rom[109187] = 12'h  0;
rom[109188] = 12'h  0;
rom[109189] = 12'h  0;
rom[109190] = 12'h  0;
rom[109191] = 12'h  0;
rom[109192] = 12'h  0;
rom[109193] = 12'h  0;
rom[109194] = 12'h  0;
rom[109195] = 12'h  0;
rom[109196] = 12'h  0;
rom[109197] = 12'h  0;
rom[109198] = 12'h  0;
rom[109199] = 12'h  0;
rom[109200] = 12'hfff;
rom[109201] = 12'hfff;
rom[109202] = 12'hfff;
rom[109203] = 12'hfff;
rom[109204] = 12'hfff;
rom[109205] = 12'hfff;
rom[109206] = 12'hfff;
rom[109207] = 12'hfff;
rom[109208] = 12'hfff;
rom[109209] = 12'hfff;
rom[109210] = 12'hfff;
rom[109211] = 12'hfff;
rom[109212] = 12'hfff;
rom[109213] = 12'hfff;
rom[109214] = 12'hfff;
rom[109215] = 12'hfff;
rom[109216] = 12'hfff;
rom[109217] = 12'hfff;
rom[109218] = 12'hfff;
rom[109219] = 12'hfff;
rom[109220] = 12'hfff;
rom[109221] = 12'hfff;
rom[109222] = 12'hfff;
rom[109223] = 12'hfff;
rom[109224] = 12'hfff;
rom[109225] = 12'hfff;
rom[109226] = 12'hfff;
rom[109227] = 12'hfff;
rom[109228] = 12'hfff;
rom[109229] = 12'hfff;
rom[109230] = 12'hfff;
rom[109231] = 12'hfff;
rom[109232] = 12'hfff;
rom[109233] = 12'hfff;
rom[109234] = 12'hfff;
rom[109235] = 12'hfff;
rom[109236] = 12'hfff;
rom[109237] = 12'hfff;
rom[109238] = 12'hfff;
rom[109239] = 12'hfff;
rom[109240] = 12'hfff;
rom[109241] = 12'hfff;
rom[109242] = 12'hfff;
rom[109243] = 12'hfff;
rom[109244] = 12'hfff;
rom[109245] = 12'hfff;
rom[109246] = 12'hfff;
rom[109247] = 12'hfff;
rom[109248] = 12'hfff;
rom[109249] = 12'hfff;
rom[109250] = 12'hfff;
rom[109251] = 12'heee;
rom[109252] = 12'heee;
rom[109253] = 12'heee;
rom[109254] = 12'heee;
rom[109255] = 12'heee;
rom[109256] = 12'heee;
rom[109257] = 12'heee;
rom[109258] = 12'heee;
rom[109259] = 12'heee;
rom[109260] = 12'heee;
rom[109261] = 12'heee;
rom[109262] = 12'heee;
rom[109263] = 12'hddd;
rom[109264] = 12'hddd;
rom[109265] = 12'hddd;
rom[109266] = 12'hddd;
rom[109267] = 12'hddd;
rom[109268] = 12'hddd;
rom[109269] = 12'hddd;
rom[109270] = 12'hddd;
rom[109271] = 12'hddd;
rom[109272] = 12'hddd;
rom[109273] = 12'hddd;
rom[109274] = 12'hddd;
rom[109275] = 12'hddd;
rom[109276] = 12'hddd;
rom[109277] = 12'hccc;
rom[109278] = 12'hccc;
rom[109279] = 12'hccc;
rom[109280] = 12'hccc;
rom[109281] = 12'hbbb;
rom[109282] = 12'hbbb;
rom[109283] = 12'hbbb;
rom[109284] = 12'hccc;
rom[109285] = 12'hccc;
rom[109286] = 12'hccc;
rom[109287] = 12'hccc;
rom[109288] = 12'hddd;
rom[109289] = 12'hddd;
rom[109290] = 12'heee;
rom[109291] = 12'hddd;
rom[109292] = 12'hddd;
rom[109293] = 12'hddd;
rom[109294] = 12'hddd;
rom[109295] = 12'heee;
rom[109296] = 12'hddd;
rom[109297] = 12'hccc;
rom[109298] = 12'hbbb;
rom[109299] = 12'hbbb;
rom[109300] = 12'hbbb;
rom[109301] = 12'hbbb;
rom[109302] = 12'haaa;
rom[109303] = 12'haaa;
rom[109304] = 12'haaa;
rom[109305] = 12'haaa;
rom[109306] = 12'haaa;
rom[109307] = 12'haaa;
rom[109308] = 12'hccc;
rom[109309] = 12'heee;
rom[109310] = 12'heee;
rom[109311] = 12'hddd;
rom[109312] = 12'haaa;
rom[109313] = 12'haaa;
rom[109314] = 12'haaa;
rom[109315] = 12'haaa;
rom[109316] = 12'h999;
rom[109317] = 12'h999;
rom[109318] = 12'h999;
rom[109319] = 12'haaa;
rom[109320] = 12'h999;
rom[109321] = 12'h888;
rom[109322] = 12'h888;
rom[109323] = 12'h999;
rom[109324] = 12'h999;
rom[109325] = 12'haaa;
rom[109326] = 12'haaa;
rom[109327] = 12'hbbb;
rom[109328] = 12'hbbb;
rom[109329] = 12'hbbb;
rom[109330] = 12'hbbb;
rom[109331] = 12'haaa;
rom[109332] = 12'haaa;
rom[109333] = 12'hbbb;
rom[109334] = 12'hbbb;
rom[109335] = 12'haaa;
rom[109336] = 12'haaa;
rom[109337] = 12'hbbb;
rom[109338] = 12'hbbb;
rom[109339] = 12'hbbb;
rom[109340] = 12'hbbb;
rom[109341] = 12'hbbb;
rom[109342] = 12'hbbb;
rom[109343] = 12'hbbb;
rom[109344] = 12'hbbb;
rom[109345] = 12'hbbb;
rom[109346] = 12'hccc;
rom[109347] = 12'hccc;
rom[109348] = 12'hccc;
rom[109349] = 12'hccc;
rom[109350] = 12'hddd;
rom[109351] = 12'hddd;
rom[109352] = 12'heee;
rom[109353] = 12'heee;
rom[109354] = 12'heee;
rom[109355] = 12'hfff;
rom[109356] = 12'hfff;
rom[109357] = 12'hfff;
rom[109358] = 12'hfff;
rom[109359] = 12'hfff;
rom[109360] = 12'hfff;
rom[109361] = 12'hfff;
rom[109362] = 12'hfff;
rom[109363] = 12'hfff;
rom[109364] = 12'hfff;
rom[109365] = 12'hfff;
rom[109366] = 12'hfff;
rom[109367] = 12'hfff;
rom[109368] = 12'hfff;
rom[109369] = 12'hfff;
rom[109370] = 12'hfff;
rom[109371] = 12'hfff;
rom[109372] = 12'hfff;
rom[109373] = 12'hfff;
rom[109374] = 12'heee;
rom[109375] = 12'heee;
rom[109376] = 12'heee;
rom[109377] = 12'heee;
rom[109378] = 12'heee;
rom[109379] = 12'heee;
rom[109380] = 12'hddd;
rom[109381] = 12'hddd;
rom[109382] = 12'hddd;
rom[109383] = 12'hddd;
rom[109384] = 12'hddd;
rom[109385] = 12'hddd;
rom[109386] = 12'hccc;
rom[109387] = 12'hccc;
rom[109388] = 12'hccc;
rom[109389] = 12'hccc;
rom[109390] = 12'hccc;
rom[109391] = 12'hccc;
rom[109392] = 12'hccc;
rom[109393] = 12'hccc;
rom[109394] = 12'hccc;
rom[109395] = 12'hccc;
rom[109396] = 12'hccc;
rom[109397] = 12'hccc;
rom[109398] = 12'hccc;
rom[109399] = 12'hccc;
rom[109400] = 12'hccc;
rom[109401] = 12'hccc;
rom[109402] = 12'hccc;
rom[109403] = 12'hbbb;
rom[109404] = 12'hbbb;
rom[109405] = 12'hbbb;
rom[109406] = 12'hbbb;
rom[109407] = 12'hbbb;
rom[109408] = 12'hbbb;
rom[109409] = 12'hccc;
rom[109410] = 12'hccc;
rom[109411] = 12'hddd;
rom[109412] = 12'hddd;
rom[109413] = 12'hddd;
rom[109414] = 12'heee;
rom[109415] = 12'heee;
rom[109416] = 12'heee;
rom[109417] = 12'hfff;
rom[109418] = 12'hfff;
rom[109419] = 12'hfff;
rom[109420] = 12'hfff;
rom[109421] = 12'hfff;
rom[109422] = 12'hfff;
rom[109423] = 12'hfff;
rom[109424] = 12'hfff;
rom[109425] = 12'hfff;
rom[109426] = 12'hfff;
rom[109427] = 12'hfff;
rom[109428] = 12'hfff;
rom[109429] = 12'hfff;
rom[109430] = 12'hfff;
rom[109431] = 12'hfff;
rom[109432] = 12'hfff;
rom[109433] = 12'heee;
rom[109434] = 12'hddd;
rom[109435] = 12'hddd;
rom[109436] = 12'hccc;
rom[109437] = 12'hbbb;
rom[109438] = 12'haaa;
rom[109439] = 12'h999;
rom[109440] = 12'h999;
rom[109441] = 12'h999;
rom[109442] = 12'h888;
rom[109443] = 12'h888;
rom[109444] = 12'h999;
rom[109445] = 12'h999;
rom[109446] = 12'hbbb;
rom[109447] = 12'hddd;
rom[109448] = 12'hfff;
rom[109449] = 12'heee;
rom[109450] = 12'hbbb;
rom[109451] = 12'h999;
rom[109452] = 12'h777;
rom[109453] = 12'h666;
rom[109454] = 12'h555;
rom[109455] = 12'h666;
rom[109456] = 12'h555;
rom[109457] = 12'h777;
rom[109458] = 12'h777;
rom[109459] = 12'h666;
rom[109460] = 12'h666;
rom[109461] = 12'h888;
rom[109462] = 12'hbbb;
rom[109463] = 12'heee;
rom[109464] = 12'hfff;
rom[109465] = 12'hddd;
rom[109466] = 12'haaa;
rom[109467] = 12'h777;
rom[109468] = 12'h666;
rom[109469] = 12'h555;
rom[109470] = 12'h555;
rom[109471] = 12'h777;
rom[109472] = 12'heee;
rom[109473] = 12'hccc;
rom[109474] = 12'h888;
rom[109475] = 12'h333;
rom[109476] = 12'h222;
rom[109477] = 12'h222;
rom[109478] = 12'h111;
rom[109479] = 12'h  0;
rom[109480] = 12'h111;
rom[109481] = 12'h111;
rom[109482] = 12'h111;
rom[109483] = 12'h222;
rom[109484] = 12'h777;
rom[109485] = 12'hccc;
rom[109486] = 12'heee;
rom[109487] = 12'hddd;
rom[109488] = 12'h888;
rom[109489] = 12'h555;
rom[109490] = 12'h333;
rom[109491] = 12'h333;
rom[109492] = 12'h333;
rom[109493] = 12'h333;
rom[109494] = 12'h222;
rom[109495] = 12'h222;
rom[109496] = 12'h222;
rom[109497] = 12'h222;
rom[109498] = 12'h111;
rom[109499] = 12'h222;
rom[109500] = 12'h555;
rom[109501] = 12'h999;
rom[109502] = 12'hbbb;
rom[109503] = 12'hccc;
rom[109504] = 12'hbbb;
rom[109505] = 12'hccc;
rom[109506] = 12'hddd;
rom[109507] = 12'hddd;
rom[109508] = 12'hbbb;
rom[109509] = 12'h777;
rom[109510] = 12'h444;
rom[109511] = 12'h333;
rom[109512] = 12'h222;
rom[109513] = 12'h222;
rom[109514] = 12'h222;
rom[109515] = 12'h111;
rom[109516] = 12'h111;
rom[109517] = 12'h111;
rom[109518] = 12'h111;
rom[109519] = 12'h111;
rom[109520] = 12'h111;
rom[109521] = 12'h111;
rom[109522] = 12'h  0;
rom[109523] = 12'h  0;
rom[109524] = 12'h111;
rom[109525] = 12'h111;
rom[109526] = 12'h111;
rom[109527] = 12'h111;
rom[109528] = 12'h111;
rom[109529] = 12'h222;
rom[109530] = 12'h222;
rom[109531] = 12'h222;
rom[109532] = 12'h222;
rom[109533] = 12'h111;
rom[109534] = 12'h111;
rom[109535] = 12'h111;
rom[109536] = 12'h  0;
rom[109537] = 12'h  0;
rom[109538] = 12'h  0;
rom[109539] = 12'h  0;
rom[109540] = 12'h  0;
rom[109541] = 12'h  0;
rom[109542] = 12'h  0;
rom[109543] = 12'h  0;
rom[109544] = 12'h  0;
rom[109545] = 12'h  0;
rom[109546] = 12'h  0;
rom[109547] = 12'h  0;
rom[109548] = 12'h  0;
rom[109549] = 12'h  0;
rom[109550] = 12'h  0;
rom[109551] = 12'h  0;
rom[109552] = 12'h111;
rom[109553] = 12'h  0;
rom[109554] = 12'h111;
rom[109555] = 12'h222;
rom[109556] = 12'h333;
rom[109557] = 12'h333;
rom[109558] = 12'h666;
rom[109559] = 12'haaa;
rom[109560] = 12'heee;
rom[109561] = 12'heee;
rom[109562] = 12'hbbb;
rom[109563] = 12'h777;
rom[109564] = 12'h555;
rom[109565] = 12'h444;
rom[109566] = 12'h222;
rom[109567] = 12'h222;
rom[109568] = 12'h222;
rom[109569] = 12'h111;
rom[109570] = 12'h  0;
rom[109571] = 12'h  0;
rom[109572] = 12'h111;
rom[109573] = 12'h  0;
rom[109574] = 12'h  0;
rom[109575] = 12'h  0;
rom[109576] = 12'h  0;
rom[109577] = 12'h  0;
rom[109578] = 12'h  0;
rom[109579] = 12'h  0;
rom[109580] = 12'h  0;
rom[109581] = 12'h  0;
rom[109582] = 12'h  0;
rom[109583] = 12'h  0;
rom[109584] = 12'h  0;
rom[109585] = 12'h  0;
rom[109586] = 12'h  0;
rom[109587] = 12'h  0;
rom[109588] = 12'h  0;
rom[109589] = 12'h  0;
rom[109590] = 12'h  0;
rom[109591] = 12'h  0;
rom[109592] = 12'h  0;
rom[109593] = 12'h  0;
rom[109594] = 12'h  0;
rom[109595] = 12'h  0;
rom[109596] = 12'h  0;
rom[109597] = 12'h  0;
rom[109598] = 12'h  0;
rom[109599] = 12'h  0;
rom[109600] = 12'hfff;
rom[109601] = 12'hfff;
rom[109602] = 12'hfff;
rom[109603] = 12'hfff;
rom[109604] = 12'hfff;
rom[109605] = 12'hfff;
rom[109606] = 12'hfff;
rom[109607] = 12'hfff;
rom[109608] = 12'hfff;
rom[109609] = 12'hfff;
rom[109610] = 12'hfff;
rom[109611] = 12'hfff;
rom[109612] = 12'hfff;
rom[109613] = 12'hfff;
rom[109614] = 12'hfff;
rom[109615] = 12'hfff;
rom[109616] = 12'hfff;
rom[109617] = 12'hfff;
rom[109618] = 12'hfff;
rom[109619] = 12'hfff;
rom[109620] = 12'hfff;
rom[109621] = 12'hfff;
rom[109622] = 12'hfff;
rom[109623] = 12'hfff;
rom[109624] = 12'hfff;
rom[109625] = 12'hfff;
rom[109626] = 12'hfff;
rom[109627] = 12'hfff;
rom[109628] = 12'hfff;
rom[109629] = 12'hfff;
rom[109630] = 12'hfff;
rom[109631] = 12'hfff;
rom[109632] = 12'hfff;
rom[109633] = 12'hfff;
rom[109634] = 12'hfff;
rom[109635] = 12'hfff;
rom[109636] = 12'hfff;
rom[109637] = 12'hfff;
rom[109638] = 12'hfff;
rom[109639] = 12'hfff;
rom[109640] = 12'hfff;
rom[109641] = 12'hfff;
rom[109642] = 12'hfff;
rom[109643] = 12'hfff;
rom[109644] = 12'hfff;
rom[109645] = 12'hfff;
rom[109646] = 12'hfff;
rom[109647] = 12'hfff;
rom[109648] = 12'hfff;
rom[109649] = 12'hfff;
rom[109650] = 12'heee;
rom[109651] = 12'heee;
rom[109652] = 12'heee;
rom[109653] = 12'heee;
rom[109654] = 12'heee;
rom[109655] = 12'heee;
rom[109656] = 12'heee;
rom[109657] = 12'heee;
rom[109658] = 12'heee;
rom[109659] = 12'heee;
rom[109660] = 12'heee;
rom[109661] = 12'heee;
rom[109662] = 12'hddd;
rom[109663] = 12'hddd;
rom[109664] = 12'hddd;
rom[109665] = 12'hddd;
rom[109666] = 12'hddd;
rom[109667] = 12'hddd;
rom[109668] = 12'hccc;
rom[109669] = 12'hccc;
rom[109670] = 12'hccc;
rom[109671] = 12'hddd;
rom[109672] = 12'hddd;
rom[109673] = 12'hddd;
rom[109674] = 12'hddd;
rom[109675] = 12'hccc;
rom[109676] = 12'hccc;
rom[109677] = 12'hccc;
rom[109678] = 12'hccc;
rom[109679] = 12'hccc;
rom[109680] = 12'hbbb;
rom[109681] = 12'hbbb;
rom[109682] = 12'hbbb;
rom[109683] = 12'hbbb;
rom[109684] = 12'hbbb;
rom[109685] = 12'hbbb;
rom[109686] = 12'hbbb;
rom[109687] = 12'hccc;
rom[109688] = 12'heee;
rom[109689] = 12'heee;
rom[109690] = 12'hddd;
rom[109691] = 12'hccc;
rom[109692] = 12'hddd;
rom[109693] = 12'heee;
rom[109694] = 12'heee;
rom[109695] = 12'hddd;
rom[109696] = 12'hbbb;
rom[109697] = 12'hbbb;
rom[109698] = 12'haaa;
rom[109699] = 12'haaa;
rom[109700] = 12'hbbb;
rom[109701] = 12'hbbb;
rom[109702] = 12'haaa;
rom[109703] = 12'haaa;
rom[109704] = 12'haaa;
rom[109705] = 12'haaa;
rom[109706] = 12'haaa;
rom[109707] = 12'haaa;
rom[109708] = 12'hccc;
rom[109709] = 12'heee;
rom[109710] = 12'hddd;
rom[109711] = 12'hbbb;
rom[109712] = 12'haaa;
rom[109713] = 12'haaa;
rom[109714] = 12'haaa;
rom[109715] = 12'h999;
rom[109716] = 12'h999;
rom[109717] = 12'h999;
rom[109718] = 12'h999;
rom[109719] = 12'haaa;
rom[109720] = 12'h999;
rom[109721] = 12'h999;
rom[109722] = 12'h999;
rom[109723] = 12'h999;
rom[109724] = 12'h999;
rom[109725] = 12'haaa;
rom[109726] = 12'haaa;
rom[109727] = 12'hbbb;
rom[109728] = 12'hbbb;
rom[109729] = 12'haaa;
rom[109730] = 12'haaa;
rom[109731] = 12'h999;
rom[109732] = 12'haaa;
rom[109733] = 12'haaa;
rom[109734] = 12'haaa;
rom[109735] = 12'haaa;
rom[109736] = 12'haaa;
rom[109737] = 12'haaa;
rom[109738] = 12'haaa;
rom[109739] = 12'haaa;
rom[109740] = 12'haaa;
rom[109741] = 12'haaa;
rom[109742] = 12'haaa;
rom[109743] = 12'haaa;
rom[109744] = 12'haaa;
rom[109745] = 12'hbbb;
rom[109746] = 12'hbbb;
rom[109747] = 12'hbbb;
rom[109748] = 12'hbbb;
rom[109749] = 12'hccc;
rom[109750] = 12'hccc;
rom[109751] = 12'hccc;
rom[109752] = 12'hddd;
rom[109753] = 12'hddd;
rom[109754] = 12'heee;
rom[109755] = 12'heee;
rom[109756] = 12'hfff;
rom[109757] = 12'hfff;
rom[109758] = 12'hfff;
rom[109759] = 12'hfff;
rom[109760] = 12'hfff;
rom[109761] = 12'hfff;
rom[109762] = 12'hfff;
rom[109763] = 12'hfff;
rom[109764] = 12'hfff;
rom[109765] = 12'hfff;
rom[109766] = 12'hfff;
rom[109767] = 12'hfff;
rom[109768] = 12'hfff;
rom[109769] = 12'hfff;
rom[109770] = 12'hfff;
rom[109771] = 12'hfff;
rom[109772] = 12'hfff;
rom[109773] = 12'hfff;
rom[109774] = 12'hfff;
rom[109775] = 12'hfff;
rom[109776] = 12'hfff;
rom[109777] = 12'hfff;
rom[109778] = 12'heee;
rom[109779] = 12'heee;
rom[109780] = 12'heee;
rom[109781] = 12'heee;
rom[109782] = 12'hddd;
rom[109783] = 12'hddd;
rom[109784] = 12'hddd;
rom[109785] = 12'hddd;
rom[109786] = 12'hddd;
rom[109787] = 12'hddd;
rom[109788] = 12'hddd;
rom[109789] = 12'hccc;
rom[109790] = 12'hccc;
rom[109791] = 12'hccc;
rom[109792] = 12'hccc;
rom[109793] = 12'hccc;
rom[109794] = 12'hccc;
rom[109795] = 12'hccc;
rom[109796] = 12'hccc;
rom[109797] = 12'hccc;
rom[109798] = 12'hccc;
rom[109799] = 12'hccc;
rom[109800] = 12'hccc;
rom[109801] = 12'hccc;
rom[109802] = 12'hccc;
rom[109803] = 12'hccc;
rom[109804] = 12'hccc;
rom[109805] = 12'hccc;
rom[109806] = 12'hccc;
rom[109807] = 12'hccc;
rom[109808] = 12'hccc;
rom[109809] = 12'hddd;
rom[109810] = 12'hddd;
rom[109811] = 12'heee;
rom[109812] = 12'heee;
rom[109813] = 12'heee;
rom[109814] = 12'hfff;
rom[109815] = 12'hfff;
rom[109816] = 12'hfff;
rom[109817] = 12'hfff;
rom[109818] = 12'hfff;
rom[109819] = 12'hfff;
rom[109820] = 12'hfff;
rom[109821] = 12'hfff;
rom[109822] = 12'hfff;
rom[109823] = 12'hfff;
rom[109824] = 12'hfff;
rom[109825] = 12'hfff;
rom[109826] = 12'hfff;
rom[109827] = 12'hfff;
rom[109828] = 12'hfff;
rom[109829] = 12'hfff;
rom[109830] = 12'heee;
rom[109831] = 12'heee;
rom[109832] = 12'hccc;
rom[109833] = 12'hbbb;
rom[109834] = 12'haaa;
rom[109835] = 12'h999;
rom[109836] = 12'h999;
rom[109837] = 12'h888;
rom[109838] = 12'h888;
rom[109839] = 12'h888;
rom[109840] = 12'h888;
rom[109841] = 12'h888;
rom[109842] = 12'h888;
rom[109843] = 12'h888;
rom[109844] = 12'h888;
rom[109845] = 12'h999;
rom[109846] = 12'hccc;
rom[109847] = 12'heee;
rom[109848] = 12'hfff;
rom[109849] = 12'hddd;
rom[109850] = 12'haaa;
rom[109851] = 12'h777;
rom[109852] = 12'h555;
rom[109853] = 12'h555;
rom[109854] = 12'h555;
rom[109855] = 12'h555;
rom[109856] = 12'h444;
rom[109857] = 12'h666;
rom[109858] = 12'h666;
rom[109859] = 12'h555;
rom[109860] = 12'h555;
rom[109861] = 12'h666;
rom[109862] = 12'haaa;
rom[109863] = 12'hddd;
rom[109864] = 12'hfff;
rom[109865] = 12'heee;
rom[109866] = 12'haaa;
rom[109867] = 12'h777;
rom[109868] = 12'h666;
rom[109869] = 12'h444;
rom[109870] = 12'h444;
rom[109871] = 12'h555;
rom[109872] = 12'hccc;
rom[109873] = 12'hddd;
rom[109874] = 12'haaa;
rom[109875] = 12'h444;
rom[109876] = 12'h222;
rom[109877] = 12'h222;
rom[109878] = 12'h111;
rom[109879] = 12'h  0;
rom[109880] = 12'h111;
rom[109881] = 12'h222;
rom[109882] = 12'h111;
rom[109883] = 12'h  0;
rom[109884] = 12'h333;
rom[109885] = 12'haaa;
rom[109886] = 12'heee;
rom[109887] = 12'heee;
rom[109888] = 12'hbbb;
rom[109889] = 12'h777;
rom[109890] = 12'h444;
rom[109891] = 12'h333;
rom[109892] = 12'h333;
rom[109893] = 12'h333;
rom[109894] = 12'h222;
rom[109895] = 12'h111;
rom[109896] = 12'h111;
rom[109897] = 12'h111;
rom[109898] = 12'h111;
rom[109899] = 12'h111;
rom[109900] = 12'h333;
rom[109901] = 12'h555;
rom[109902] = 12'h999;
rom[109903] = 12'hbbb;
rom[109904] = 12'hccc;
rom[109905] = 12'hbbb;
rom[109906] = 12'hccc;
rom[109907] = 12'hddd;
rom[109908] = 12'hddd;
rom[109909] = 12'haaa;
rom[109910] = 12'h666;
rom[109911] = 12'h333;
rom[109912] = 12'h222;
rom[109913] = 12'h222;
rom[109914] = 12'h222;
rom[109915] = 12'h111;
rom[109916] = 12'h111;
rom[109917] = 12'h111;
rom[109918] = 12'h111;
rom[109919] = 12'h111;
rom[109920] = 12'h111;
rom[109921] = 12'h111;
rom[109922] = 12'h111;
rom[109923] = 12'h  0;
rom[109924] = 12'h  0;
rom[109925] = 12'h111;
rom[109926] = 12'h111;
rom[109927] = 12'h111;
rom[109928] = 12'h111;
rom[109929] = 12'h111;
rom[109930] = 12'h222;
rom[109931] = 12'h222;
rom[109932] = 12'h222;
rom[109933] = 12'h111;
rom[109934] = 12'h111;
rom[109935] = 12'h111;
rom[109936] = 12'h  0;
rom[109937] = 12'h  0;
rom[109938] = 12'h  0;
rom[109939] = 12'h  0;
rom[109940] = 12'h  0;
rom[109941] = 12'h  0;
rom[109942] = 12'h  0;
rom[109943] = 12'h  0;
rom[109944] = 12'h  0;
rom[109945] = 12'h  0;
rom[109946] = 12'h  0;
rom[109947] = 12'h  0;
rom[109948] = 12'h  0;
rom[109949] = 12'h  0;
rom[109950] = 12'h  0;
rom[109951] = 12'h  0;
rom[109952] = 12'h111;
rom[109953] = 12'h  0;
rom[109954] = 12'h  0;
rom[109955] = 12'h222;
rom[109956] = 12'h222;
rom[109957] = 12'h111;
rom[109958] = 12'h333;
rom[109959] = 12'h666;
rom[109960] = 12'hbbb;
rom[109961] = 12'heee;
rom[109962] = 12'heee;
rom[109963] = 12'haaa;
rom[109964] = 12'h777;
rom[109965] = 12'h555;
rom[109966] = 12'h333;
rom[109967] = 12'h222;
rom[109968] = 12'h222;
rom[109969] = 12'h111;
rom[109970] = 12'h  0;
rom[109971] = 12'h  0;
rom[109972] = 12'h  0;
rom[109973] = 12'h  0;
rom[109974] = 12'h  0;
rom[109975] = 12'h  0;
rom[109976] = 12'h  0;
rom[109977] = 12'h  0;
rom[109978] = 12'h  0;
rom[109979] = 12'h  0;
rom[109980] = 12'h  0;
rom[109981] = 12'h  0;
rom[109982] = 12'h  0;
rom[109983] = 12'h  0;
rom[109984] = 12'h  0;
rom[109985] = 12'h  0;
rom[109986] = 12'h  0;
rom[109987] = 12'h  0;
rom[109988] = 12'h  0;
rom[109989] = 12'h  0;
rom[109990] = 12'h  0;
rom[109991] = 12'h  0;
rom[109992] = 12'h  0;
rom[109993] = 12'h  0;
rom[109994] = 12'h  0;
rom[109995] = 12'h  0;
rom[109996] = 12'h  0;
rom[109997] = 12'h  0;
rom[109998] = 12'h  0;
rom[109999] = 12'h  0;
rom[110000] = 12'hfff;
rom[110001] = 12'hfff;
rom[110002] = 12'hfff;
rom[110003] = 12'hfff;
rom[110004] = 12'hfff;
rom[110005] = 12'hfff;
rom[110006] = 12'hfff;
rom[110007] = 12'hfff;
rom[110008] = 12'hfff;
rom[110009] = 12'hfff;
rom[110010] = 12'hfff;
rom[110011] = 12'hfff;
rom[110012] = 12'hfff;
rom[110013] = 12'hfff;
rom[110014] = 12'hfff;
rom[110015] = 12'hfff;
rom[110016] = 12'hfff;
rom[110017] = 12'hfff;
rom[110018] = 12'hfff;
rom[110019] = 12'hfff;
rom[110020] = 12'hfff;
rom[110021] = 12'hfff;
rom[110022] = 12'hfff;
rom[110023] = 12'hfff;
rom[110024] = 12'hfff;
rom[110025] = 12'hfff;
rom[110026] = 12'hfff;
rom[110027] = 12'hfff;
rom[110028] = 12'hfff;
rom[110029] = 12'hfff;
rom[110030] = 12'hfff;
rom[110031] = 12'hfff;
rom[110032] = 12'hfff;
rom[110033] = 12'hfff;
rom[110034] = 12'hfff;
rom[110035] = 12'hfff;
rom[110036] = 12'hfff;
rom[110037] = 12'hfff;
rom[110038] = 12'hfff;
rom[110039] = 12'hfff;
rom[110040] = 12'hfff;
rom[110041] = 12'hfff;
rom[110042] = 12'hfff;
rom[110043] = 12'hfff;
rom[110044] = 12'hfff;
rom[110045] = 12'hfff;
rom[110046] = 12'hfff;
rom[110047] = 12'heee;
rom[110048] = 12'hfff;
rom[110049] = 12'hfff;
rom[110050] = 12'heee;
rom[110051] = 12'heee;
rom[110052] = 12'heee;
rom[110053] = 12'heee;
rom[110054] = 12'heee;
rom[110055] = 12'heee;
rom[110056] = 12'heee;
rom[110057] = 12'heee;
rom[110058] = 12'heee;
rom[110059] = 12'hddd;
rom[110060] = 12'hddd;
rom[110061] = 12'hddd;
rom[110062] = 12'hddd;
rom[110063] = 12'hddd;
rom[110064] = 12'hccc;
rom[110065] = 12'hccc;
rom[110066] = 12'hccc;
rom[110067] = 12'hccc;
rom[110068] = 12'hccc;
rom[110069] = 12'hccc;
rom[110070] = 12'hddd;
rom[110071] = 12'hddd;
rom[110072] = 12'hddd;
rom[110073] = 12'hddd;
rom[110074] = 12'hccc;
rom[110075] = 12'hccc;
rom[110076] = 12'hccc;
rom[110077] = 12'hccc;
rom[110078] = 12'hccc;
rom[110079] = 12'hbbb;
rom[110080] = 12'hbbb;
rom[110081] = 12'hbbb;
rom[110082] = 12'hbbb;
rom[110083] = 12'hbbb;
rom[110084] = 12'hbbb;
rom[110085] = 12'hbbb;
rom[110086] = 12'hccc;
rom[110087] = 12'hddd;
rom[110088] = 12'heee;
rom[110089] = 12'heee;
rom[110090] = 12'hddd;
rom[110091] = 12'hddd;
rom[110092] = 12'heee;
rom[110093] = 12'heee;
rom[110094] = 12'heee;
rom[110095] = 12'hccc;
rom[110096] = 12'hbbb;
rom[110097] = 12'haaa;
rom[110098] = 12'haaa;
rom[110099] = 12'haaa;
rom[110100] = 12'hbbb;
rom[110101] = 12'haaa;
rom[110102] = 12'haaa;
rom[110103] = 12'haaa;
rom[110104] = 12'h999;
rom[110105] = 12'haaa;
rom[110106] = 12'hbbb;
rom[110107] = 12'hbbb;
rom[110108] = 12'hddd;
rom[110109] = 12'heee;
rom[110110] = 12'hccc;
rom[110111] = 12'haaa;
rom[110112] = 12'h999;
rom[110113] = 12'h999;
rom[110114] = 12'h999;
rom[110115] = 12'h999;
rom[110116] = 12'h999;
rom[110117] = 12'h999;
rom[110118] = 12'h999;
rom[110119] = 12'h999;
rom[110120] = 12'h999;
rom[110121] = 12'h999;
rom[110122] = 12'h999;
rom[110123] = 12'h999;
rom[110124] = 12'h999;
rom[110125] = 12'haaa;
rom[110126] = 12'hbbb;
rom[110127] = 12'hbbb;
rom[110128] = 12'haaa;
rom[110129] = 12'haaa;
rom[110130] = 12'h999;
rom[110131] = 12'h999;
rom[110132] = 12'haaa;
rom[110133] = 12'haaa;
rom[110134] = 12'haaa;
rom[110135] = 12'haaa;
rom[110136] = 12'haaa;
rom[110137] = 12'haaa;
rom[110138] = 12'haaa;
rom[110139] = 12'h999;
rom[110140] = 12'h999;
rom[110141] = 12'h999;
rom[110142] = 12'h999;
rom[110143] = 12'h999;
rom[110144] = 12'haaa;
rom[110145] = 12'haaa;
rom[110146] = 12'hbbb;
rom[110147] = 12'hbbb;
rom[110148] = 12'hbbb;
rom[110149] = 12'hbbb;
rom[110150] = 12'hbbb;
rom[110151] = 12'hbbb;
rom[110152] = 12'hccc;
rom[110153] = 12'hccc;
rom[110154] = 12'hddd;
rom[110155] = 12'hddd;
rom[110156] = 12'heee;
rom[110157] = 12'heee;
rom[110158] = 12'hfff;
rom[110159] = 12'hfff;
rom[110160] = 12'hfff;
rom[110161] = 12'hfff;
rom[110162] = 12'hfff;
rom[110163] = 12'hfff;
rom[110164] = 12'hfff;
rom[110165] = 12'hfff;
rom[110166] = 12'hfff;
rom[110167] = 12'hfff;
rom[110168] = 12'hfff;
rom[110169] = 12'hfff;
rom[110170] = 12'hfff;
rom[110171] = 12'hfff;
rom[110172] = 12'hfff;
rom[110173] = 12'hfff;
rom[110174] = 12'hfff;
rom[110175] = 12'hfff;
rom[110176] = 12'hfff;
rom[110177] = 12'hfff;
rom[110178] = 12'hfff;
rom[110179] = 12'hfff;
rom[110180] = 12'heee;
rom[110181] = 12'heee;
rom[110182] = 12'heee;
rom[110183] = 12'heee;
rom[110184] = 12'hddd;
rom[110185] = 12'hddd;
rom[110186] = 12'hddd;
rom[110187] = 12'hddd;
rom[110188] = 12'hddd;
rom[110189] = 12'hddd;
rom[110190] = 12'hccc;
rom[110191] = 12'hccc;
rom[110192] = 12'hccc;
rom[110193] = 12'hccc;
rom[110194] = 12'hccc;
rom[110195] = 12'hccc;
rom[110196] = 12'hccc;
rom[110197] = 12'hccc;
rom[110198] = 12'hccc;
rom[110199] = 12'hccc;
rom[110200] = 12'hccc;
rom[110201] = 12'hccc;
rom[110202] = 12'hccc;
rom[110203] = 12'hccc;
rom[110204] = 12'hddd;
rom[110205] = 12'hddd;
rom[110206] = 12'hddd;
rom[110207] = 12'hddd;
rom[110208] = 12'heee;
rom[110209] = 12'heee;
rom[110210] = 12'heee;
rom[110211] = 12'hfff;
rom[110212] = 12'hfff;
rom[110213] = 12'hfff;
rom[110214] = 12'hfff;
rom[110215] = 12'hfff;
rom[110216] = 12'hfff;
rom[110217] = 12'hfff;
rom[110218] = 12'hfff;
rom[110219] = 12'hfff;
rom[110220] = 12'hfff;
rom[110221] = 12'hfff;
rom[110222] = 12'hfff;
rom[110223] = 12'hfff;
rom[110224] = 12'hfff;
rom[110225] = 12'hfff;
rom[110226] = 12'hfff;
rom[110227] = 12'heee;
rom[110228] = 12'heee;
rom[110229] = 12'hddd;
rom[110230] = 12'hccc;
rom[110231] = 12'hbbb;
rom[110232] = 12'h999;
rom[110233] = 12'h888;
rom[110234] = 12'h888;
rom[110235] = 12'h777;
rom[110236] = 12'h777;
rom[110237] = 12'h777;
rom[110238] = 12'h777;
rom[110239] = 12'h777;
rom[110240] = 12'h888;
rom[110241] = 12'h888;
rom[110242] = 12'h888;
rom[110243] = 12'h777;
rom[110244] = 12'h888;
rom[110245] = 12'haaa;
rom[110246] = 12'hccc;
rom[110247] = 12'heee;
rom[110248] = 12'heee;
rom[110249] = 12'hbbb;
rom[110250] = 12'h888;
rom[110251] = 12'h555;
rom[110252] = 12'h444;
rom[110253] = 12'h444;
rom[110254] = 12'h444;
rom[110255] = 12'h444;
rom[110256] = 12'h444;
rom[110257] = 12'h555;
rom[110258] = 12'h555;
rom[110259] = 12'h555;
rom[110260] = 12'h444;
rom[110261] = 12'h555;
rom[110262] = 12'h888;
rom[110263] = 12'hddd;
rom[110264] = 12'hfff;
rom[110265] = 12'heee;
rom[110266] = 12'haaa;
rom[110267] = 12'h777;
rom[110268] = 12'h666;
rom[110269] = 12'h444;
rom[110270] = 12'h333;
rom[110271] = 12'h444;
rom[110272] = 12'haaa;
rom[110273] = 12'heee;
rom[110274] = 12'hbbb;
rom[110275] = 12'h555;
rom[110276] = 12'h222;
rom[110277] = 12'h222;
rom[110278] = 12'h111;
rom[110279] = 12'h111;
rom[110280] = 12'h111;
rom[110281] = 12'h111;
rom[110282] = 12'h111;
rom[110283] = 12'h  0;
rom[110284] = 12'h222;
rom[110285] = 12'h777;
rom[110286] = 12'hccc;
rom[110287] = 12'heee;
rom[110288] = 12'hddd;
rom[110289] = 12'h999;
rom[110290] = 12'h444;
rom[110291] = 12'h222;
rom[110292] = 12'h222;
rom[110293] = 12'h333;
rom[110294] = 12'h222;
rom[110295] = 12'h111;
rom[110296] = 12'h111;
rom[110297] = 12'h111;
rom[110298] = 12'h222;
rom[110299] = 12'h222;
rom[110300] = 12'h222;
rom[110301] = 12'h333;
rom[110302] = 12'h666;
rom[110303] = 12'h888;
rom[110304] = 12'hccc;
rom[110305] = 12'hbbb;
rom[110306] = 12'hbbb;
rom[110307] = 12'hddd;
rom[110308] = 12'hddd;
rom[110309] = 12'hccc;
rom[110310] = 12'h888;
rom[110311] = 12'h555;
rom[110312] = 12'h333;
rom[110313] = 12'h333;
rom[110314] = 12'h222;
rom[110315] = 12'h222;
rom[110316] = 12'h111;
rom[110317] = 12'h111;
rom[110318] = 12'h111;
rom[110319] = 12'h111;
rom[110320] = 12'h111;
rom[110321] = 12'h111;
rom[110322] = 12'h111;
rom[110323] = 12'h111;
rom[110324] = 12'h111;
rom[110325] = 12'h111;
rom[110326] = 12'h111;
rom[110327] = 12'h111;
rom[110328] = 12'h111;
rom[110329] = 12'h111;
rom[110330] = 12'h111;
rom[110331] = 12'h111;
rom[110332] = 12'h111;
rom[110333] = 12'h111;
rom[110334] = 12'h111;
rom[110335] = 12'h111;
rom[110336] = 12'h  0;
rom[110337] = 12'h  0;
rom[110338] = 12'h  0;
rom[110339] = 12'h  0;
rom[110340] = 12'h  0;
rom[110341] = 12'h  0;
rom[110342] = 12'h  0;
rom[110343] = 12'h  0;
rom[110344] = 12'h  0;
rom[110345] = 12'h  0;
rom[110346] = 12'h  0;
rom[110347] = 12'h  0;
rom[110348] = 12'h  0;
rom[110349] = 12'h  0;
rom[110350] = 12'h  0;
rom[110351] = 12'h  0;
rom[110352] = 12'h  0;
rom[110353] = 12'h  0;
rom[110354] = 12'h  0;
rom[110355] = 12'h111;
rom[110356] = 12'h111;
rom[110357] = 12'h111;
rom[110358] = 12'h222;
rom[110359] = 12'h444;
rom[110360] = 12'h777;
rom[110361] = 12'hbbb;
rom[110362] = 12'heee;
rom[110363] = 12'hddd;
rom[110364] = 12'h999;
rom[110365] = 12'h666;
rom[110366] = 12'h444;
rom[110367] = 12'h333;
rom[110368] = 12'h222;
rom[110369] = 12'h222;
rom[110370] = 12'h111;
rom[110371] = 12'h111;
rom[110372] = 12'h  0;
rom[110373] = 12'h  0;
rom[110374] = 12'h  0;
rom[110375] = 12'h  0;
rom[110376] = 12'h  0;
rom[110377] = 12'h  0;
rom[110378] = 12'h  0;
rom[110379] = 12'h  0;
rom[110380] = 12'h  0;
rom[110381] = 12'h  0;
rom[110382] = 12'h  0;
rom[110383] = 12'h  0;
rom[110384] = 12'h  0;
rom[110385] = 12'h  0;
rom[110386] = 12'h  0;
rom[110387] = 12'h  0;
rom[110388] = 12'h  0;
rom[110389] = 12'h  0;
rom[110390] = 12'h  0;
rom[110391] = 12'h  0;
rom[110392] = 12'h  0;
rom[110393] = 12'h  0;
rom[110394] = 12'h  0;
rom[110395] = 12'h  0;
rom[110396] = 12'h  0;
rom[110397] = 12'h  0;
rom[110398] = 12'h  0;
rom[110399] = 12'h  0;
rom[110400] = 12'hfff;
rom[110401] = 12'hfff;
rom[110402] = 12'hfff;
rom[110403] = 12'hfff;
rom[110404] = 12'hfff;
rom[110405] = 12'hfff;
rom[110406] = 12'hfff;
rom[110407] = 12'hfff;
rom[110408] = 12'hfff;
rom[110409] = 12'hfff;
rom[110410] = 12'hfff;
rom[110411] = 12'hfff;
rom[110412] = 12'hfff;
rom[110413] = 12'hfff;
rom[110414] = 12'hfff;
rom[110415] = 12'hfff;
rom[110416] = 12'hfff;
rom[110417] = 12'hfff;
rom[110418] = 12'hfff;
rom[110419] = 12'hfff;
rom[110420] = 12'hfff;
rom[110421] = 12'hfff;
rom[110422] = 12'hfff;
rom[110423] = 12'hfff;
rom[110424] = 12'hfff;
rom[110425] = 12'hfff;
rom[110426] = 12'hfff;
rom[110427] = 12'hfff;
rom[110428] = 12'hfff;
rom[110429] = 12'hfff;
rom[110430] = 12'hfff;
rom[110431] = 12'hfff;
rom[110432] = 12'hfff;
rom[110433] = 12'hfff;
rom[110434] = 12'hfff;
rom[110435] = 12'hfff;
rom[110436] = 12'hfff;
rom[110437] = 12'hfff;
rom[110438] = 12'hfff;
rom[110439] = 12'hfff;
rom[110440] = 12'hfff;
rom[110441] = 12'hfff;
rom[110442] = 12'hfff;
rom[110443] = 12'hfff;
rom[110444] = 12'hfff;
rom[110445] = 12'hfff;
rom[110446] = 12'hfff;
rom[110447] = 12'heee;
rom[110448] = 12'heee;
rom[110449] = 12'heee;
rom[110450] = 12'heee;
rom[110451] = 12'heee;
rom[110452] = 12'heee;
rom[110453] = 12'heee;
rom[110454] = 12'heee;
rom[110455] = 12'heee;
rom[110456] = 12'hddd;
rom[110457] = 12'hddd;
rom[110458] = 12'hddd;
rom[110459] = 12'hddd;
rom[110460] = 12'hddd;
rom[110461] = 12'hddd;
rom[110462] = 12'hddd;
rom[110463] = 12'hddd;
rom[110464] = 12'hccc;
rom[110465] = 12'hccc;
rom[110466] = 12'hccc;
rom[110467] = 12'hccc;
rom[110468] = 12'hccc;
rom[110469] = 12'hccc;
rom[110470] = 12'hddd;
rom[110471] = 12'hddd;
rom[110472] = 12'hddd;
rom[110473] = 12'hddd;
rom[110474] = 12'hccc;
rom[110475] = 12'hccc;
rom[110476] = 12'hccc;
rom[110477] = 12'hccc;
rom[110478] = 12'hbbb;
rom[110479] = 12'hbbb;
rom[110480] = 12'hbbb;
rom[110481] = 12'hbbb;
rom[110482] = 12'hbbb;
rom[110483] = 12'hbbb;
rom[110484] = 12'hbbb;
rom[110485] = 12'hbbb;
rom[110486] = 12'hddd;
rom[110487] = 12'heee;
rom[110488] = 12'heee;
rom[110489] = 12'hddd;
rom[110490] = 12'hddd;
rom[110491] = 12'heee;
rom[110492] = 12'hfff;
rom[110493] = 12'heee;
rom[110494] = 12'hccc;
rom[110495] = 12'hbbb;
rom[110496] = 12'hbbb;
rom[110497] = 12'haaa;
rom[110498] = 12'haaa;
rom[110499] = 12'haaa;
rom[110500] = 12'haaa;
rom[110501] = 12'haaa;
rom[110502] = 12'haaa;
rom[110503] = 12'haaa;
rom[110504] = 12'h999;
rom[110505] = 12'haaa;
rom[110506] = 12'hbbb;
rom[110507] = 12'hddd;
rom[110508] = 12'hddd;
rom[110509] = 12'hccc;
rom[110510] = 12'hbbb;
rom[110511] = 12'haaa;
rom[110512] = 12'h999;
rom[110513] = 12'h999;
rom[110514] = 12'h999;
rom[110515] = 12'h999;
rom[110516] = 12'h999;
rom[110517] = 12'h999;
rom[110518] = 12'h999;
rom[110519] = 12'h999;
rom[110520] = 12'h999;
rom[110521] = 12'h999;
rom[110522] = 12'h999;
rom[110523] = 12'h999;
rom[110524] = 12'h999;
rom[110525] = 12'haaa;
rom[110526] = 12'haaa;
rom[110527] = 12'hbbb;
rom[110528] = 12'haaa;
rom[110529] = 12'h999;
rom[110530] = 12'h999;
rom[110531] = 12'haaa;
rom[110532] = 12'haaa;
rom[110533] = 12'h999;
rom[110534] = 12'h999;
rom[110535] = 12'h999;
rom[110536] = 12'haaa;
rom[110537] = 12'h999;
rom[110538] = 12'h999;
rom[110539] = 12'h999;
rom[110540] = 12'h888;
rom[110541] = 12'h888;
rom[110542] = 12'h999;
rom[110543] = 12'h999;
rom[110544] = 12'haaa;
rom[110545] = 12'haaa;
rom[110546] = 12'haaa;
rom[110547] = 12'haaa;
rom[110548] = 12'haaa;
rom[110549] = 12'haaa;
rom[110550] = 12'haaa;
rom[110551] = 12'haaa;
rom[110552] = 12'hbbb;
rom[110553] = 12'hbbb;
rom[110554] = 12'hbbb;
rom[110555] = 12'hccc;
rom[110556] = 12'hddd;
rom[110557] = 12'hddd;
rom[110558] = 12'heee;
rom[110559] = 12'heee;
rom[110560] = 12'hfff;
rom[110561] = 12'hfff;
rom[110562] = 12'hfff;
rom[110563] = 12'hfff;
rom[110564] = 12'hfff;
rom[110565] = 12'hfff;
rom[110566] = 12'hfff;
rom[110567] = 12'hfff;
rom[110568] = 12'hfff;
rom[110569] = 12'hfff;
rom[110570] = 12'hfff;
rom[110571] = 12'hfff;
rom[110572] = 12'hfff;
rom[110573] = 12'hfff;
rom[110574] = 12'hfff;
rom[110575] = 12'hfff;
rom[110576] = 12'hfff;
rom[110577] = 12'hfff;
rom[110578] = 12'hfff;
rom[110579] = 12'hfff;
rom[110580] = 12'hfff;
rom[110581] = 12'hfff;
rom[110582] = 12'hfff;
rom[110583] = 12'hfff;
rom[110584] = 12'heee;
rom[110585] = 12'heee;
rom[110586] = 12'heee;
rom[110587] = 12'heee;
rom[110588] = 12'heee;
rom[110589] = 12'heee;
rom[110590] = 12'hddd;
rom[110591] = 12'hddd;
rom[110592] = 12'hddd;
rom[110593] = 12'hddd;
rom[110594] = 12'hddd;
rom[110595] = 12'hddd;
rom[110596] = 12'hddd;
rom[110597] = 12'hddd;
rom[110598] = 12'hddd;
rom[110599] = 12'hddd;
rom[110600] = 12'hddd;
rom[110601] = 12'hddd;
rom[110602] = 12'hddd;
rom[110603] = 12'heee;
rom[110604] = 12'heee;
rom[110605] = 12'heee;
rom[110606] = 12'heee;
rom[110607] = 12'heee;
rom[110608] = 12'hfff;
rom[110609] = 12'hfff;
rom[110610] = 12'hfff;
rom[110611] = 12'hfff;
rom[110612] = 12'hfff;
rom[110613] = 12'hfff;
rom[110614] = 12'hfff;
rom[110615] = 12'hfff;
rom[110616] = 12'hfff;
rom[110617] = 12'hfff;
rom[110618] = 12'hfff;
rom[110619] = 12'hfff;
rom[110620] = 12'hfff;
rom[110621] = 12'hfff;
rom[110622] = 12'hfff;
rom[110623] = 12'hfff;
rom[110624] = 12'hfff;
rom[110625] = 12'heee;
rom[110626] = 12'hddd;
rom[110627] = 12'hccc;
rom[110628] = 12'hbbb;
rom[110629] = 12'haaa;
rom[110630] = 12'h999;
rom[110631] = 12'h888;
rom[110632] = 12'h777;
rom[110633] = 12'h777;
rom[110634] = 12'h666;
rom[110635] = 12'h666;
rom[110636] = 12'h666;
rom[110637] = 12'h666;
rom[110638] = 12'h666;
rom[110639] = 12'h666;
rom[110640] = 12'h666;
rom[110641] = 12'h777;
rom[110642] = 12'h777;
rom[110643] = 12'h666;
rom[110644] = 12'h777;
rom[110645] = 12'haaa;
rom[110646] = 12'hddd;
rom[110647] = 12'heee;
rom[110648] = 12'hddd;
rom[110649] = 12'h999;
rom[110650] = 12'h666;
rom[110651] = 12'h444;
rom[110652] = 12'h333;
rom[110653] = 12'h333;
rom[110654] = 12'h444;
rom[110655] = 12'h333;
rom[110656] = 12'h333;
rom[110657] = 12'h444;
rom[110658] = 12'h555;
rom[110659] = 12'h555;
rom[110660] = 12'h444;
rom[110661] = 12'h444;
rom[110662] = 12'h777;
rom[110663] = 12'hccc;
rom[110664] = 12'hfff;
rom[110665] = 12'heee;
rom[110666] = 12'haaa;
rom[110667] = 12'h666;
rom[110668] = 12'h555;
rom[110669] = 12'h444;
rom[110670] = 12'h333;
rom[110671] = 12'h333;
rom[110672] = 12'h888;
rom[110673] = 12'heee;
rom[110674] = 12'hddd;
rom[110675] = 12'h666;
rom[110676] = 12'h222;
rom[110677] = 12'h111;
rom[110678] = 12'h111;
rom[110679] = 12'h111;
rom[110680] = 12'h  0;
rom[110681] = 12'h  0;
rom[110682] = 12'h  0;
rom[110683] = 12'h  0;
rom[110684] = 12'h111;
rom[110685] = 12'h444;
rom[110686] = 12'h999;
rom[110687] = 12'heee;
rom[110688] = 12'hfff;
rom[110689] = 12'hbbb;
rom[110690] = 12'h666;
rom[110691] = 12'h333;
rom[110692] = 12'h222;
rom[110693] = 12'h222;
rom[110694] = 12'h222;
rom[110695] = 12'h222;
rom[110696] = 12'h111;
rom[110697] = 12'h111;
rom[110698] = 12'h222;
rom[110699] = 12'h222;
rom[110700] = 12'h111;
rom[110701] = 12'h111;
rom[110702] = 12'h333;
rom[110703] = 12'h666;
rom[110704] = 12'haaa;
rom[110705] = 12'hbbb;
rom[110706] = 12'hccc;
rom[110707] = 12'hccc;
rom[110708] = 12'hddd;
rom[110709] = 12'hccc;
rom[110710] = 12'haaa;
rom[110711] = 12'h777;
rom[110712] = 12'h444;
rom[110713] = 12'h333;
rom[110714] = 12'h222;
rom[110715] = 12'h222;
rom[110716] = 12'h222;
rom[110717] = 12'h111;
rom[110718] = 12'h111;
rom[110719] = 12'h111;
rom[110720] = 12'h111;
rom[110721] = 12'h111;
rom[110722] = 12'h111;
rom[110723] = 12'h111;
rom[110724] = 12'h111;
rom[110725] = 12'h111;
rom[110726] = 12'h111;
rom[110727] = 12'h111;
rom[110728] = 12'h111;
rom[110729] = 12'h111;
rom[110730] = 12'h111;
rom[110731] = 12'h111;
rom[110732] = 12'h111;
rom[110733] = 12'h111;
rom[110734] = 12'h111;
rom[110735] = 12'h111;
rom[110736] = 12'h  0;
rom[110737] = 12'h  0;
rom[110738] = 12'h  0;
rom[110739] = 12'h  0;
rom[110740] = 12'h  0;
rom[110741] = 12'h  0;
rom[110742] = 12'h  0;
rom[110743] = 12'h  0;
rom[110744] = 12'h  0;
rom[110745] = 12'h  0;
rom[110746] = 12'h  0;
rom[110747] = 12'h  0;
rom[110748] = 12'h  0;
rom[110749] = 12'h  0;
rom[110750] = 12'h  0;
rom[110751] = 12'h  0;
rom[110752] = 12'h  0;
rom[110753] = 12'h  0;
rom[110754] = 12'h  0;
rom[110755] = 12'h  0;
rom[110756] = 12'h  0;
rom[110757] = 12'h222;
rom[110758] = 12'h222;
rom[110759] = 12'h222;
rom[110760] = 12'h444;
rom[110761] = 12'h777;
rom[110762] = 12'hccc;
rom[110763] = 12'heee;
rom[110764] = 12'hccc;
rom[110765] = 12'h888;
rom[110766] = 12'h555;
rom[110767] = 12'h333;
rom[110768] = 12'h222;
rom[110769] = 12'h222;
rom[110770] = 12'h222;
rom[110771] = 12'h111;
rom[110772] = 12'h  0;
rom[110773] = 12'h  0;
rom[110774] = 12'h  0;
rom[110775] = 12'h  0;
rom[110776] = 12'h  0;
rom[110777] = 12'h  0;
rom[110778] = 12'h  0;
rom[110779] = 12'h  0;
rom[110780] = 12'h  0;
rom[110781] = 12'h  0;
rom[110782] = 12'h  0;
rom[110783] = 12'h  0;
rom[110784] = 12'h  0;
rom[110785] = 12'h  0;
rom[110786] = 12'h  0;
rom[110787] = 12'h  0;
rom[110788] = 12'h  0;
rom[110789] = 12'h  0;
rom[110790] = 12'h  0;
rom[110791] = 12'h  0;
rom[110792] = 12'h  0;
rom[110793] = 12'h  0;
rom[110794] = 12'h  0;
rom[110795] = 12'h  0;
rom[110796] = 12'h  0;
rom[110797] = 12'h  0;
rom[110798] = 12'h  0;
rom[110799] = 12'h  0;
rom[110800] = 12'hfff;
rom[110801] = 12'hfff;
rom[110802] = 12'hfff;
rom[110803] = 12'hfff;
rom[110804] = 12'hfff;
rom[110805] = 12'hfff;
rom[110806] = 12'hfff;
rom[110807] = 12'hfff;
rom[110808] = 12'hfff;
rom[110809] = 12'hfff;
rom[110810] = 12'hfff;
rom[110811] = 12'hfff;
rom[110812] = 12'hfff;
rom[110813] = 12'hfff;
rom[110814] = 12'hfff;
rom[110815] = 12'hfff;
rom[110816] = 12'hfff;
rom[110817] = 12'hfff;
rom[110818] = 12'hfff;
rom[110819] = 12'hfff;
rom[110820] = 12'hfff;
rom[110821] = 12'hfff;
rom[110822] = 12'hfff;
rom[110823] = 12'hfff;
rom[110824] = 12'hfff;
rom[110825] = 12'hfff;
rom[110826] = 12'hfff;
rom[110827] = 12'hfff;
rom[110828] = 12'hfff;
rom[110829] = 12'hfff;
rom[110830] = 12'hfff;
rom[110831] = 12'hfff;
rom[110832] = 12'hfff;
rom[110833] = 12'hfff;
rom[110834] = 12'hfff;
rom[110835] = 12'hfff;
rom[110836] = 12'hfff;
rom[110837] = 12'hfff;
rom[110838] = 12'hfff;
rom[110839] = 12'hfff;
rom[110840] = 12'hfff;
rom[110841] = 12'hfff;
rom[110842] = 12'hfff;
rom[110843] = 12'hfff;
rom[110844] = 12'hfff;
rom[110845] = 12'hfff;
rom[110846] = 12'heee;
rom[110847] = 12'heee;
rom[110848] = 12'heee;
rom[110849] = 12'heee;
rom[110850] = 12'heee;
rom[110851] = 12'heee;
rom[110852] = 12'heee;
rom[110853] = 12'heee;
rom[110854] = 12'hddd;
rom[110855] = 12'hddd;
rom[110856] = 12'hddd;
rom[110857] = 12'hddd;
rom[110858] = 12'hddd;
rom[110859] = 12'hddd;
rom[110860] = 12'hddd;
rom[110861] = 12'hddd;
rom[110862] = 12'hccc;
rom[110863] = 12'hccc;
rom[110864] = 12'hccc;
rom[110865] = 12'hccc;
rom[110866] = 12'hccc;
rom[110867] = 12'hccc;
rom[110868] = 12'hccc;
rom[110869] = 12'hddd;
rom[110870] = 12'hddd;
rom[110871] = 12'hddd;
rom[110872] = 12'hccc;
rom[110873] = 12'hccc;
rom[110874] = 12'hccc;
rom[110875] = 12'hccc;
rom[110876] = 12'hccc;
rom[110877] = 12'hbbb;
rom[110878] = 12'hbbb;
rom[110879] = 12'hbbb;
rom[110880] = 12'hbbb;
rom[110881] = 12'hbbb;
rom[110882] = 12'hbbb;
rom[110883] = 12'hbbb;
rom[110884] = 12'hbbb;
rom[110885] = 12'hccc;
rom[110886] = 12'heee;
rom[110887] = 12'hfff;
rom[110888] = 12'heee;
rom[110889] = 12'hddd;
rom[110890] = 12'heee;
rom[110891] = 12'hfff;
rom[110892] = 12'heee;
rom[110893] = 12'hccc;
rom[110894] = 12'hbbb;
rom[110895] = 12'hbbb;
rom[110896] = 12'haaa;
rom[110897] = 12'haaa;
rom[110898] = 12'haaa;
rom[110899] = 12'haaa;
rom[110900] = 12'haaa;
rom[110901] = 12'haaa;
rom[110902] = 12'haaa;
rom[110903] = 12'h999;
rom[110904] = 12'haaa;
rom[110905] = 12'haaa;
rom[110906] = 12'hccc;
rom[110907] = 12'heee;
rom[110908] = 12'hddd;
rom[110909] = 12'hbbb;
rom[110910] = 12'haaa;
rom[110911] = 12'haaa;
rom[110912] = 12'h999;
rom[110913] = 12'h999;
rom[110914] = 12'h888;
rom[110915] = 12'h999;
rom[110916] = 12'h999;
rom[110917] = 12'h999;
rom[110918] = 12'h999;
rom[110919] = 12'h999;
rom[110920] = 12'h999;
rom[110921] = 12'h999;
rom[110922] = 12'h999;
rom[110923] = 12'h999;
rom[110924] = 12'h999;
rom[110925] = 12'haaa;
rom[110926] = 12'haaa;
rom[110927] = 12'haaa;
rom[110928] = 12'h999;
rom[110929] = 12'h999;
rom[110930] = 12'h999;
rom[110931] = 12'h999;
rom[110932] = 12'h999;
rom[110933] = 12'h999;
rom[110934] = 12'h999;
rom[110935] = 12'h999;
rom[110936] = 12'h999;
rom[110937] = 12'h999;
rom[110938] = 12'h888;
rom[110939] = 12'h888;
rom[110940] = 12'h888;
rom[110941] = 12'h888;
rom[110942] = 12'h888;
rom[110943] = 12'h999;
rom[110944] = 12'haaa;
rom[110945] = 12'haaa;
rom[110946] = 12'h999;
rom[110947] = 12'h999;
rom[110948] = 12'h999;
rom[110949] = 12'h999;
rom[110950] = 12'h999;
rom[110951] = 12'h999;
rom[110952] = 12'h999;
rom[110953] = 12'haaa;
rom[110954] = 12'haaa;
rom[110955] = 12'hbbb;
rom[110956] = 12'hbbb;
rom[110957] = 12'hccc;
rom[110958] = 12'hccc;
rom[110959] = 12'hddd;
rom[110960] = 12'heee;
rom[110961] = 12'heee;
rom[110962] = 12'hfff;
rom[110963] = 12'hfff;
rom[110964] = 12'hfff;
rom[110965] = 12'hfff;
rom[110966] = 12'hfff;
rom[110967] = 12'hfff;
rom[110968] = 12'hfff;
rom[110969] = 12'hfff;
rom[110970] = 12'hfff;
rom[110971] = 12'hfff;
rom[110972] = 12'hfff;
rom[110973] = 12'hfff;
rom[110974] = 12'hfff;
rom[110975] = 12'hfff;
rom[110976] = 12'hfff;
rom[110977] = 12'hfff;
rom[110978] = 12'hfff;
rom[110979] = 12'hfff;
rom[110980] = 12'hfff;
rom[110981] = 12'hfff;
rom[110982] = 12'hfff;
rom[110983] = 12'hfff;
rom[110984] = 12'hfff;
rom[110985] = 12'hfff;
rom[110986] = 12'hfff;
rom[110987] = 12'hfff;
rom[110988] = 12'hfff;
rom[110989] = 12'hfff;
rom[110990] = 12'heee;
rom[110991] = 12'heee;
rom[110992] = 12'heee;
rom[110993] = 12'heee;
rom[110994] = 12'heee;
rom[110995] = 12'heee;
rom[110996] = 12'heee;
rom[110997] = 12'heee;
rom[110998] = 12'heee;
rom[110999] = 12'heee;
rom[111000] = 12'heee;
rom[111001] = 12'heee;
rom[111002] = 12'heee;
rom[111003] = 12'hfff;
rom[111004] = 12'hfff;
rom[111005] = 12'hfff;
rom[111006] = 12'hfff;
rom[111007] = 12'hfff;
rom[111008] = 12'hfff;
rom[111009] = 12'hfff;
rom[111010] = 12'hfff;
rom[111011] = 12'hfff;
rom[111012] = 12'hfff;
rom[111013] = 12'hfff;
rom[111014] = 12'hfff;
rom[111015] = 12'hfff;
rom[111016] = 12'hfff;
rom[111017] = 12'hfff;
rom[111018] = 12'hfff;
rom[111019] = 12'hfff;
rom[111020] = 12'hfff;
rom[111021] = 12'hfff;
rom[111022] = 12'heee;
rom[111023] = 12'hddd;
rom[111024] = 12'hddd;
rom[111025] = 12'hccc;
rom[111026] = 12'haaa;
rom[111027] = 12'haaa;
rom[111028] = 12'h999;
rom[111029] = 12'h999;
rom[111030] = 12'h888;
rom[111031] = 12'h777;
rom[111032] = 12'h666;
rom[111033] = 12'h666;
rom[111034] = 12'h555;
rom[111035] = 12'h555;
rom[111036] = 12'h555;
rom[111037] = 12'h555;
rom[111038] = 12'h555;
rom[111039] = 12'h555;
rom[111040] = 12'h555;
rom[111041] = 12'h666;
rom[111042] = 12'h666;
rom[111043] = 12'h666;
rom[111044] = 12'h888;
rom[111045] = 12'hbbb;
rom[111046] = 12'heee;
rom[111047] = 12'heee;
rom[111048] = 12'haaa;
rom[111049] = 12'h777;
rom[111050] = 12'h444;
rom[111051] = 12'h333;
rom[111052] = 12'h222;
rom[111053] = 12'h333;
rom[111054] = 12'h333;
rom[111055] = 12'h222;
rom[111056] = 12'h333;
rom[111057] = 12'h333;
rom[111058] = 12'h444;
rom[111059] = 12'h555;
rom[111060] = 12'h444;
rom[111061] = 12'h333;
rom[111062] = 12'h666;
rom[111063] = 12'hbbb;
rom[111064] = 12'hfff;
rom[111065] = 12'heee;
rom[111066] = 12'haaa;
rom[111067] = 12'h666;
rom[111068] = 12'h555;
rom[111069] = 12'h444;
rom[111070] = 12'h333;
rom[111071] = 12'h222;
rom[111072] = 12'h666;
rom[111073] = 12'hddd;
rom[111074] = 12'heee;
rom[111075] = 12'h888;
rom[111076] = 12'h222;
rom[111077] = 12'h111;
rom[111078] = 12'h111;
rom[111079] = 12'h111;
rom[111080] = 12'h  0;
rom[111081] = 12'h  0;
rom[111082] = 12'h  0;
rom[111083] = 12'h111;
rom[111084] = 12'h  0;
rom[111085] = 12'h111;
rom[111086] = 12'h666;
rom[111087] = 12'hccc;
rom[111088] = 12'hfff;
rom[111089] = 12'hddd;
rom[111090] = 12'h888;
rom[111091] = 12'h444;
rom[111092] = 12'h222;
rom[111093] = 12'h222;
rom[111094] = 12'h222;
rom[111095] = 12'h222;
rom[111096] = 12'h222;
rom[111097] = 12'h111;
rom[111098] = 12'h111;
rom[111099] = 12'h111;
rom[111100] = 12'h111;
rom[111101] = 12'h111;
rom[111102] = 12'h222;
rom[111103] = 12'h444;
rom[111104] = 12'h666;
rom[111105] = 12'h999;
rom[111106] = 12'hccc;
rom[111107] = 12'hccc;
rom[111108] = 12'hccc;
rom[111109] = 12'hddd;
rom[111110] = 12'hbbb;
rom[111111] = 12'h999;
rom[111112] = 12'h555;
rom[111113] = 12'h444;
rom[111114] = 12'h333;
rom[111115] = 12'h333;
rom[111116] = 12'h222;
rom[111117] = 12'h222;
rom[111118] = 12'h111;
rom[111119] = 12'h111;
rom[111120] = 12'h111;
rom[111121] = 12'h111;
rom[111122] = 12'h111;
rom[111123] = 12'h111;
rom[111124] = 12'h111;
rom[111125] = 12'h111;
rom[111126] = 12'h111;
rom[111127] = 12'h111;
rom[111128] = 12'h111;
rom[111129] = 12'h111;
rom[111130] = 12'h  0;
rom[111131] = 12'h111;
rom[111132] = 12'h111;
rom[111133] = 12'h111;
rom[111134] = 12'h111;
rom[111135] = 12'h  0;
rom[111136] = 12'h  0;
rom[111137] = 12'h  0;
rom[111138] = 12'h  0;
rom[111139] = 12'h  0;
rom[111140] = 12'h  0;
rom[111141] = 12'h  0;
rom[111142] = 12'h  0;
rom[111143] = 12'h  0;
rom[111144] = 12'h  0;
rom[111145] = 12'h  0;
rom[111146] = 12'h  0;
rom[111147] = 12'h  0;
rom[111148] = 12'h  0;
rom[111149] = 12'h  0;
rom[111150] = 12'h  0;
rom[111151] = 12'h  0;
rom[111152] = 12'h  0;
rom[111153] = 12'h  0;
rom[111154] = 12'h  0;
rom[111155] = 12'h  0;
rom[111156] = 12'h  0;
rom[111157] = 12'h111;
rom[111158] = 12'h222;
rom[111159] = 12'h111;
rom[111160] = 12'h333;
rom[111161] = 12'h444;
rom[111162] = 12'h888;
rom[111163] = 12'hddd;
rom[111164] = 12'heee;
rom[111165] = 12'hccc;
rom[111166] = 12'h888;
rom[111167] = 12'h444;
rom[111168] = 12'h222;
rom[111169] = 12'h222;
rom[111170] = 12'h222;
rom[111171] = 12'h111;
rom[111172] = 12'h111;
rom[111173] = 12'h  0;
rom[111174] = 12'h  0;
rom[111175] = 12'h  0;
rom[111176] = 12'h  0;
rom[111177] = 12'h  0;
rom[111178] = 12'h  0;
rom[111179] = 12'h  0;
rom[111180] = 12'h  0;
rom[111181] = 12'h  0;
rom[111182] = 12'h  0;
rom[111183] = 12'h  0;
rom[111184] = 12'h  0;
rom[111185] = 12'h  0;
rom[111186] = 12'h  0;
rom[111187] = 12'h  0;
rom[111188] = 12'h  0;
rom[111189] = 12'h  0;
rom[111190] = 12'h  0;
rom[111191] = 12'h  0;
rom[111192] = 12'h  0;
rom[111193] = 12'h  0;
rom[111194] = 12'h  0;
rom[111195] = 12'h  0;
rom[111196] = 12'h  0;
rom[111197] = 12'h  0;
rom[111198] = 12'h  0;
rom[111199] = 12'h  0;
rom[111200] = 12'hfff;
rom[111201] = 12'hfff;
rom[111202] = 12'hfff;
rom[111203] = 12'hfff;
rom[111204] = 12'hfff;
rom[111205] = 12'hfff;
rom[111206] = 12'hfff;
rom[111207] = 12'hfff;
rom[111208] = 12'hfff;
rom[111209] = 12'hfff;
rom[111210] = 12'hfff;
rom[111211] = 12'hfff;
rom[111212] = 12'hfff;
rom[111213] = 12'hfff;
rom[111214] = 12'hfff;
rom[111215] = 12'hfff;
rom[111216] = 12'hfff;
rom[111217] = 12'hfff;
rom[111218] = 12'hfff;
rom[111219] = 12'hfff;
rom[111220] = 12'hfff;
rom[111221] = 12'hfff;
rom[111222] = 12'hfff;
rom[111223] = 12'hfff;
rom[111224] = 12'hfff;
rom[111225] = 12'hfff;
rom[111226] = 12'hfff;
rom[111227] = 12'hfff;
rom[111228] = 12'hfff;
rom[111229] = 12'hfff;
rom[111230] = 12'hfff;
rom[111231] = 12'hfff;
rom[111232] = 12'hfff;
rom[111233] = 12'hfff;
rom[111234] = 12'hfff;
rom[111235] = 12'hfff;
rom[111236] = 12'hfff;
rom[111237] = 12'hfff;
rom[111238] = 12'hfff;
rom[111239] = 12'hfff;
rom[111240] = 12'hfff;
rom[111241] = 12'hfff;
rom[111242] = 12'hfff;
rom[111243] = 12'hfff;
rom[111244] = 12'heee;
rom[111245] = 12'heee;
rom[111246] = 12'heee;
rom[111247] = 12'heee;
rom[111248] = 12'heee;
rom[111249] = 12'heee;
rom[111250] = 12'heee;
rom[111251] = 12'heee;
rom[111252] = 12'heee;
rom[111253] = 12'heee;
rom[111254] = 12'hddd;
rom[111255] = 12'hddd;
rom[111256] = 12'hddd;
rom[111257] = 12'hddd;
rom[111258] = 12'hddd;
rom[111259] = 12'hddd;
rom[111260] = 12'hccc;
rom[111261] = 12'hccc;
rom[111262] = 12'hccc;
rom[111263] = 12'hccc;
rom[111264] = 12'hccc;
rom[111265] = 12'hccc;
rom[111266] = 12'hccc;
rom[111267] = 12'hccc;
rom[111268] = 12'hddd;
rom[111269] = 12'hddd;
rom[111270] = 12'hddd;
rom[111271] = 12'hccc;
rom[111272] = 12'hccc;
rom[111273] = 12'hccc;
rom[111274] = 12'hccc;
rom[111275] = 12'hccc;
rom[111276] = 12'hccc;
rom[111277] = 12'hbbb;
rom[111278] = 12'hbbb;
rom[111279] = 12'hbbb;
rom[111280] = 12'hbbb;
rom[111281] = 12'hbbb;
rom[111282] = 12'hbbb;
rom[111283] = 12'hbbb;
rom[111284] = 12'hccc;
rom[111285] = 12'hddd;
rom[111286] = 12'heee;
rom[111287] = 12'heee;
rom[111288] = 12'hddd;
rom[111289] = 12'heee;
rom[111290] = 12'heee;
rom[111291] = 12'heee;
rom[111292] = 12'hddd;
rom[111293] = 12'hbbb;
rom[111294] = 12'haaa;
rom[111295] = 12'haaa;
rom[111296] = 12'haaa;
rom[111297] = 12'haaa;
rom[111298] = 12'haaa;
rom[111299] = 12'haaa;
rom[111300] = 12'haaa;
rom[111301] = 12'haaa;
rom[111302] = 12'haaa;
rom[111303] = 12'h999;
rom[111304] = 12'haaa;
rom[111305] = 12'hbbb;
rom[111306] = 12'hddd;
rom[111307] = 12'hddd;
rom[111308] = 12'hccc;
rom[111309] = 12'haaa;
rom[111310] = 12'h999;
rom[111311] = 12'h999;
rom[111312] = 12'h999;
rom[111313] = 12'h999;
rom[111314] = 12'h999;
rom[111315] = 12'h999;
rom[111316] = 12'h999;
rom[111317] = 12'h999;
rom[111318] = 12'h999;
rom[111319] = 12'h999;
rom[111320] = 12'h999;
rom[111321] = 12'h999;
rom[111322] = 12'h999;
rom[111323] = 12'h999;
rom[111324] = 12'h999;
rom[111325] = 12'haaa;
rom[111326] = 12'haaa;
rom[111327] = 12'h999;
rom[111328] = 12'h888;
rom[111329] = 12'h888;
rom[111330] = 12'h888;
rom[111331] = 12'h888;
rom[111332] = 12'h999;
rom[111333] = 12'h999;
rom[111334] = 12'h999;
rom[111335] = 12'h999;
rom[111336] = 12'h888;
rom[111337] = 12'h888;
rom[111338] = 12'h777;
rom[111339] = 12'h777;
rom[111340] = 12'h777;
rom[111341] = 12'h888;
rom[111342] = 12'h888;
rom[111343] = 12'h999;
rom[111344] = 12'h999;
rom[111345] = 12'h999;
rom[111346] = 12'h888;
rom[111347] = 12'h888;
rom[111348] = 12'h888;
rom[111349] = 12'h888;
rom[111350] = 12'h888;
rom[111351] = 12'h888;
rom[111352] = 12'h999;
rom[111353] = 12'h999;
rom[111354] = 12'h999;
rom[111355] = 12'haaa;
rom[111356] = 12'haaa;
rom[111357] = 12'hbbb;
rom[111358] = 12'hbbb;
rom[111359] = 12'hbbb;
rom[111360] = 12'hccc;
rom[111361] = 12'hddd;
rom[111362] = 12'hddd;
rom[111363] = 12'heee;
rom[111364] = 12'hfff;
rom[111365] = 12'hfff;
rom[111366] = 12'hfff;
rom[111367] = 12'hfff;
rom[111368] = 12'hfff;
rom[111369] = 12'hfff;
rom[111370] = 12'hfff;
rom[111371] = 12'hfff;
rom[111372] = 12'hfff;
rom[111373] = 12'hfff;
rom[111374] = 12'hfff;
rom[111375] = 12'hfff;
rom[111376] = 12'hfff;
rom[111377] = 12'hfff;
rom[111378] = 12'hfff;
rom[111379] = 12'hfff;
rom[111380] = 12'hfff;
rom[111381] = 12'hfff;
rom[111382] = 12'hfff;
rom[111383] = 12'hfff;
rom[111384] = 12'hfff;
rom[111385] = 12'hfff;
rom[111386] = 12'hfff;
rom[111387] = 12'hfff;
rom[111388] = 12'hfff;
rom[111389] = 12'hfff;
rom[111390] = 12'hfff;
rom[111391] = 12'hfff;
rom[111392] = 12'hfff;
rom[111393] = 12'hfff;
rom[111394] = 12'hfff;
rom[111395] = 12'hfff;
rom[111396] = 12'hfff;
rom[111397] = 12'hfff;
rom[111398] = 12'hfff;
rom[111399] = 12'hfff;
rom[111400] = 12'hfff;
rom[111401] = 12'hfff;
rom[111402] = 12'hfff;
rom[111403] = 12'hfff;
rom[111404] = 12'hfff;
rom[111405] = 12'hfff;
rom[111406] = 12'hfff;
rom[111407] = 12'hfff;
rom[111408] = 12'hfff;
rom[111409] = 12'hfff;
rom[111410] = 12'hfff;
rom[111411] = 12'hfff;
rom[111412] = 12'hfff;
rom[111413] = 12'hfff;
rom[111414] = 12'hfff;
rom[111415] = 12'hfff;
rom[111416] = 12'hfff;
rom[111417] = 12'hfff;
rom[111418] = 12'hfff;
rom[111419] = 12'heee;
rom[111420] = 12'heee;
rom[111421] = 12'hddd;
rom[111422] = 12'hccc;
rom[111423] = 12'hbbb;
rom[111424] = 12'haaa;
rom[111425] = 12'h999;
rom[111426] = 12'h888;
rom[111427] = 12'h777;
rom[111428] = 12'h888;
rom[111429] = 12'h888;
rom[111430] = 12'h777;
rom[111431] = 12'h777;
rom[111432] = 12'h666;
rom[111433] = 12'h555;
rom[111434] = 12'h444;
rom[111435] = 12'h444;
rom[111436] = 12'h444;
rom[111437] = 12'h444;
rom[111438] = 12'h555;
rom[111439] = 12'h555;
rom[111440] = 12'h555;
rom[111441] = 12'h666;
rom[111442] = 12'h666;
rom[111443] = 12'h666;
rom[111444] = 12'h999;
rom[111445] = 12'hddd;
rom[111446] = 12'heee;
rom[111447] = 12'hddd;
rom[111448] = 12'h888;
rom[111449] = 12'h555;
rom[111450] = 12'h333;
rom[111451] = 12'h333;
rom[111452] = 12'h222;
rom[111453] = 12'h222;
rom[111454] = 12'h333;
rom[111455] = 12'h222;
rom[111456] = 12'h222;
rom[111457] = 12'h222;
rom[111458] = 12'h333;
rom[111459] = 12'h444;
rom[111460] = 12'h444;
rom[111461] = 12'h333;
rom[111462] = 12'h555;
rom[111463] = 12'haaa;
rom[111464] = 12'hfff;
rom[111465] = 12'heee;
rom[111466] = 12'hbbb;
rom[111467] = 12'h666;
rom[111468] = 12'h444;
rom[111469] = 12'h444;
rom[111470] = 12'h333;
rom[111471] = 12'h222;
rom[111472] = 12'h555;
rom[111473] = 12'hbbb;
rom[111474] = 12'heee;
rom[111475] = 12'haaa;
rom[111476] = 12'h333;
rom[111477] = 12'h111;
rom[111478] = 12'h111;
rom[111479] = 12'h111;
rom[111480] = 12'h  0;
rom[111481] = 12'h  0;
rom[111482] = 12'h  0;
rom[111483] = 12'h  0;
rom[111484] = 12'h  0;
rom[111485] = 12'h111;
rom[111486] = 12'h444;
rom[111487] = 12'h999;
rom[111488] = 12'hddd;
rom[111489] = 12'heee;
rom[111490] = 12'hbbb;
rom[111491] = 12'h666;
rom[111492] = 12'h222;
rom[111493] = 12'h222;
rom[111494] = 12'h222;
rom[111495] = 12'h111;
rom[111496] = 12'h222;
rom[111497] = 12'h111;
rom[111498] = 12'h111;
rom[111499] = 12'h111;
rom[111500] = 12'h111;
rom[111501] = 12'h111;
rom[111502] = 12'h222;
rom[111503] = 12'h222;
rom[111504] = 12'h444;
rom[111505] = 12'h777;
rom[111506] = 12'haaa;
rom[111507] = 12'hbbb;
rom[111508] = 12'hccc;
rom[111509] = 12'hddd;
rom[111510] = 12'hccc;
rom[111511] = 12'hbbb;
rom[111512] = 12'h777;
rom[111513] = 12'h555;
rom[111514] = 12'h333;
rom[111515] = 12'h333;
rom[111516] = 12'h333;
rom[111517] = 12'h222;
rom[111518] = 12'h111;
rom[111519] = 12'h222;
rom[111520] = 12'h111;
rom[111521] = 12'h111;
rom[111522] = 12'h111;
rom[111523] = 12'h111;
rom[111524] = 12'h111;
rom[111525] = 12'h111;
rom[111526] = 12'h111;
rom[111527] = 12'h111;
rom[111528] = 12'h111;
rom[111529] = 12'h  0;
rom[111530] = 12'h  0;
rom[111531] = 12'h  0;
rom[111532] = 12'h  0;
rom[111533] = 12'h111;
rom[111534] = 12'h  0;
rom[111535] = 12'h  0;
rom[111536] = 12'h  0;
rom[111537] = 12'h  0;
rom[111538] = 12'h  0;
rom[111539] = 12'h  0;
rom[111540] = 12'h  0;
rom[111541] = 12'h  0;
rom[111542] = 12'h  0;
rom[111543] = 12'h  0;
rom[111544] = 12'h  0;
rom[111545] = 12'h  0;
rom[111546] = 12'h  0;
rom[111547] = 12'h  0;
rom[111548] = 12'h  0;
rom[111549] = 12'h  0;
rom[111550] = 12'h  0;
rom[111551] = 12'h  0;
rom[111552] = 12'h  0;
rom[111553] = 12'h  0;
rom[111554] = 12'h  0;
rom[111555] = 12'h  0;
rom[111556] = 12'h  0;
rom[111557] = 12'h  0;
rom[111558] = 12'h111;
rom[111559] = 12'h111;
rom[111560] = 12'h222;
rom[111561] = 12'h222;
rom[111562] = 12'h555;
rom[111563] = 12'h999;
rom[111564] = 12'hccc;
rom[111565] = 12'hddd;
rom[111566] = 12'haaa;
rom[111567] = 12'h666;
rom[111568] = 12'h444;
rom[111569] = 12'h333;
rom[111570] = 12'h222;
rom[111571] = 12'h222;
rom[111572] = 12'h111;
rom[111573] = 12'h111;
rom[111574] = 12'h  0;
rom[111575] = 12'h  0;
rom[111576] = 12'h  0;
rom[111577] = 12'h  0;
rom[111578] = 12'h  0;
rom[111579] = 12'h  0;
rom[111580] = 12'h  0;
rom[111581] = 12'h  0;
rom[111582] = 12'h  0;
rom[111583] = 12'h  0;
rom[111584] = 12'h  0;
rom[111585] = 12'h  0;
rom[111586] = 12'h  0;
rom[111587] = 12'h  0;
rom[111588] = 12'h  0;
rom[111589] = 12'h  0;
rom[111590] = 12'h  0;
rom[111591] = 12'h  0;
rom[111592] = 12'h  0;
rom[111593] = 12'h  0;
rom[111594] = 12'h  0;
rom[111595] = 12'h  0;
rom[111596] = 12'h  0;
rom[111597] = 12'h  0;
rom[111598] = 12'h  0;
rom[111599] = 12'h  0;
rom[111600] = 12'hfff;
rom[111601] = 12'hfff;
rom[111602] = 12'hfff;
rom[111603] = 12'hfff;
rom[111604] = 12'hfff;
rom[111605] = 12'hfff;
rom[111606] = 12'hfff;
rom[111607] = 12'hfff;
rom[111608] = 12'hfff;
rom[111609] = 12'hfff;
rom[111610] = 12'hfff;
rom[111611] = 12'hfff;
rom[111612] = 12'hfff;
rom[111613] = 12'hfff;
rom[111614] = 12'hfff;
rom[111615] = 12'hfff;
rom[111616] = 12'hfff;
rom[111617] = 12'hfff;
rom[111618] = 12'hfff;
rom[111619] = 12'hfff;
rom[111620] = 12'hfff;
rom[111621] = 12'hfff;
rom[111622] = 12'hfff;
rom[111623] = 12'hfff;
rom[111624] = 12'hfff;
rom[111625] = 12'hfff;
rom[111626] = 12'hfff;
rom[111627] = 12'hfff;
rom[111628] = 12'hfff;
rom[111629] = 12'hfff;
rom[111630] = 12'hfff;
rom[111631] = 12'hfff;
rom[111632] = 12'hfff;
rom[111633] = 12'hfff;
rom[111634] = 12'hfff;
rom[111635] = 12'hfff;
rom[111636] = 12'hfff;
rom[111637] = 12'hfff;
rom[111638] = 12'hfff;
rom[111639] = 12'hfff;
rom[111640] = 12'hfff;
rom[111641] = 12'hfff;
rom[111642] = 12'hfff;
rom[111643] = 12'heee;
rom[111644] = 12'heee;
rom[111645] = 12'heee;
rom[111646] = 12'heee;
rom[111647] = 12'heee;
rom[111648] = 12'heee;
rom[111649] = 12'heee;
rom[111650] = 12'heee;
rom[111651] = 12'heee;
rom[111652] = 12'heee;
rom[111653] = 12'heee;
rom[111654] = 12'hddd;
rom[111655] = 12'hddd;
rom[111656] = 12'hddd;
rom[111657] = 12'hddd;
rom[111658] = 12'hddd;
rom[111659] = 12'hddd;
rom[111660] = 12'hccc;
rom[111661] = 12'hccc;
rom[111662] = 12'hccc;
rom[111663] = 12'hccc;
rom[111664] = 12'hccc;
rom[111665] = 12'hccc;
rom[111666] = 12'hccc;
rom[111667] = 12'hccc;
rom[111668] = 12'hddd;
rom[111669] = 12'hddd;
rom[111670] = 12'hccc;
rom[111671] = 12'hccc;
rom[111672] = 12'hccc;
rom[111673] = 12'hccc;
rom[111674] = 12'hccc;
rom[111675] = 12'hccc;
rom[111676] = 12'hccc;
rom[111677] = 12'hbbb;
rom[111678] = 12'hbbb;
rom[111679] = 12'hbbb;
rom[111680] = 12'hbbb;
rom[111681] = 12'hbbb;
rom[111682] = 12'hbbb;
rom[111683] = 12'hbbb;
rom[111684] = 12'hccc;
rom[111685] = 12'heee;
rom[111686] = 12'heee;
rom[111687] = 12'hddd;
rom[111688] = 12'heee;
rom[111689] = 12'heee;
rom[111690] = 12'heee;
rom[111691] = 12'hddd;
rom[111692] = 12'hbbb;
rom[111693] = 12'haaa;
rom[111694] = 12'haaa;
rom[111695] = 12'haaa;
rom[111696] = 12'haaa;
rom[111697] = 12'haaa;
rom[111698] = 12'haaa;
rom[111699] = 12'haaa;
rom[111700] = 12'haaa;
rom[111701] = 12'haaa;
rom[111702] = 12'haaa;
rom[111703] = 12'haaa;
rom[111704] = 12'hbbb;
rom[111705] = 12'hccc;
rom[111706] = 12'hddd;
rom[111707] = 12'hccc;
rom[111708] = 12'hbbb;
rom[111709] = 12'haaa;
rom[111710] = 12'h999;
rom[111711] = 12'h999;
rom[111712] = 12'h999;
rom[111713] = 12'h999;
rom[111714] = 12'h999;
rom[111715] = 12'h999;
rom[111716] = 12'h999;
rom[111717] = 12'h999;
rom[111718] = 12'h999;
rom[111719] = 12'h999;
rom[111720] = 12'h999;
rom[111721] = 12'h999;
rom[111722] = 12'h999;
rom[111723] = 12'h999;
rom[111724] = 12'h999;
rom[111725] = 12'haaa;
rom[111726] = 12'h999;
rom[111727] = 12'h888;
rom[111728] = 12'h888;
rom[111729] = 12'h888;
rom[111730] = 12'h888;
rom[111731] = 12'h888;
rom[111732] = 12'h888;
rom[111733] = 12'h999;
rom[111734] = 12'h999;
rom[111735] = 12'h888;
rom[111736] = 12'h888;
rom[111737] = 12'h777;
rom[111738] = 12'h777;
rom[111739] = 12'h777;
rom[111740] = 12'h777;
rom[111741] = 12'h777;
rom[111742] = 12'h888;
rom[111743] = 12'h999;
rom[111744] = 12'h999;
rom[111745] = 12'h888;
rom[111746] = 12'h777;
rom[111747] = 12'h777;
rom[111748] = 12'h777;
rom[111749] = 12'h888;
rom[111750] = 12'h888;
rom[111751] = 12'h888;
rom[111752] = 12'h888;
rom[111753] = 12'h888;
rom[111754] = 12'h999;
rom[111755] = 12'h999;
rom[111756] = 12'h999;
rom[111757] = 12'haaa;
rom[111758] = 12'haaa;
rom[111759] = 12'hbbb;
rom[111760] = 12'hbbb;
rom[111761] = 12'hbbb;
rom[111762] = 12'hccc;
rom[111763] = 12'hddd;
rom[111764] = 12'hddd;
rom[111765] = 12'heee;
rom[111766] = 12'heee;
rom[111767] = 12'heee;
rom[111768] = 12'hfff;
rom[111769] = 12'hfff;
rom[111770] = 12'hfff;
rom[111771] = 12'hfff;
rom[111772] = 12'hfff;
rom[111773] = 12'hfff;
rom[111774] = 12'hfff;
rom[111775] = 12'hfff;
rom[111776] = 12'hfff;
rom[111777] = 12'hfff;
rom[111778] = 12'hfff;
rom[111779] = 12'hfff;
rom[111780] = 12'hfff;
rom[111781] = 12'hfff;
rom[111782] = 12'hfff;
rom[111783] = 12'hfff;
rom[111784] = 12'hfff;
rom[111785] = 12'hfff;
rom[111786] = 12'hfff;
rom[111787] = 12'hfff;
rom[111788] = 12'hfff;
rom[111789] = 12'hfff;
rom[111790] = 12'hfff;
rom[111791] = 12'hfff;
rom[111792] = 12'hfff;
rom[111793] = 12'hfff;
rom[111794] = 12'hfff;
rom[111795] = 12'hfff;
rom[111796] = 12'hfff;
rom[111797] = 12'hfff;
rom[111798] = 12'hfff;
rom[111799] = 12'hfff;
rom[111800] = 12'hfff;
rom[111801] = 12'hfff;
rom[111802] = 12'hfff;
rom[111803] = 12'hfff;
rom[111804] = 12'hfff;
rom[111805] = 12'hfff;
rom[111806] = 12'hfff;
rom[111807] = 12'hfff;
rom[111808] = 12'hfff;
rom[111809] = 12'hfff;
rom[111810] = 12'hfff;
rom[111811] = 12'hfff;
rom[111812] = 12'hfff;
rom[111813] = 12'hfff;
rom[111814] = 12'hfff;
rom[111815] = 12'hfff;
rom[111816] = 12'hfff;
rom[111817] = 12'hfff;
rom[111818] = 12'heee;
rom[111819] = 12'hddd;
rom[111820] = 12'hccc;
rom[111821] = 12'hbbb;
rom[111822] = 12'haaa;
rom[111823] = 12'h999;
rom[111824] = 12'h888;
rom[111825] = 12'h777;
rom[111826] = 12'h666;
rom[111827] = 12'h666;
rom[111828] = 12'h777;
rom[111829] = 12'h777;
rom[111830] = 12'h777;
rom[111831] = 12'h777;
rom[111832] = 12'h666;
rom[111833] = 12'h555;
rom[111834] = 12'h444;
rom[111835] = 12'h333;
rom[111836] = 12'h333;
rom[111837] = 12'h444;
rom[111838] = 12'h444;
rom[111839] = 12'h555;
rom[111840] = 12'h555;
rom[111841] = 12'h666;
rom[111842] = 12'h666;
rom[111843] = 12'h666;
rom[111844] = 12'h999;
rom[111845] = 12'hddd;
rom[111846] = 12'hddd;
rom[111847] = 12'hbbb;
rom[111848] = 12'h777;
rom[111849] = 12'h333;
rom[111850] = 12'h222;
rom[111851] = 12'h222;
rom[111852] = 12'h111;
rom[111853] = 12'h111;
rom[111854] = 12'h222;
rom[111855] = 12'h111;
rom[111856] = 12'h111;
rom[111857] = 12'h222;
rom[111858] = 12'h333;
rom[111859] = 12'h444;
rom[111860] = 12'h333;
rom[111861] = 12'h222;
rom[111862] = 12'h555;
rom[111863] = 12'h999;
rom[111864] = 12'hfff;
rom[111865] = 12'hfff;
rom[111866] = 12'hbbb;
rom[111867] = 12'h666;
rom[111868] = 12'h444;
rom[111869] = 12'h444;
rom[111870] = 12'h222;
rom[111871] = 12'h222;
rom[111872] = 12'h333;
rom[111873] = 12'haaa;
rom[111874] = 12'heee;
rom[111875] = 12'hbbb;
rom[111876] = 12'h444;
rom[111877] = 12'h111;
rom[111878] = 12'h111;
rom[111879] = 12'h111;
rom[111880] = 12'h  0;
rom[111881] = 12'h  0;
rom[111882] = 12'h111;
rom[111883] = 12'h111;
rom[111884] = 12'h  0;
rom[111885] = 12'h  0;
rom[111886] = 12'h333;
rom[111887] = 12'h777;
rom[111888] = 12'hccc;
rom[111889] = 12'heee;
rom[111890] = 12'hddd;
rom[111891] = 12'h888;
rom[111892] = 12'h333;
rom[111893] = 12'h222;
rom[111894] = 12'h222;
rom[111895] = 12'h111;
rom[111896] = 12'h111;
rom[111897] = 12'h111;
rom[111898] = 12'h111;
rom[111899] = 12'h111;
rom[111900] = 12'h111;
rom[111901] = 12'h111;
rom[111902] = 12'h111;
rom[111903] = 12'h111;
rom[111904] = 12'h333;
rom[111905] = 12'h555;
rom[111906] = 12'h888;
rom[111907] = 12'haaa;
rom[111908] = 12'hbbb;
rom[111909] = 12'hccc;
rom[111910] = 12'hccc;
rom[111911] = 12'hccc;
rom[111912] = 12'h999;
rom[111913] = 12'h666;
rom[111914] = 12'h333;
rom[111915] = 12'h333;
rom[111916] = 12'h333;
rom[111917] = 12'h222;
rom[111918] = 12'h111;
rom[111919] = 12'h222;
rom[111920] = 12'h111;
rom[111921] = 12'h111;
rom[111922] = 12'h111;
rom[111923] = 12'h111;
rom[111924] = 12'h111;
rom[111925] = 12'h111;
rom[111926] = 12'h111;
rom[111927] = 12'h111;
rom[111928] = 12'h  0;
rom[111929] = 12'h  0;
rom[111930] = 12'h  0;
rom[111931] = 12'h  0;
rom[111932] = 12'h  0;
rom[111933] = 12'h  0;
rom[111934] = 12'h  0;
rom[111935] = 12'h  0;
rom[111936] = 12'h  0;
rom[111937] = 12'h  0;
rom[111938] = 12'h  0;
rom[111939] = 12'h  0;
rom[111940] = 12'h  0;
rom[111941] = 12'h  0;
rom[111942] = 12'h  0;
rom[111943] = 12'h  0;
rom[111944] = 12'h  0;
rom[111945] = 12'h  0;
rom[111946] = 12'h  0;
rom[111947] = 12'h  0;
rom[111948] = 12'h  0;
rom[111949] = 12'h  0;
rom[111950] = 12'h  0;
rom[111951] = 12'h  0;
rom[111952] = 12'h  0;
rom[111953] = 12'h  0;
rom[111954] = 12'h  0;
rom[111955] = 12'h111;
rom[111956] = 12'h111;
rom[111957] = 12'h  0;
rom[111958] = 12'h  0;
rom[111959] = 12'h111;
rom[111960] = 12'h111;
rom[111961] = 12'h111;
rom[111962] = 12'h333;
rom[111963] = 12'h666;
rom[111964] = 12'h999;
rom[111965] = 12'hccc;
rom[111966] = 12'hddd;
rom[111967] = 12'haaa;
rom[111968] = 12'h555;
rom[111969] = 12'h444;
rom[111970] = 12'h222;
rom[111971] = 12'h111;
rom[111972] = 12'h111;
rom[111973] = 12'h111;
rom[111974] = 12'h  0;
rom[111975] = 12'h  0;
rom[111976] = 12'h  0;
rom[111977] = 12'h  0;
rom[111978] = 12'h  0;
rom[111979] = 12'h  0;
rom[111980] = 12'h  0;
rom[111981] = 12'h  0;
rom[111982] = 12'h  0;
rom[111983] = 12'h  0;
rom[111984] = 12'h  0;
rom[111985] = 12'h  0;
rom[111986] = 12'h  0;
rom[111987] = 12'h  0;
rom[111988] = 12'h  0;
rom[111989] = 12'h  0;
rom[111990] = 12'h  0;
rom[111991] = 12'h  0;
rom[111992] = 12'h  0;
rom[111993] = 12'h  0;
rom[111994] = 12'h  0;
rom[111995] = 12'h  0;
rom[111996] = 12'h  0;
rom[111997] = 12'h  0;
rom[111998] = 12'h  0;
rom[111999] = 12'h  0;
rom[112000] = 12'hfff;
rom[112001] = 12'hfff;
rom[112002] = 12'hfff;
rom[112003] = 12'hfff;
rom[112004] = 12'hfff;
rom[112005] = 12'hfff;
rom[112006] = 12'hfff;
rom[112007] = 12'hfff;
rom[112008] = 12'hfff;
rom[112009] = 12'hfff;
rom[112010] = 12'hfff;
rom[112011] = 12'hfff;
rom[112012] = 12'hfff;
rom[112013] = 12'hfff;
rom[112014] = 12'hfff;
rom[112015] = 12'hfff;
rom[112016] = 12'hfff;
rom[112017] = 12'hfff;
rom[112018] = 12'hfff;
rom[112019] = 12'hfff;
rom[112020] = 12'hfff;
rom[112021] = 12'hfff;
rom[112022] = 12'hfff;
rom[112023] = 12'hfff;
rom[112024] = 12'hfff;
rom[112025] = 12'hfff;
rom[112026] = 12'hfff;
rom[112027] = 12'hfff;
rom[112028] = 12'hfff;
rom[112029] = 12'hfff;
rom[112030] = 12'hfff;
rom[112031] = 12'hfff;
rom[112032] = 12'hfff;
rom[112033] = 12'hfff;
rom[112034] = 12'hfff;
rom[112035] = 12'heee;
rom[112036] = 12'heee;
rom[112037] = 12'heee;
rom[112038] = 12'heee;
rom[112039] = 12'hfff;
rom[112040] = 12'hfff;
rom[112041] = 12'hfff;
rom[112042] = 12'heee;
rom[112043] = 12'heee;
rom[112044] = 12'heee;
rom[112045] = 12'heee;
rom[112046] = 12'heee;
rom[112047] = 12'heee;
rom[112048] = 12'heee;
rom[112049] = 12'heee;
rom[112050] = 12'heee;
rom[112051] = 12'heee;
rom[112052] = 12'hddd;
rom[112053] = 12'hddd;
rom[112054] = 12'hddd;
rom[112055] = 12'hddd;
rom[112056] = 12'hddd;
rom[112057] = 12'hddd;
rom[112058] = 12'hddd;
rom[112059] = 12'hccc;
rom[112060] = 12'hccc;
rom[112061] = 12'hccc;
rom[112062] = 12'hccc;
rom[112063] = 12'hccc;
rom[112064] = 12'hccc;
rom[112065] = 12'hccc;
rom[112066] = 12'hddd;
rom[112067] = 12'hddd;
rom[112068] = 12'hddd;
rom[112069] = 12'hccc;
rom[112070] = 12'hccc;
rom[112071] = 12'hbbb;
rom[112072] = 12'hccc;
rom[112073] = 12'hccc;
rom[112074] = 12'hccc;
rom[112075] = 12'hbbb;
rom[112076] = 12'hbbb;
rom[112077] = 12'hbbb;
rom[112078] = 12'hbbb;
rom[112079] = 12'hbbb;
rom[112080] = 12'hbbb;
rom[112081] = 12'haaa;
rom[112082] = 12'hbbb;
rom[112083] = 12'hccc;
rom[112084] = 12'heee;
rom[112085] = 12'heee;
rom[112086] = 12'heee;
rom[112087] = 12'hddd;
rom[112088] = 12'heee;
rom[112089] = 12'heee;
rom[112090] = 12'hddd;
rom[112091] = 12'hbbb;
rom[112092] = 12'haaa;
rom[112093] = 12'haaa;
rom[112094] = 12'haaa;
rom[112095] = 12'haaa;
rom[112096] = 12'h999;
rom[112097] = 12'h999;
rom[112098] = 12'h999;
rom[112099] = 12'h999;
rom[112100] = 12'h999;
rom[112101] = 12'h999;
rom[112102] = 12'haaa;
rom[112103] = 12'hbbb;
rom[112104] = 12'hccc;
rom[112105] = 12'hddd;
rom[112106] = 12'hddd;
rom[112107] = 12'hccc;
rom[112108] = 12'haaa;
rom[112109] = 12'h999;
rom[112110] = 12'h999;
rom[112111] = 12'h999;
rom[112112] = 12'h999;
rom[112113] = 12'h999;
rom[112114] = 12'h999;
rom[112115] = 12'h999;
rom[112116] = 12'h999;
rom[112117] = 12'h999;
rom[112118] = 12'h999;
rom[112119] = 12'h999;
rom[112120] = 12'h999;
rom[112121] = 12'h999;
rom[112122] = 12'h999;
rom[112123] = 12'h999;
rom[112124] = 12'haaa;
rom[112125] = 12'haaa;
rom[112126] = 12'h999;
rom[112127] = 12'h888;
rom[112128] = 12'h777;
rom[112129] = 12'h777;
rom[112130] = 12'h777;
rom[112131] = 12'h777;
rom[112132] = 12'h888;
rom[112133] = 12'h888;
rom[112134] = 12'h888;
rom[112135] = 12'h888;
rom[112136] = 12'h777;
rom[112137] = 12'h777;
rom[112138] = 12'h666;
rom[112139] = 12'h666;
rom[112140] = 12'h777;
rom[112141] = 12'h777;
rom[112142] = 12'h888;
rom[112143] = 12'h999;
rom[112144] = 12'h888;
rom[112145] = 12'h777;
rom[112146] = 12'h666;
rom[112147] = 12'h666;
rom[112148] = 12'h777;
rom[112149] = 12'h777;
rom[112150] = 12'h777;
rom[112151] = 12'h777;
rom[112152] = 12'h777;
rom[112153] = 12'h888;
rom[112154] = 12'h888;
rom[112155] = 12'h888;
rom[112156] = 12'h999;
rom[112157] = 12'h999;
rom[112158] = 12'haaa;
rom[112159] = 12'haaa;
rom[112160] = 12'haaa;
rom[112161] = 12'haaa;
rom[112162] = 12'hbbb;
rom[112163] = 12'hbbb;
rom[112164] = 12'hbbb;
rom[112165] = 12'hccc;
rom[112166] = 12'hddd;
rom[112167] = 12'hddd;
rom[112168] = 12'heee;
rom[112169] = 12'heee;
rom[112170] = 12'hfff;
rom[112171] = 12'hfff;
rom[112172] = 12'hfff;
rom[112173] = 12'hfff;
rom[112174] = 12'hfff;
rom[112175] = 12'hfff;
rom[112176] = 12'hfff;
rom[112177] = 12'hfff;
rom[112178] = 12'hfff;
rom[112179] = 12'hfff;
rom[112180] = 12'hfff;
rom[112181] = 12'hfff;
rom[112182] = 12'hfff;
rom[112183] = 12'hfff;
rom[112184] = 12'hfff;
rom[112185] = 12'hfff;
rom[112186] = 12'hfff;
rom[112187] = 12'hfff;
rom[112188] = 12'hfff;
rom[112189] = 12'hfff;
rom[112190] = 12'hfff;
rom[112191] = 12'hfff;
rom[112192] = 12'hfff;
rom[112193] = 12'hfff;
rom[112194] = 12'hfff;
rom[112195] = 12'hfff;
rom[112196] = 12'hfff;
rom[112197] = 12'hfff;
rom[112198] = 12'hfff;
rom[112199] = 12'hfff;
rom[112200] = 12'hfff;
rom[112201] = 12'hfff;
rom[112202] = 12'hfff;
rom[112203] = 12'hfff;
rom[112204] = 12'hfff;
rom[112205] = 12'hfff;
rom[112206] = 12'hfff;
rom[112207] = 12'hfff;
rom[112208] = 12'hfff;
rom[112209] = 12'hfff;
rom[112210] = 12'hfff;
rom[112211] = 12'hfff;
rom[112212] = 12'hfff;
rom[112213] = 12'hfff;
rom[112214] = 12'heee;
rom[112215] = 12'hddd;
rom[112216] = 12'hddd;
rom[112217] = 12'hddd;
rom[112218] = 12'hbbb;
rom[112219] = 12'hbbb;
rom[112220] = 12'hbbb;
rom[112221] = 12'hbbb;
rom[112222] = 12'h999;
rom[112223] = 12'h888;
rom[112224] = 12'h777;
rom[112225] = 12'h666;
rom[112226] = 12'h555;
rom[112227] = 12'h555;
rom[112228] = 12'h555;
rom[112229] = 12'h666;
rom[112230] = 12'h777;
rom[112231] = 12'h777;
rom[112232] = 12'h666;
rom[112233] = 12'h555;
rom[112234] = 12'h444;
rom[112235] = 12'h333;
rom[112236] = 12'h222;
rom[112237] = 12'h333;
rom[112238] = 12'h333;
rom[112239] = 12'h444;
rom[112240] = 12'h555;
rom[112241] = 12'h555;
rom[112242] = 12'h555;
rom[112243] = 12'h777;
rom[112244] = 12'hbbb;
rom[112245] = 12'hddd;
rom[112246] = 12'hccc;
rom[112247] = 12'h999;
rom[112248] = 12'h555;
rom[112249] = 12'h333;
rom[112250] = 12'h111;
rom[112251] = 12'h111;
rom[112252] = 12'h111;
rom[112253] = 12'h111;
rom[112254] = 12'h111;
rom[112255] = 12'h111;
rom[112256] = 12'h111;
rom[112257] = 12'h  0;
rom[112258] = 12'h222;
rom[112259] = 12'h333;
rom[112260] = 12'h333;
rom[112261] = 12'h222;
rom[112262] = 12'h333;
rom[112263] = 12'h888;
rom[112264] = 12'heee;
rom[112265] = 12'hfff;
rom[112266] = 12'hccc;
rom[112267] = 12'h666;
rom[112268] = 12'h444;
rom[112269] = 12'h333;
rom[112270] = 12'h222;
rom[112271] = 12'h222;
rom[112272] = 12'h333;
rom[112273] = 12'h888;
rom[112274] = 12'hccc;
rom[112275] = 12'hddd;
rom[112276] = 12'h666;
rom[112277] = 12'h222;
rom[112278] = 12'h111;
rom[112279] = 12'h111;
rom[112280] = 12'h  0;
rom[112281] = 12'h  0;
rom[112282] = 12'h  0;
rom[112283] = 12'h  0;
rom[112284] = 12'h  0;
rom[112285] = 12'h  0;
rom[112286] = 12'h111;
rom[112287] = 12'h555;
rom[112288] = 12'haaa;
rom[112289] = 12'hddd;
rom[112290] = 12'heee;
rom[112291] = 12'hbbb;
rom[112292] = 12'h444;
rom[112293] = 12'h111;
rom[112294] = 12'h111;
rom[112295] = 12'h222;
rom[112296] = 12'h222;
rom[112297] = 12'h111;
rom[112298] = 12'h111;
rom[112299] = 12'h111;
rom[112300] = 12'h222;
rom[112301] = 12'h111;
rom[112302] = 12'h111;
rom[112303] = 12'h111;
rom[112304] = 12'h222;
rom[112305] = 12'h222;
rom[112306] = 12'h444;
rom[112307] = 12'h888;
rom[112308] = 12'hbbb;
rom[112309] = 12'hccc;
rom[112310] = 12'hccc;
rom[112311] = 12'hccc;
rom[112312] = 12'hbbb;
rom[112313] = 12'h888;
rom[112314] = 12'h444;
rom[112315] = 12'h333;
rom[112316] = 12'h333;
rom[112317] = 12'h222;
rom[112318] = 12'h222;
rom[112319] = 12'h222;
rom[112320] = 12'h111;
rom[112321] = 12'h111;
rom[112322] = 12'h111;
rom[112323] = 12'h111;
rom[112324] = 12'h111;
rom[112325] = 12'h111;
rom[112326] = 12'h111;
rom[112327] = 12'h111;
rom[112328] = 12'h  0;
rom[112329] = 12'h  0;
rom[112330] = 12'h  0;
rom[112331] = 12'h  0;
rom[112332] = 12'h  0;
rom[112333] = 12'h  0;
rom[112334] = 12'h  0;
rom[112335] = 12'h  0;
rom[112336] = 12'h  0;
rom[112337] = 12'h  0;
rom[112338] = 12'h  0;
rom[112339] = 12'h  0;
rom[112340] = 12'h  0;
rom[112341] = 12'h  0;
rom[112342] = 12'h  0;
rom[112343] = 12'h  0;
rom[112344] = 12'h  0;
rom[112345] = 12'h  0;
rom[112346] = 12'h  0;
rom[112347] = 12'h  0;
rom[112348] = 12'h  0;
rom[112349] = 12'h  0;
rom[112350] = 12'h  0;
rom[112351] = 12'h  0;
rom[112352] = 12'h  0;
rom[112353] = 12'h  0;
rom[112354] = 12'h  0;
rom[112355] = 12'h  0;
rom[112356] = 12'h  0;
rom[112357] = 12'h  0;
rom[112358] = 12'h  0;
rom[112359] = 12'h  0;
rom[112360] = 12'h  0;
rom[112361] = 12'h111;
rom[112362] = 12'h111;
rom[112363] = 12'h333;
rom[112364] = 12'h666;
rom[112365] = 12'hbbb;
rom[112366] = 12'hddd;
rom[112367] = 12'hccc;
rom[112368] = 12'h888;
rom[112369] = 12'h555;
rom[112370] = 12'h222;
rom[112371] = 12'h222;
rom[112372] = 12'h222;
rom[112373] = 12'h111;
rom[112374] = 12'h  0;
rom[112375] = 12'h111;
rom[112376] = 12'h  0;
rom[112377] = 12'h  0;
rom[112378] = 12'h  0;
rom[112379] = 12'h  0;
rom[112380] = 12'h  0;
rom[112381] = 12'h  0;
rom[112382] = 12'h  0;
rom[112383] = 12'h  0;
rom[112384] = 12'h  0;
rom[112385] = 12'h  0;
rom[112386] = 12'h  0;
rom[112387] = 12'h  0;
rom[112388] = 12'h  0;
rom[112389] = 12'h  0;
rom[112390] = 12'h  0;
rom[112391] = 12'h  0;
rom[112392] = 12'h  0;
rom[112393] = 12'h  0;
rom[112394] = 12'h  0;
rom[112395] = 12'h  0;
rom[112396] = 12'h  0;
rom[112397] = 12'h  0;
rom[112398] = 12'h  0;
rom[112399] = 12'h  0;
rom[112400] = 12'hfff;
rom[112401] = 12'hfff;
rom[112402] = 12'hfff;
rom[112403] = 12'hfff;
rom[112404] = 12'hfff;
rom[112405] = 12'hfff;
rom[112406] = 12'hfff;
rom[112407] = 12'hfff;
rom[112408] = 12'hfff;
rom[112409] = 12'hfff;
rom[112410] = 12'hfff;
rom[112411] = 12'hfff;
rom[112412] = 12'hfff;
rom[112413] = 12'hfff;
rom[112414] = 12'hfff;
rom[112415] = 12'hfff;
rom[112416] = 12'hfff;
rom[112417] = 12'hfff;
rom[112418] = 12'hfff;
rom[112419] = 12'hfff;
rom[112420] = 12'hfff;
rom[112421] = 12'hfff;
rom[112422] = 12'hfff;
rom[112423] = 12'hfff;
rom[112424] = 12'hfff;
rom[112425] = 12'hfff;
rom[112426] = 12'hfff;
rom[112427] = 12'hfff;
rom[112428] = 12'hfff;
rom[112429] = 12'hfff;
rom[112430] = 12'hfff;
rom[112431] = 12'hfff;
rom[112432] = 12'hfff;
rom[112433] = 12'hfff;
rom[112434] = 12'hfff;
rom[112435] = 12'heee;
rom[112436] = 12'heee;
rom[112437] = 12'heee;
rom[112438] = 12'heee;
rom[112439] = 12'hfff;
rom[112440] = 12'hfff;
rom[112441] = 12'hfff;
rom[112442] = 12'heee;
rom[112443] = 12'heee;
rom[112444] = 12'heee;
rom[112445] = 12'heee;
rom[112446] = 12'heee;
rom[112447] = 12'heee;
rom[112448] = 12'heee;
rom[112449] = 12'heee;
rom[112450] = 12'heee;
rom[112451] = 12'heee;
rom[112452] = 12'hddd;
rom[112453] = 12'hddd;
rom[112454] = 12'hddd;
rom[112455] = 12'hddd;
rom[112456] = 12'hddd;
rom[112457] = 12'hddd;
rom[112458] = 12'hccc;
rom[112459] = 12'hccc;
rom[112460] = 12'hccc;
rom[112461] = 12'hccc;
rom[112462] = 12'hccc;
rom[112463] = 12'hccc;
rom[112464] = 12'hccc;
rom[112465] = 12'hccc;
rom[112466] = 12'hddd;
rom[112467] = 12'hddd;
rom[112468] = 12'hccc;
rom[112469] = 12'hccc;
rom[112470] = 12'hccc;
rom[112471] = 12'hccc;
rom[112472] = 12'hbbb;
rom[112473] = 12'hccc;
rom[112474] = 12'hccc;
rom[112475] = 12'hbbb;
rom[112476] = 12'hbbb;
rom[112477] = 12'hbbb;
rom[112478] = 12'hbbb;
rom[112479] = 12'hbbb;
rom[112480] = 12'hbbb;
rom[112481] = 12'hbbb;
rom[112482] = 12'hbbb;
rom[112483] = 12'hddd;
rom[112484] = 12'heee;
rom[112485] = 12'heee;
rom[112486] = 12'heee;
rom[112487] = 12'hfff;
rom[112488] = 12'heee;
rom[112489] = 12'hddd;
rom[112490] = 12'hccc;
rom[112491] = 12'hbbb;
rom[112492] = 12'haaa;
rom[112493] = 12'h999;
rom[112494] = 12'h999;
rom[112495] = 12'h999;
rom[112496] = 12'h999;
rom[112497] = 12'h999;
rom[112498] = 12'h999;
rom[112499] = 12'h999;
rom[112500] = 12'h999;
rom[112501] = 12'h999;
rom[112502] = 12'haaa;
rom[112503] = 12'hbbb;
rom[112504] = 12'hccc;
rom[112505] = 12'hddd;
rom[112506] = 12'hccc;
rom[112507] = 12'hbbb;
rom[112508] = 12'haaa;
rom[112509] = 12'h999;
rom[112510] = 12'h999;
rom[112511] = 12'h999;
rom[112512] = 12'h999;
rom[112513] = 12'h999;
rom[112514] = 12'h999;
rom[112515] = 12'h999;
rom[112516] = 12'h999;
rom[112517] = 12'h999;
rom[112518] = 12'h999;
rom[112519] = 12'h999;
rom[112520] = 12'h888;
rom[112521] = 12'h888;
rom[112522] = 12'h888;
rom[112523] = 12'h999;
rom[112524] = 12'h999;
rom[112525] = 12'h999;
rom[112526] = 12'h888;
rom[112527] = 12'h777;
rom[112528] = 12'h777;
rom[112529] = 12'h777;
rom[112530] = 12'h777;
rom[112531] = 12'h777;
rom[112532] = 12'h888;
rom[112533] = 12'h888;
rom[112534] = 12'h888;
rom[112535] = 12'h888;
rom[112536] = 12'h777;
rom[112537] = 12'h666;
rom[112538] = 12'h666;
rom[112539] = 12'h666;
rom[112540] = 12'h777;
rom[112541] = 12'h777;
rom[112542] = 12'h888;
rom[112543] = 12'h888;
rom[112544] = 12'h777;
rom[112545] = 12'h666;
rom[112546] = 12'h666;
rom[112547] = 12'h666;
rom[112548] = 12'h666;
rom[112549] = 12'h666;
rom[112550] = 12'h777;
rom[112551] = 12'h777;
rom[112552] = 12'h777;
rom[112553] = 12'h777;
rom[112554] = 12'h888;
rom[112555] = 12'h888;
rom[112556] = 12'h888;
rom[112557] = 12'h999;
rom[112558] = 12'h999;
rom[112559] = 12'h999;
rom[112560] = 12'h999;
rom[112561] = 12'haaa;
rom[112562] = 12'haaa;
rom[112563] = 12'haaa;
rom[112564] = 12'haaa;
rom[112565] = 12'hbbb;
rom[112566] = 12'hbbb;
rom[112567] = 12'hbbb;
rom[112568] = 12'hccc;
rom[112569] = 12'hddd;
rom[112570] = 12'hddd;
rom[112571] = 12'heee;
rom[112572] = 12'heee;
rom[112573] = 12'heee;
rom[112574] = 12'hfff;
rom[112575] = 12'hfff;
rom[112576] = 12'hfff;
rom[112577] = 12'hfff;
rom[112578] = 12'hfff;
rom[112579] = 12'hfff;
rom[112580] = 12'hfff;
rom[112581] = 12'hfff;
rom[112582] = 12'hfff;
rom[112583] = 12'hfff;
rom[112584] = 12'hfff;
rom[112585] = 12'hfff;
rom[112586] = 12'hfff;
rom[112587] = 12'hfff;
rom[112588] = 12'hfff;
rom[112589] = 12'hfff;
rom[112590] = 12'hfff;
rom[112591] = 12'hfff;
rom[112592] = 12'hfff;
rom[112593] = 12'hfff;
rom[112594] = 12'hfff;
rom[112595] = 12'hfff;
rom[112596] = 12'hfff;
rom[112597] = 12'hfff;
rom[112598] = 12'hfff;
rom[112599] = 12'hfff;
rom[112600] = 12'hfff;
rom[112601] = 12'hfff;
rom[112602] = 12'hfff;
rom[112603] = 12'hfff;
rom[112604] = 12'hfff;
rom[112605] = 12'hfff;
rom[112606] = 12'hfff;
rom[112607] = 12'hfff;
rom[112608] = 12'hfff;
rom[112609] = 12'hfff;
rom[112610] = 12'hfff;
rom[112611] = 12'heee;
rom[112612] = 12'heee;
rom[112613] = 12'heee;
rom[112614] = 12'hddd;
rom[112615] = 12'hbbb;
rom[112616] = 12'hbbb;
rom[112617] = 12'haaa;
rom[112618] = 12'h999;
rom[112619] = 12'h999;
rom[112620] = 12'haaa;
rom[112621] = 12'hbbb;
rom[112622] = 12'haaa;
rom[112623] = 12'h888;
rom[112624] = 12'h666;
rom[112625] = 12'h555;
rom[112626] = 12'h555;
rom[112627] = 12'h444;
rom[112628] = 12'h555;
rom[112629] = 12'h555;
rom[112630] = 12'h666;
rom[112631] = 12'h777;
rom[112632] = 12'h666;
rom[112633] = 12'h555;
rom[112634] = 12'h444;
rom[112635] = 12'h333;
rom[112636] = 12'h222;
rom[112637] = 12'h222;
rom[112638] = 12'h333;
rom[112639] = 12'h444;
rom[112640] = 12'h444;
rom[112641] = 12'h444;
rom[112642] = 12'h555;
rom[112643] = 12'h888;
rom[112644] = 12'hccc;
rom[112645] = 12'heee;
rom[112646] = 12'hbbb;
rom[112647] = 12'h777;
rom[112648] = 12'h444;
rom[112649] = 12'h222;
rom[112650] = 12'h111;
rom[112651] = 12'h111;
rom[112652] = 12'h111;
rom[112653] = 12'h111;
rom[112654] = 12'h  0;
rom[112655] = 12'h111;
rom[112656] = 12'h  0;
rom[112657] = 12'h  0;
rom[112658] = 12'h222;
rom[112659] = 12'h333;
rom[112660] = 12'h333;
rom[112661] = 12'h222;
rom[112662] = 12'h333;
rom[112663] = 12'h777;
rom[112664] = 12'heee;
rom[112665] = 12'hfff;
rom[112666] = 12'hccc;
rom[112667] = 12'h666;
rom[112668] = 12'h444;
rom[112669] = 12'h333;
rom[112670] = 12'h222;
rom[112671] = 12'h222;
rom[112672] = 12'h222;
rom[112673] = 12'h666;
rom[112674] = 12'hbbb;
rom[112675] = 12'hddd;
rom[112676] = 12'h777;
rom[112677] = 12'h333;
rom[112678] = 12'h  0;
rom[112679] = 12'h111;
rom[112680] = 12'h  0;
rom[112681] = 12'h  0;
rom[112682] = 12'h  0;
rom[112683] = 12'h  0;
rom[112684] = 12'h  0;
rom[112685] = 12'h  0;
rom[112686] = 12'h111;
rom[112687] = 12'h333;
rom[112688] = 12'h888;
rom[112689] = 12'haaa;
rom[112690] = 12'hddd;
rom[112691] = 12'hddd;
rom[112692] = 12'h777;
rom[112693] = 12'h222;
rom[112694] = 12'h111;
rom[112695] = 12'h111;
rom[112696] = 12'h111;
rom[112697] = 12'h111;
rom[112698] = 12'h111;
rom[112699] = 12'h111;
rom[112700] = 12'h111;
rom[112701] = 12'h111;
rom[112702] = 12'h111;
rom[112703] = 12'h222;
rom[112704] = 12'h111;
rom[112705] = 12'h222;
rom[112706] = 12'h333;
rom[112707] = 12'h666;
rom[112708] = 12'h999;
rom[112709] = 12'haaa;
rom[112710] = 12'hccc;
rom[112711] = 12'hccc;
rom[112712] = 12'hccc;
rom[112713] = 12'h999;
rom[112714] = 12'h666;
rom[112715] = 12'h444;
rom[112716] = 12'h333;
rom[112717] = 12'h222;
rom[112718] = 12'h222;
rom[112719] = 12'h222;
rom[112720] = 12'h111;
rom[112721] = 12'h111;
rom[112722] = 12'h111;
rom[112723] = 12'h111;
rom[112724] = 12'h111;
rom[112725] = 12'h111;
rom[112726] = 12'h111;
rom[112727] = 12'h111;
rom[112728] = 12'h  0;
rom[112729] = 12'h  0;
rom[112730] = 12'h  0;
rom[112731] = 12'h  0;
rom[112732] = 12'h  0;
rom[112733] = 12'h  0;
rom[112734] = 12'h  0;
rom[112735] = 12'h  0;
rom[112736] = 12'h  0;
rom[112737] = 12'h  0;
rom[112738] = 12'h  0;
rom[112739] = 12'h  0;
rom[112740] = 12'h  0;
rom[112741] = 12'h  0;
rom[112742] = 12'h  0;
rom[112743] = 12'h  0;
rom[112744] = 12'h  0;
rom[112745] = 12'h  0;
rom[112746] = 12'h  0;
rom[112747] = 12'h  0;
rom[112748] = 12'h  0;
rom[112749] = 12'h  0;
rom[112750] = 12'h  0;
rom[112751] = 12'h  0;
rom[112752] = 12'h  0;
rom[112753] = 12'h  0;
rom[112754] = 12'h  0;
rom[112755] = 12'h  0;
rom[112756] = 12'h  0;
rom[112757] = 12'h  0;
rom[112758] = 12'h  0;
rom[112759] = 12'h  0;
rom[112760] = 12'h  0;
rom[112761] = 12'h111;
rom[112762] = 12'h111;
rom[112763] = 12'h222;
rom[112764] = 12'h444;
rom[112765] = 12'h888;
rom[112766] = 12'hbbb;
rom[112767] = 12'hccc;
rom[112768] = 12'h999;
rom[112769] = 12'h666;
rom[112770] = 12'h444;
rom[112771] = 12'h222;
rom[112772] = 12'h222;
rom[112773] = 12'h111;
rom[112774] = 12'h  0;
rom[112775] = 12'h  0;
rom[112776] = 12'h  0;
rom[112777] = 12'h  0;
rom[112778] = 12'h  0;
rom[112779] = 12'h  0;
rom[112780] = 12'h  0;
rom[112781] = 12'h  0;
rom[112782] = 12'h  0;
rom[112783] = 12'h  0;
rom[112784] = 12'h  0;
rom[112785] = 12'h  0;
rom[112786] = 12'h  0;
rom[112787] = 12'h  0;
rom[112788] = 12'h  0;
rom[112789] = 12'h  0;
rom[112790] = 12'h  0;
rom[112791] = 12'h  0;
rom[112792] = 12'h  0;
rom[112793] = 12'h  0;
rom[112794] = 12'h  0;
rom[112795] = 12'h  0;
rom[112796] = 12'h  0;
rom[112797] = 12'h  0;
rom[112798] = 12'h  0;
rom[112799] = 12'h  0;
rom[112800] = 12'hfff;
rom[112801] = 12'hfff;
rom[112802] = 12'hfff;
rom[112803] = 12'hfff;
rom[112804] = 12'hfff;
rom[112805] = 12'hfff;
rom[112806] = 12'hfff;
rom[112807] = 12'hfff;
rom[112808] = 12'hfff;
rom[112809] = 12'hfff;
rom[112810] = 12'hfff;
rom[112811] = 12'hfff;
rom[112812] = 12'hfff;
rom[112813] = 12'hfff;
rom[112814] = 12'hfff;
rom[112815] = 12'hfff;
rom[112816] = 12'hfff;
rom[112817] = 12'hfff;
rom[112818] = 12'hfff;
rom[112819] = 12'hfff;
rom[112820] = 12'hfff;
rom[112821] = 12'hfff;
rom[112822] = 12'hfff;
rom[112823] = 12'hfff;
rom[112824] = 12'hfff;
rom[112825] = 12'hfff;
rom[112826] = 12'hfff;
rom[112827] = 12'hfff;
rom[112828] = 12'hfff;
rom[112829] = 12'hfff;
rom[112830] = 12'hfff;
rom[112831] = 12'hfff;
rom[112832] = 12'hfff;
rom[112833] = 12'hfff;
rom[112834] = 12'hfff;
rom[112835] = 12'heee;
rom[112836] = 12'heee;
rom[112837] = 12'heee;
rom[112838] = 12'heee;
rom[112839] = 12'hfff;
rom[112840] = 12'heee;
rom[112841] = 12'heee;
rom[112842] = 12'heee;
rom[112843] = 12'heee;
rom[112844] = 12'heee;
rom[112845] = 12'heee;
rom[112846] = 12'heee;
rom[112847] = 12'heee;
rom[112848] = 12'heee;
rom[112849] = 12'heee;
rom[112850] = 12'heee;
rom[112851] = 12'hddd;
rom[112852] = 12'hddd;
rom[112853] = 12'hddd;
rom[112854] = 12'hddd;
rom[112855] = 12'hddd;
rom[112856] = 12'hddd;
rom[112857] = 12'hddd;
rom[112858] = 12'hccc;
rom[112859] = 12'hccc;
rom[112860] = 12'hccc;
rom[112861] = 12'hccc;
rom[112862] = 12'hccc;
rom[112863] = 12'hccc;
rom[112864] = 12'hccc;
rom[112865] = 12'hccc;
rom[112866] = 12'hddd;
rom[112867] = 12'hddd;
rom[112868] = 12'hccc;
rom[112869] = 12'hccc;
rom[112870] = 12'hccc;
rom[112871] = 12'hccc;
rom[112872] = 12'hbbb;
rom[112873] = 12'hccc;
rom[112874] = 12'hbbb;
rom[112875] = 12'hbbb;
rom[112876] = 12'hbbb;
rom[112877] = 12'hbbb;
rom[112878] = 12'hbbb;
rom[112879] = 12'haaa;
rom[112880] = 12'hbbb;
rom[112881] = 12'hbbb;
rom[112882] = 12'hccc;
rom[112883] = 12'heee;
rom[112884] = 12'heee;
rom[112885] = 12'heee;
rom[112886] = 12'heee;
rom[112887] = 12'hfff;
rom[112888] = 12'hddd;
rom[112889] = 12'hbbb;
rom[112890] = 12'haaa;
rom[112891] = 12'haaa;
rom[112892] = 12'haaa;
rom[112893] = 12'h999;
rom[112894] = 12'h999;
rom[112895] = 12'h999;
rom[112896] = 12'h999;
rom[112897] = 12'h999;
rom[112898] = 12'h999;
rom[112899] = 12'h999;
rom[112900] = 12'h999;
rom[112901] = 12'haaa;
rom[112902] = 12'hbbb;
rom[112903] = 12'hbbb;
rom[112904] = 12'hccc;
rom[112905] = 12'hccc;
rom[112906] = 12'hccc;
rom[112907] = 12'haaa;
rom[112908] = 12'h999;
rom[112909] = 12'h999;
rom[112910] = 12'h999;
rom[112911] = 12'h999;
rom[112912] = 12'h999;
rom[112913] = 12'h999;
rom[112914] = 12'h999;
rom[112915] = 12'h999;
rom[112916] = 12'h999;
rom[112917] = 12'h999;
rom[112918] = 12'h888;
rom[112919] = 12'h888;
rom[112920] = 12'h888;
rom[112921] = 12'h888;
rom[112922] = 12'h888;
rom[112923] = 12'h888;
rom[112924] = 12'h999;
rom[112925] = 12'h999;
rom[112926] = 12'h777;
rom[112927] = 12'h666;
rom[112928] = 12'h666;
rom[112929] = 12'h666;
rom[112930] = 12'h777;
rom[112931] = 12'h777;
rom[112932] = 12'h888;
rom[112933] = 12'h888;
rom[112934] = 12'h777;
rom[112935] = 12'h777;
rom[112936] = 12'h666;
rom[112937] = 12'h666;
rom[112938] = 12'h666;
rom[112939] = 12'h666;
rom[112940] = 12'h777;
rom[112941] = 12'h888;
rom[112942] = 12'h888;
rom[112943] = 12'h777;
rom[112944] = 12'h666;
rom[112945] = 12'h666;
rom[112946] = 12'h666;
rom[112947] = 12'h666;
rom[112948] = 12'h666;
rom[112949] = 12'h666;
rom[112950] = 12'h666;
rom[112951] = 12'h777;
rom[112952] = 12'h777;
rom[112953] = 12'h777;
rom[112954] = 12'h777;
rom[112955] = 12'h777;
rom[112956] = 12'h888;
rom[112957] = 12'h888;
rom[112958] = 12'h888;
rom[112959] = 12'h999;
rom[112960] = 12'h999;
rom[112961] = 12'h999;
rom[112962] = 12'h999;
rom[112963] = 12'haaa;
rom[112964] = 12'haaa;
rom[112965] = 12'haaa;
rom[112966] = 12'haaa;
rom[112967] = 12'haaa;
rom[112968] = 12'hbbb;
rom[112969] = 12'hbbb;
rom[112970] = 12'hccc;
rom[112971] = 12'hccc;
rom[112972] = 12'hddd;
rom[112973] = 12'hddd;
rom[112974] = 12'hddd;
rom[112975] = 12'heee;
rom[112976] = 12'heee;
rom[112977] = 12'heee;
rom[112978] = 12'hfff;
rom[112979] = 12'hfff;
rom[112980] = 12'hfff;
rom[112981] = 12'hfff;
rom[112982] = 12'hfff;
rom[112983] = 12'hfff;
rom[112984] = 12'hfff;
rom[112985] = 12'hfff;
rom[112986] = 12'hfff;
rom[112987] = 12'hfff;
rom[112988] = 12'hfff;
rom[112989] = 12'hfff;
rom[112990] = 12'hfff;
rom[112991] = 12'hfff;
rom[112992] = 12'hfff;
rom[112993] = 12'hfff;
rom[112994] = 12'hfff;
rom[112995] = 12'hfff;
rom[112996] = 12'hfff;
rom[112997] = 12'hfff;
rom[112998] = 12'hfff;
rom[112999] = 12'hfff;
rom[113000] = 12'hfff;
rom[113001] = 12'hfff;
rom[113002] = 12'hfff;
rom[113003] = 12'hfff;
rom[113004] = 12'hfff;
rom[113005] = 12'hfff;
rom[113006] = 12'hfff;
rom[113007] = 12'hfff;
rom[113008] = 12'hfff;
rom[113009] = 12'heee;
rom[113010] = 12'hddd;
rom[113011] = 12'hddd;
rom[113012] = 12'hccc;
rom[113013] = 12'hccc;
rom[113014] = 12'hbbb;
rom[113015] = 12'haaa;
rom[113016] = 12'h999;
rom[113017] = 12'h888;
rom[113018] = 12'h888;
rom[113019] = 12'h888;
rom[113020] = 12'haaa;
rom[113021] = 12'hbbb;
rom[113022] = 12'hbbb;
rom[113023] = 12'h999;
rom[113024] = 12'h666;
rom[113025] = 12'h555;
rom[113026] = 12'h444;
rom[113027] = 12'h444;
rom[113028] = 12'h444;
rom[113029] = 12'h444;
rom[113030] = 12'h555;
rom[113031] = 12'h666;
rom[113032] = 12'h666;
rom[113033] = 12'h555;
rom[113034] = 12'h444;
rom[113035] = 12'h333;
rom[113036] = 12'h222;
rom[113037] = 12'h222;
rom[113038] = 12'h333;
rom[113039] = 12'h333;
rom[113040] = 12'h444;
rom[113041] = 12'h444;
rom[113042] = 12'h555;
rom[113043] = 12'h999;
rom[113044] = 12'hddd;
rom[113045] = 12'hddd;
rom[113046] = 12'h999;
rom[113047] = 12'h555;
rom[113048] = 12'h222;
rom[113049] = 12'h111;
rom[113050] = 12'h111;
rom[113051] = 12'h111;
rom[113052] = 12'h111;
rom[113053] = 12'h  0;
rom[113054] = 12'h  0;
rom[113055] = 12'h  0;
rom[113056] = 12'h111;
rom[113057] = 12'h  0;
rom[113058] = 12'h111;
rom[113059] = 12'h222;
rom[113060] = 12'h222;
rom[113061] = 12'h222;
rom[113062] = 12'h222;
rom[113063] = 12'h777;
rom[113064] = 12'heee;
rom[113065] = 12'hfff;
rom[113066] = 12'hccc;
rom[113067] = 12'h666;
rom[113068] = 12'h444;
rom[113069] = 12'h333;
rom[113070] = 12'h222;
rom[113071] = 12'h111;
rom[113072] = 12'h111;
rom[113073] = 12'h555;
rom[113074] = 12'haaa;
rom[113075] = 12'heee;
rom[113076] = 12'h999;
rom[113077] = 12'h333;
rom[113078] = 12'h  0;
rom[113079] = 12'h  0;
rom[113080] = 12'h  0;
rom[113081] = 12'h111;
rom[113082] = 12'h  0;
rom[113083] = 12'h111;
rom[113084] = 12'h111;
rom[113085] = 12'h  0;
rom[113086] = 12'h  0;
rom[113087] = 12'h222;
rom[113088] = 12'h777;
rom[113089] = 12'h888;
rom[113090] = 12'hccc;
rom[113091] = 12'heee;
rom[113092] = 12'haaa;
rom[113093] = 12'h444;
rom[113094] = 12'h222;
rom[113095] = 12'h111;
rom[113096] = 12'h  0;
rom[113097] = 12'h111;
rom[113098] = 12'h111;
rom[113099] = 12'h111;
rom[113100] = 12'h111;
rom[113101] = 12'h111;
rom[113102] = 12'h222;
rom[113103] = 12'h222;
rom[113104] = 12'h111;
rom[113105] = 12'h111;
rom[113106] = 12'h222;
rom[113107] = 12'h444;
rom[113108] = 12'h666;
rom[113109] = 12'h888;
rom[113110] = 12'haaa;
rom[113111] = 12'hccc;
rom[113112] = 12'hccc;
rom[113113] = 12'hbbb;
rom[113114] = 12'h888;
rom[113115] = 12'h555;
rom[113116] = 12'h333;
rom[113117] = 12'h222;
rom[113118] = 12'h222;
rom[113119] = 12'h222;
rom[113120] = 12'h111;
rom[113121] = 12'h111;
rom[113122] = 12'h222;
rom[113123] = 12'h222;
rom[113124] = 12'h111;
rom[113125] = 12'h111;
rom[113126] = 12'h  0;
rom[113127] = 12'h  0;
rom[113128] = 12'h  0;
rom[113129] = 12'h  0;
rom[113130] = 12'h  0;
rom[113131] = 12'h  0;
rom[113132] = 12'h  0;
rom[113133] = 12'h  0;
rom[113134] = 12'h  0;
rom[113135] = 12'h  0;
rom[113136] = 12'h  0;
rom[113137] = 12'h  0;
rom[113138] = 12'h  0;
rom[113139] = 12'h  0;
rom[113140] = 12'h  0;
rom[113141] = 12'h  0;
rom[113142] = 12'h  0;
rom[113143] = 12'h  0;
rom[113144] = 12'h  0;
rom[113145] = 12'h  0;
rom[113146] = 12'h  0;
rom[113147] = 12'h  0;
rom[113148] = 12'h  0;
rom[113149] = 12'h  0;
rom[113150] = 12'h  0;
rom[113151] = 12'h  0;
rom[113152] = 12'h  0;
rom[113153] = 12'h  0;
rom[113154] = 12'h  0;
rom[113155] = 12'h  0;
rom[113156] = 12'h  0;
rom[113157] = 12'h  0;
rom[113158] = 12'h  0;
rom[113159] = 12'h  0;
rom[113160] = 12'h  0;
rom[113161] = 12'h111;
rom[113162] = 12'h111;
rom[113163] = 12'h111;
rom[113164] = 12'h222;
rom[113165] = 12'h555;
rom[113166] = 12'h888;
rom[113167] = 12'hbbb;
rom[113168] = 12'hbbb;
rom[113169] = 12'h999;
rom[113170] = 12'h555;
rom[113171] = 12'h333;
rom[113172] = 12'h222;
rom[113173] = 12'h111;
rom[113174] = 12'h111;
rom[113175] = 12'h  0;
rom[113176] = 12'h  0;
rom[113177] = 12'h  0;
rom[113178] = 12'h  0;
rom[113179] = 12'h  0;
rom[113180] = 12'h  0;
rom[113181] = 12'h  0;
rom[113182] = 12'h  0;
rom[113183] = 12'h  0;
rom[113184] = 12'h  0;
rom[113185] = 12'h  0;
rom[113186] = 12'h  0;
rom[113187] = 12'h  0;
rom[113188] = 12'h  0;
rom[113189] = 12'h  0;
rom[113190] = 12'h  0;
rom[113191] = 12'h  0;
rom[113192] = 12'h  0;
rom[113193] = 12'h  0;
rom[113194] = 12'h  0;
rom[113195] = 12'h  0;
rom[113196] = 12'h  0;
rom[113197] = 12'h  0;
rom[113198] = 12'h  0;
rom[113199] = 12'h  0;
rom[113200] = 12'hfff;
rom[113201] = 12'hfff;
rom[113202] = 12'hfff;
rom[113203] = 12'hfff;
rom[113204] = 12'hfff;
rom[113205] = 12'hfff;
rom[113206] = 12'hfff;
rom[113207] = 12'hfff;
rom[113208] = 12'hfff;
rom[113209] = 12'hfff;
rom[113210] = 12'hfff;
rom[113211] = 12'hfff;
rom[113212] = 12'hfff;
rom[113213] = 12'hfff;
rom[113214] = 12'hfff;
rom[113215] = 12'hfff;
rom[113216] = 12'hfff;
rom[113217] = 12'hfff;
rom[113218] = 12'hfff;
rom[113219] = 12'hfff;
rom[113220] = 12'hfff;
rom[113221] = 12'hfff;
rom[113222] = 12'hfff;
rom[113223] = 12'hfff;
rom[113224] = 12'hfff;
rom[113225] = 12'hfff;
rom[113226] = 12'hfff;
rom[113227] = 12'hfff;
rom[113228] = 12'hfff;
rom[113229] = 12'hfff;
rom[113230] = 12'hfff;
rom[113231] = 12'hfff;
rom[113232] = 12'hfff;
rom[113233] = 12'hfff;
rom[113234] = 12'hfff;
rom[113235] = 12'heee;
rom[113236] = 12'heee;
rom[113237] = 12'heee;
rom[113238] = 12'heee;
rom[113239] = 12'heee;
rom[113240] = 12'heee;
rom[113241] = 12'heee;
rom[113242] = 12'heee;
rom[113243] = 12'heee;
rom[113244] = 12'heee;
rom[113245] = 12'heee;
rom[113246] = 12'heee;
rom[113247] = 12'heee;
rom[113248] = 12'heee;
rom[113249] = 12'hddd;
rom[113250] = 12'hddd;
rom[113251] = 12'hddd;
rom[113252] = 12'hddd;
rom[113253] = 12'hddd;
rom[113254] = 12'hddd;
rom[113255] = 12'hddd;
rom[113256] = 12'hccc;
rom[113257] = 12'hccc;
rom[113258] = 12'hccc;
rom[113259] = 12'hccc;
rom[113260] = 12'hccc;
rom[113261] = 12'hccc;
rom[113262] = 12'hccc;
rom[113263] = 12'hccc;
rom[113264] = 12'hccc;
rom[113265] = 12'hccc;
rom[113266] = 12'hddd;
rom[113267] = 12'hccc;
rom[113268] = 12'hccc;
rom[113269] = 12'hbbb;
rom[113270] = 12'hbbb;
rom[113271] = 12'hccc;
rom[113272] = 12'hccc;
rom[113273] = 12'hbbb;
rom[113274] = 12'hbbb;
rom[113275] = 12'hbbb;
rom[113276] = 12'hbbb;
rom[113277] = 12'hbbb;
rom[113278] = 12'hbbb;
rom[113279] = 12'haaa;
rom[113280] = 12'hbbb;
rom[113281] = 12'hccc;
rom[113282] = 12'hddd;
rom[113283] = 12'heee;
rom[113284] = 12'heee;
rom[113285] = 12'heee;
rom[113286] = 12'heee;
rom[113287] = 12'heee;
rom[113288] = 12'hccc;
rom[113289] = 12'haaa;
rom[113290] = 12'h999;
rom[113291] = 12'h999;
rom[113292] = 12'haaa;
rom[113293] = 12'haaa;
rom[113294] = 12'h999;
rom[113295] = 12'h999;
rom[113296] = 12'h999;
rom[113297] = 12'h999;
rom[113298] = 12'h999;
rom[113299] = 12'h999;
rom[113300] = 12'haaa;
rom[113301] = 12'hbbb;
rom[113302] = 12'hbbb;
rom[113303] = 12'hccc;
rom[113304] = 12'hccc;
rom[113305] = 12'hccc;
rom[113306] = 12'hbbb;
rom[113307] = 12'haaa;
rom[113308] = 12'h999;
rom[113309] = 12'h999;
rom[113310] = 12'h999;
rom[113311] = 12'h999;
rom[113312] = 12'h999;
rom[113313] = 12'h999;
rom[113314] = 12'h999;
rom[113315] = 12'h999;
rom[113316] = 12'h888;
rom[113317] = 12'h888;
rom[113318] = 12'h888;
rom[113319] = 12'h888;
rom[113320] = 12'h888;
rom[113321] = 12'h777;
rom[113322] = 12'h888;
rom[113323] = 12'h888;
rom[113324] = 12'h999;
rom[113325] = 12'h888;
rom[113326] = 12'h777;
rom[113327] = 12'h666;
rom[113328] = 12'h666;
rom[113329] = 12'h666;
rom[113330] = 12'h777;
rom[113331] = 12'h777;
rom[113332] = 12'h888;
rom[113333] = 12'h777;
rom[113334] = 12'h777;
rom[113335] = 12'h777;
rom[113336] = 12'h666;
rom[113337] = 12'h666;
rom[113338] = 12'h666;
rom[113339] = 12'h666;
rom[113340] = 12'h777;
rom[113341] = 12'h888;
rom[113342] = 12'h777;
rom[113343] = 12'h666;
rom[113344] = 12'h555;
rom[113345] = 12'h555;
rom[113346] = 12'h555;
rom[113347] = 12'h666;
rom[113348] = 12'h666;
rom[113349] = 12'h666;
rom[113350] = 12'h666;
rom[113351] = 12'h666;
rom[113352] = 12'h777;
rom[113353] = 12'h777;
rom[113354] = 12'h777;
rom[113355] = 12'h777;
rom[113356] = 12'h777;
rom[113357] = 12'h777;
rom[113358] = 12'h888;
rom[113359] = 12'h888;
rom[113360] = 12'h888;
rom[113361] = 12'h999;
rom[113362] = 12'h999;
rom[113363] = 12'h999;
rom[113364] = 12'haaa;
rom[113365] = 12'haaa;
rom[113366] = 12'haaa;
rom[113367] = 12'haaa;
rom[113368] = 12'haaa;
rom[113369] = 12'haaa;
rom[113370] = 12'hbbb;
rom[113371] = 12'hbbb;
rom[113372] = 12'hbbb;
rom[113373] = 12'hccc;
rom[113374] = 12'hccc;
rom[113375] = 12'hccc;
rom[113376] = 12'hddd;
rom[113377] = 12'hddd;
rom[113378] = 12'hddd;
rom[113379] = 12'heee;
rom[113380] = 12'heee;
rom[113381] = 12'heee;
rom[113382] = 12'hfff;
rom[113383] = 12'hfff;
rom[113384] = 12'hfff;
rom[113385] = 12'hfff;
rom[113386] = 12'hfff;
rom[113387] = 12'hfff;
rom[113388] = 12'hfff;
rom[113389] = 12'hfff;
rom[113390] = 12'hfff;
rom[113391] = 12'hfff;
rom[113392] = 12'hfff;
rom[113393] = 12'hfff;
rom[113394] = 12'hfff;
rom[113395] = 12'hfff;
rom[113396] = 12'hfff;
rom[113397] = 12'hfff;
rom[113398] = 12'hfff;
rom[113399] = 12'hfff;
rom[113400] = 12'hfff;
rom[113401] = 12'hfff;
rom[113402] = 12'hfff;
rom[113403] = 12'hfff;
rom[113404] = 12'hfff;
rom[113405] = 12'heee;
rom[113406] = 12'heee;
rom[113407] = 12'hddd;
rom[113408] = 12'hddd;
rom[113409] = 12'hccc;
rom[113410] = 12'hbbb;
rom[113411] = 12'hbbb;
rom[113412] = 12'haaa;
rom[113413] = 12'haaa;
rom[113414] = 12'h999;
rom[113415] = 12'h999;
rom[113416] = 12'h888;
rom[113417] = 12'h888;
rom[113418] = 12'h777;
rom[113419] = 12'h666;
rom[113420] = 12'h888;
rom[113421] = 12'haaa;
rom[113422] = 12'hbbb;
rom[113423] = 12'haaa;
rom[113424] = 12'h666;
rom[113425] = 12'h555;
rom[113426] = 12'h444;
rom[113427] = 12'h333;
rom[113428] = 12'h333;
rom[113429] = 12'h333;
rom[113430] = 12'h444;
rom[113431] = 12'h555;
rom[113432] = 12'h555;
rom[113433] = 12'h444;
rom[113434] = 12'h444;
rom[113435] = 12'h333;
rom[113436] = 12'h222;
rom[113437] = 12'h222;
rom[113438] = 12'h333;
rom[113439] = 12'h333;
rom[113440] = 12'h333;
rom[113441] = 12'h333;
rom[113442] = 12'h666;
rom[113443] = 12'haaa;
rom[113444] = 12'hddd;
rom[113445] = 12'hccc;
rom[113446] = 12'h777;
rom[113447] = 12'h333;
rom[113448] = 12'h222;
rom[113449] = 12'h111;
rom[113450] = 12'h111;
rom[113451] = 12'h111;
rom[113452] = 12'h111;
rom[113453] = 12'h  0;
rom[113454] = 12'h  0;
rom[113455] = 12'h111;
rom[113456] = 12'h111;
rom[113457] = 12'h  0;
rom[113458] = 12'h111;
rom[113459] = 12'h222;
rom[113460] = 12'h222;
rom[113461] = 12'h222;
rom[113462] = 12'h222;
rom[113463] = 12'h666;
rom[113464] = 12'hddd;
rom[113465] = 12'hfff;
rom[113466] = 12'hccc;
rom[113467] = 12'h666;
rom[113468] = 12'h333;
rom[113469] = 12'h333;
rom[113470] = 12'h222;
rom[113471] = 12'h111;
rom[113472] = 12'h111;
rom[113473] = 12'h333;
rom[113474] = 12'h999;
rom[113475] = 12'heee;
rom[113476] = 12'hbbb;
rom[113477] = 12'h555;
rom[113478] = 12'h  0;
rom[113479] = 12'h  0;
rom[113480] = 12'h111;
rom[113481] = 12'h111;
rom[113482] = 12'h  0;
rom[113483] = 12'h  0;
rom[113484] = 12'h111;
rom[113485] = 12'h  0;
rom[113486] = 12'h  0;
rom[113487] = 12'h111;
rom[113488] = 12'h666;
rom[113489] = 12'h888;
rom[113490] = 12'hbbb;
rom[113491] = 12'hccc;
rom[113492] = 12'hccc;
rom[113493] = 12'h777;
rom[113494] = 12'h222;
rom[113495] = 12'h111;
rom[113496] = 12'h  0;
rom[113497] = 12'h111;
rom[113498] = 12'h111;
rom[113499] = 12'h111;
rom[113500] = 12'h111;
rom[113501] = 12'h222;
rom[113502] = 12'h222;
rom[113503] = 12'h111;
rom[113504] = 12'h111;
rom[113505] = 12'h222;
rom[113506] = 12'h222;
rom[113507] = 12'h222;
rom[113508] = 12'h444;
rom[113509] = 12'h666;
rom[113510] = 12'h999;
rom[113511] = 12'haaa;
rom[113512] = 12'hccc;
rom[113513] = 12'hccc;
rom[113514] = 12'haaa;
rom[113515] = 12'h777;
rom[113516] = 12'h333;
rom[113517] = 12'h222;
rom[113518] = 12'h222;
rom[113519] = 12'h222;
rom[113520] = 12'h111;
rom[113521] = 12'h222;
rom[113522] = 12'h222;
rom[113523] = 12'h222;
rom[113524] = 12'h111;
rom[113525] = 12'h111;
rom[113526] = 12'h  0;
rom[113527] = 12'h  0;
rom[113528] = 12'h  0;
rom[113529] = 12'h  0;
rom[113530] = 12'h  0;
rom[113531] = 12'h  0;
rom[113532] = 12'h  0;
rom[113533] = 12'h  0;
rom[113534] = 12'h  0;
rom[113535] = 12'h  0;
rom[113536] = 12'h  0;
rom[113537] = 12'h  0;
rom[113538] = 12'h  0;
rom[113539] = 12'h  0;
rom[113540] = 12'h  0;
rom[113541] = 12'h  0;
rom[113542] = 12'h  0;
rom[113543] = 12'h  0;
rom[113544] = 12'h  0;
rom[113545] = 12'h  0;
rom[113546] = 12'h  0;
rom[113547] = 12'h  0;
rom[113548] = 12'h  0;
rom[113549] = 12'h  0;
rom[113550] = 12'h  0;
rom[113551] = 12'h  0;
rom[113552] = 12'h  0;
rom[113553] = 12'h  0;
rom[113554] = 12'h  0;
rom[113555] = 12'h  0;
rom[113556] = 12'h  0;
rom[113557] = 12'h  0;
rom[113558] = 12'h  0;
rom[113559] = 12'h  0;
rom[113560] = 12'h  0;
rom[113561] = 12'h  0;
rom[113562] = 12'h111;
rom[113563] = 12'h111;
rom[113564] = 12'h222;
rom[113565] = 12'h333;
rom[113566] = 12'h666;
rom[113567] = 12'h999;
rom[113568] = 12'hbbb;
rom[113569] = 12'haaa;
rom[113570] = 12'h777;
rom[113571] = 12'h444;
rom[113572] = 12'h222;
rom[113573] = 12'h222;
rom[113574] = 12'h222;
rom[113575] = 12'h111;
rom[113576] = 12'h111;
rom[113577] = 12'h  0;
rom[113578] = 12'h  0;
rom[113579] = 12'h  0;
rom[113580] = 12'h  0;
rom[113581] = 12'h  0;
rom[113582] = 12'h  0;
rom[113583] = 12'h  0;
rom[113584] = 12'h  0;
rom[113585] = 12'h  0;
rom[113586] = 12'h  0;
rom[113587] = 12'h  0;
rom[113588] = 12'h  0;
rom[113589] = 12'h  0;
rom[113590] = 12'h  0;
rom[113591] = 12'h  0;
rom[113592] = 12'h  0;
rom[113593] = 12'h  0;
rom[113594] = 12'h  0;
rom[113595] = 12'h  0;
rom[113596] = 12'h  0;
rom[113597] = 12'h  0;
rom[113598] = 12'h  0;
rom[113599] = 12'h  0;
rom[113600] = 12'hfff;
rom[113601] = 12'hfff;
rom[113602] = 12'hfff;
rom[113603] = 12'hfff;
rom[113604] = 12'hfff;
rom[113605] = 12'hfff;
rom[113606] = 12'hfff;
rom[113607] = 12'hfff;
rom[113608] = 12'hfff;
rom[113609] = 12'hfff;
rom[113610] = 12'hfff;
rom[113611] = 12'hfff;
rom[113612] = 12'hfff;
rom[113613] = 12'hfff;
rom[113614] = 12'hfff;
rom[113615] = 12'hfff;
rom[113616] = 12'hfff;
rom[113617] = 12'hfff;
rom[113618] = 12'hfff;
rom[113619] = 12'hfff;
rom[113620] = 12'hfff;
rom[113621] = 12'hfff;
rom[113622] = 12'hfff;
rom[113623] = 12'hfff;
rom[113624] = 12'hfff;
rom[113625] = 12'hfff;
rom[113626] = 12'hfff;
rom[113627] = 12'hfff;
rom[113628] = 12'hfff;
rom[113629] = 12'hfff;
rom[113630] = 12'hfff;
rom[113631] = 12'hfff;
rom[113632] = 12'hfff;
rom[113633] = 12'hfff;
rom[113634] = 12'heee;
rom[113635] = 12'heee;
rom[113636] = 12'heee;
rom[113637] = 12'heee;
rom[113638] = 12'heee;
rom[113639] = 12'heee;
rom[113640] = 12'heee;
rom[113641] = 12'heee;
rom[113642] = 12'heee;
rom[113643] = 12'heee;
rom[113644] = 12'heee;
rom[113645] = 12'heee;
rom[113646] = 12'hddd;
rom[113647] = 12'hddd;
rom[113648] = 12'hddd;
rom[113649] = 12'hddd;
rom[113650] = 12'hddd;
rom[113651] = 12'hddd;
rom[113652] = 12'hddd;
rom[113653] = 12'hddd;
rom[113654] = 12'hddd;
rom[113655] = 12'hddd;
rom[113656] = 12'hccc;
rom[113657] = 12'hccc;
rom[113658] = 12'hccc;
rom[113659] = 12'hccc;
rom[113660] = 12'hccc;
rom[113661] = 12'hccc;
rom[113662] = 12'hccc;
rom[113663] = 12'hccc;
rom[113664] = 12'hccc;
rom[113665] = 12'hccc;
rom[113666] = 12'hccc;
rom[113667] = 12'hccc;
rom[113668] = 12'hccc;
rom[113669] = 12'hbbb;
rom[113670] = 12'hbbb;
rom[113671] = 12'hccc;
rom[113672] = 12'hbbb;
rom[113673] = 12'hbbb;
rom[113674] = 12'hbbb;
rom[113675] = 12'hbbb;
rom[113676] = 12'hbbb;
rom[113677] = 12'hbbb;
rom[113678] = 12'hbbb;
rom[113679] = 12'hbbb;
rom[113680] = 12'hccc;
rom[113681] = 12'hddd;
rom[113682] = 12'heee;
rom[113683] = 12'heee;
rom[113684] = 12'heee;
rom[113685] = 12'heee;
rom[113686] = 12'heee;
rom[113687] = 12'hccc;
rom[113688] = 12'haaa;
rom[113689] = 12'haaa;
rom[113690] = 12'haaa;
rom[113691] = 12'h999;
rom[113692] = 12'haaa;
rom[113693] = 12'haaa;
rom[113694] = 12'haaa;
rom[113695] = 12'h999;
rom[113696] = 12'haaa;
rom[113697] = 12'h999;
rom[113698] = 12'h999;
rom[113699] = 12'haaa;
rom[113700] = 12'hbbb;
rom[113701] = 12'hbbb;
rom[113702] = 12'hccc;
rom[113703] = 12'hccc;
rom[113704] = 12'hccc;
rom[113705] = 12'hbbb;
rom[113706] = 12'haaa;
rom[113707] = 12'h999;
rom[113708] = 12'h999;
rom[113709] = 12'h999;
rom[113710] = 12'h999;
rom[113711] = 12'h999;
rom[113712] = 12'h888;
rom[113713] = 12'h888;
rom[113714] = 12'h888;
rom[113715] = 12'h888;
rom[113716] = 12'h888;
rom[113717] = 12'h888;
rom[113718] = 12'h888;
rom[113719] = 12'h888;
rom[113720] = 12'h888;
rom[113721] = 12'h777;
rom[113722] = 12'h888;
rom[113723] = 12'h888;
rom[113724] = 12'h888;
rom[113725] = 12'h777;
rom[113726] = 12'h666;
rom[113727] = 12'h555;
rom[113728] = 12'h666;
rom[113729] = 12'h666;
rom[113730] = 12'h777;
rom[113731] = 12'h777;
rom[113732] = 12'h777;
rom[113733] = 12'h777;
rom[113734] = 12'h666;
rom[113735] = 12'h666;
rom[113736] = 12'h666;
rom[113737] = 12'h666;
rom[113738] = 12'h666;
rom[113739] = 12'h666;
rom[113740] = 12'h777;
rom[113741] = 12'h777;
rom[113742] = 12'h666;
rom[113743] = 12'h555;
rom[113744] = 12'h555;
rom[113745] = 12'h555;
rom[113746] = 12'h555;
rom[113747] = 12'h555;
rom[113748] = 12'h555;
rom[113749] = 12'h666;
rom[113750] = 12'h666;
rom[113751] = 12'h666;
rom[113752] = 12'h666;
rom[113753] = 12'h666;
rom[113754] = 12'h666;
rom[113755] = 12'h666;
rom[113756] = 12'h777;
rom[113757] = 12'h777;
rom[113758] = 12'h777;
rom[113759] = 12'h777;
rom[113760] = 12'h888;
rom[113761] = 12'h888;
rom[113762] = 12'h888;
rom[113763] = 12'h999;
rom[113764] = 12'h999;
rom[113765] = 12'h999;
rom[113766] = 12'h999;
rom[113767] = 12'haaa;
rom[113768] = 12'h999;
rom[113769] = 12'haaa;
rom[113770] = 12'haaa;
rom[113771] = 12'haaa;
rom[113772] = 12'haaa;
rom[113773] = 12'hbbb;
rom[113774] = 12'hbbb;
rom[113775] = 12'hbbb;
rom[113776] = 12'hbbb;
rom[113777] = 12'hbbb;
rom[113778] = 12'hccc;
rom[113779] = 12'hccc;
rom[113780] = 12'hccc;
rom[113781] = 12'hddd;
rom[113782] = 12'hddd;
rom[113783] = 12'hddd;
rom[113784] = 12'hddd;
rom[113785] = 12'hddd;
rom[113786] = 12'heee;
rom[113787] = 12'heee;
rom[113788] = 12'heee;
rom[113789] = 12'heee;
rom[113790] = 12'heee;
rom[113791] = 12'heee;
rom[113792] = 12'hfff;
rom[113793] = 12'hfff;
rom[113794] = 12'hfff;
rom[113795] = 12'hfff;
rom[113796] = 12'hfff;
rom[113797] = 12'heee;
rom[113798] = 12'heee;
rom[113799] = 12'heee;
rom[113800] = 12'heee;
rom[113801] = 12'heee;
rom[113802] = 12'heee;
rom[113803] = 12'hddd;
rom[113804] = 12'hddd;
rom[113805] = 12'hddd;
rom[113806] = 12'hccc;
rom[113807] = 12'hccc;
rom[113808] = 12'hbbb;
rom[113809] = 12'haaa;
rom[113810] = 12'h999;
rom[113811] = 12'h999;
rom[113812] = 12'h888;
rom[113813] = 12'h888;
rom[113814] = 12'h888;
rom[113815] = 12'h888;
rom[113816] = 12'h888;
rom[113817] = 12'h777;
rom[113818] = 12'h666;
rom[113819] = 12'h555;
rom[113820] = 12'h666;
rom[113821] = 12'h888;
rom[113822] = 12'haaa;
rom[113823] = 12'haaa;
rom[113824] = 12'h777;
rom[113825] = 12'h555;
rom[113826] = 12'h444;
rom[113827] = 12'h333;
rom[113828] = 12'h222;
rom[113829] = 12'h222;
rom[113830] = 12'h333;
rom[113831] = 12'h333;
rom[113832] = 12'h444;
rom[113833] = 12'h444;
rom[113834] = 12'h444;
rom[113835] = 12'h333;
rom[113836] = 12'h222;
rom[113837] = 12'h222;
rom[113838] = 12'h222;
rom[113839] = 12'h333;
rom[113840] = 12'h333;
rom[113841] = 12'h444;
rom[113842] = 12'h777;
rom[113843] = 12'hccc;
rom[113844] = 12'hddd;
rom[113845] = 12'h999;
rom[113846] = 12'h444;
rom[113847] = 12'h111;
rom[113848] = 12'h111;
rom[113849] = 12'h111;
rom[113850] = 12'h111;
rom[113851] = 12'h  0;
rom[113852] = 12'h  0;
rom[113853] = 12'h  0;
rom[113854] = 12'h  0;
rom[113855] = 12'h  0;
rom[113856] = 12'h111;
rom[113857] = 12'h  0;
rom[113858] = 12'h  0;
rom[113859] = 12'h111;
rom[113860] = 12'h222;
rom[113861] = 12'h222;
rom[113862] = 12'h222;
rom[113863] = 12'h555;
rom[113864] = 12'hddd;
rom[113865] = 12'heee;
rom[113866] = 12'hbbb;
rom[113867] = 12'h666;
rom[113868] = 12'h333;
rom[113869] = 12'h222;
rom[113870] = 12'h111;
rom[113871] = 12'h111;
rom[113872] = 12'h111;
rom[113873] = 12'h222;
rom[113874] = 12'h777;
rom[113875] = 12'hddd;
rom[113876] = 12'hddd;
rom[113877] = 12'h666;
rom[113878] = 12'h111;
rom[113879] = 12'h  0;
rom[113880] = 12'h111;
rom[113881] = 12'h111;
rom[113882] = 12'h  0;
rom[113883] = 12'h  0;
rom[113884] = 12'h111;
rom[113885] = 12'h  0;
rom[113886] = 12'h  0;
rom[113887] = 12'h111;
rom[113888] = 12'h444;
rom[113889] = 12'h888;
rom[113890] = 12'h999;
rom[113891] = 12'h999;
rom[113892] = 12'hddd;
rom[113893] = 12'haaa;
rom[113894] = 12'h444;
rom[113895] = 12'h111;
rom[113896] = 12'h111;
rom[113897] = 12'h111;
rom[113898] = 12'h111;
rom[113899] = 12'h111;
rom[113900] = 12'h111;
rom[113901] = 12'h222;
rom[113902] = 12'h111;
rom[113903] = 12'h111;
rom[113904] = 12'h111;
rom[113905] = 12'h222;
rom[113906] = 12'h222;
rom[113907] = 12'h222;
rom[113908] = 12'h333;
rom[113909] = 12'h555;
rom[113910] = 12'h777;
rom[113911] = 12'h999;
rom[113912] = 12'hbbb;
rom[113913] = 12'hccc;
rom[113914] = 12'hbbb;
rom[113915] = 12'h888;
rom[113916] = 12'h555;
rom[113917] = 12'h333;
rom[113918] = 12'h222;
rom[113919] = 12'h222;
rom[113920] = 12'h222;
rom[113921] = 12'h222;
rom[113922] = 12'h222;
rom[113923] = 12'h111;
rom[113924] = 12'h111;
rom[113925] = 12'h111;
rom[113926] = 12'h  0;
rom[113927] = 12'h  0;
rom[113928] = 12'h  0;
rom[113929] = 12'h  0;
rom[113930] = 12'h  0;
rom[113931] = 12'h  0;
rom[113932] = 12'h  0;
rom[113933] = 12'h  0;
rom[113934] = 12'h  0;
rom[113935] = 12'h  0;
rom[113936] = 12'h  0;
rom[113937] = 12'h  0;
rom[113938] = 12'h  0;
rom[113939] = 12'h  0;
rom[113940] = 12'h  0;
rom[113941] = 12'h  0;
rom[113942] = 12'h  0;
rom[113943] = 12'h  0;
rom[113944] = 12'h  0;
rom[113945] = 12'h  0;
rom[113946] = 12'h  0;
rom[113947] = 12'h  0;
rom[113948] = 12'h  0;
rom[113949] = 12'h  0;
rom[113950] = 12'h  0;
rom[113951] = 12'h  0;
rom[113952] = 12'h  0;
rom[113953] = 12'h  0;
rom[113954] = 12'h  0;
rom[113955] = 12'h  0;
rom[113956] = 12'h  0;
rom[113957] = 12'h  0;
rom[113958] = 12'h  0;
rom[113959] = 12'h  0;
rom[113960] = 12'h  0;
rom[113961] = 12'h  0;
rom[113962] = 12'h  0;
rom[113963] = 12'h111;
rom[113964] = 12'h111;
rom[113965] = 12'h222;
rom[113966] = 12'h444;
rom[113967] = 12'h777;
rom[113968] = 12'hbbb;
rom[113969] = 12'hbbb;
rom[113970] = 12'h999;
rom[113971] = 12'h555;
rom[113972] = 12'h222;
rom[113973] = 12'h222;
rom[113974] = 12'h222;
rom[113975] = 12'h111;
rom[113976] = 12'h111;
rom[113977] = 12'h111;
rom[113978] = 12'h  0;
rom[113979] = 12'h  0;
rom[113980] = 12'h  0;
rom[113981] = 12'h  0;
rom[113982] = 12'h  0;
rom[113983] = 12'h  0;
rom[113984] = 12'h  0;
rom[113985] = 12'h  0;
rom[113986] = 12'h  0;
rom[113987] = 12'h  0;
rom[113988] = 12'h  0;
rom[113989] = 12'h  0;
rom[113990] = 12'h  0;
rom[113991] = 12'h  0;
rom[113992] = 12'h  0;
rom[113993] = 12'h  0;
rom[113994] = 12'h  0;
rom[113995] = 12'h  0;
rom[113996] = 12'h  0;
rom[113997] = 12'h  0;
rom[113998] = 12'h  0;
rom[113999] = 12'h  0;
rom[114000] = 12'hfff;
rom[114001] = 12'hfff;
rom[114002] = 12'hfff;
rom[114003] = 12'hfff;
rom[114004] = 12'hfff;
rom[114005] = 12'hfff;
rom[114006] = 12'hfff;
rom[114007] = 12'hfff;
rom[114008] = 12'hfff;
rom[114009] = 12'hfff;
rom[114010] = 12'hfff;
rom[114011] = 12'hfff;
rom[114012] = 12'hfff;
rom[114013] = 12'hfff;
rom[114014] = 12'hfff;
rom[114015] = 12'hfff;
rom[114016] = 12'hfff;
rom[114017] = 12'hfff;
rom[114018] = 12'hfff;
rom[114019] = 12'hfff;
rom[114020] = 12'hfff;
rom[114021] = 12'hfff;
rom[114022] = 12'hfff;
rom[114023] = 12'hfff;
rom[114024] = 12'hfff;
rom[114025] = 12'hfff;
rom[114026] = 12'hfff;
rom[114027] = 12'hfff;
rom[114028] = 12'hfff;
rom[114029] = 12'hfff;
rom[114030] = 12'hfff;
rom[114031] = 12'hfff;
rom[114032] = 12'heee;
rom[114033] = 12'heee;
rom[114034] = 12'heee;
rom[114035] = 12'heee;
rom[114036] = 12'heee;
rom[114037] = 12'heee;
rom[114038] = 12'heee;
rom[114039] = 12'heee;
rom[114040] = 12'heee;
rom[114041] = 12'heee;
rom[114042] = 12'heee;
rom[114043] = 12'heee;
rom[114044] = 12'heee;
rom[114045] = 12'hddd;
rom[114046] = 12'hddd;
rom[114047] = 12'hddd;
rom[114048] = 12'hddd;
rom[114049] = 12'hddd;
rom[114050] = 12'hddd;
rom[114051] = 12'hddd;
rom[114052] = 12'hddd;
rom[114053] = 12'hddd;
rom[114054] = 12'hccc;
rom[114055] = 12'hccc;
rom[114056] = 12'hccc;
rom[114057] = 12'hccc;
rom[114058] = 12'hccc;
rom[114059] = 12'hccc;
rom[114060] = 12'hccc;
rom[114061] = 12'hccc;
rom[114062] = 12'hccc;
rom[114063] = 12'hccc;
rom[114064] = 12'hccc;
rom[114065] = 12'hccc;
rom[114066] = 12'hccc;
rom[114067] = 12'hccc;
rom[114068] = 12'hbbb;
rom[114069] = 12'hbbb;
rom[114070] = 12'hbbb;
rom[114071] = 12'hbbb;
rom[114072] = 12'hbbb;
rom[114073] = 12'hbbb;
rom[114074] = 12'hbbb;
rom[114075] = 12'hbbb;
rom[114076] = 12'hbbb;
rom[114077] = 12'hbbb;
rom[114078] = 12'hbbb;
rom[114079] = 12'hbbb;
rom[114080] = 12'hddd;
rom[114081] = 12'heee;
rom[114082] = 12'hfff;
rom[114083] = 12'heee;
rom[114084] = 12'heee;
rom[114085] = 12'heee;
rom[114086] = 12'hddd;
rom[114087] = 12'haaa;
rom[114088] = 12'haaa;
rom[114089] = 12'haaa;
rom[114090] = 12'haaa;
rom[114091] = 12'haaa;
rom[114092] = 12'h999;
rom[114093] = 12'haaa;
rom[114094] = 12'haaa;
rom[114095] = 12'haaa;
rom[114096] = 12'haaa;
rom[114097] = 12'h999;
rom[114098] = 12'h999;
rom[114099] = 12'haaa;
rom[114100] = 12'hbbb;
rom[114101] = 12'hccc;
rom[114102] = 12'hccc;
rom[114103] = 12'hccc;
rom[114104] = 12'hbbb;
rom[114105] = 12'hbbb;
rom[114106] = 12'haaa;
rom[114107] = 12'h999;
rom[114108] = 12'h888;
rom[114109] = 12'h999;
rom[114110] = 12'h999;
rom[114111] = 12'h888;
rom[114112] = 12'h888;
rom[114113] = 12'h888;
rom[114114] = 12'h888;
rom[114115] = 12'h888;
rom[114116] = 12'h777;
rom[114117] = 12'h777;
rom[114118] = 12'h777;
rom[114119] = 12'h888;
rom[114120] = 12'h777;
rom[114121] = 12'h777;
rom[114122] = 12'h888;
rom[114123] = 12'h888;
rom[114124] = 12'h888;
rom[114125] = 12'h777;
rom[114126] = 12'h666;
rom[114127] = 12'h666;
rom[114128] = 12'h666;
rom[114129] = 12'h666;
rom[114130] = 12'h777;
rom[114131] = 12'h777;
rom[114132] = 12'h777;
rom[114133] = 12'h666;
rom[114134] = 12'h666;
rom[114135] = 12'h666;
rom[114136] = 12'h666;
rom[114137] = 12'h666;
rom[114138] = 12'h666;
rom[114139] = 12'h777;
rom[114140] = 12'h777;
rom[114141] = 12'h666;
rom[114142] = 12'h666;
rom[114143] = 12'h555;
rom[114144] = 12'h555;
rom[114145] = 12'h555;
rom[114146] = 12'h555;
rom[114147] = 12'h555;
rom[114148] = 12'h555;
rom[114149] = 12'h555;
rom[114150] = 12'h666;
rom[114151] = 12'h666;
rom[114152] = 12'h666;
rom[114153] = 12'h666;
rom[114154] = 12'h666;
rom[114155] = 12'h666;
rom[114156] = 12'h666;
rom[114157] = 12'h777;
rom[114158] = 12'h777;
rom[114159] = 12'h777;
rom[114160] = 12'h888;
rom[114161] = 12'h888;
rom[114162] = 12'h888;
rom[114163] = 12'h888;
rom[114164] = 12'h888;
rom[114165] = 12'h888;
rom[114166] = 12'h888;
rom[114167] = 12'h999;
rom[114168] = 12'h888;
rom[114169] = 12'h888;
rom[114170] = 12'h999;
rom[114171] = 12'h999;
rom[114172] = 12'h999;
rom[114173] = 12'haaa;
rom[114174] = 12'haaa;
rom[114175] = 12'haaa;
rom[114176] = 12'haaa;
rom[114177] = 12'haaa;
rom[114178] = 12'haaa;
rom[114179] = 12'haaa;
rom[114180] = 12'hbbb;
rom[114181] = 12'hbbb;
rom[114182] = 12'hbbb;
rom[114183] = 12'hbbb;
rom[114184] = 12'hbbb;
rom[114185] = 12'hccc;
rom[114186] = 12'hccc;
rom[114187] = 12'hccc;
rom[114188] = 12'hccc;
rom[114189] = 12'hddd;
rom[114190] = 12'hddd;
rom[114191] = 12'hddd;
rom[114192] = 12'hddd;
rom[114193] = 12'hddd;
rom[114194] = 12'hddd;
rom[114195] = 12'hddd;
rom[114196] = 12'hddd;
rom[114197] = 12'hddd;
rom[114198] = 12'hddd;
rom[114199] = 12'hccc;
rom[114200] = 12'hccc;
rom[114201] = 12'hccc;
rom[114202] = 12'hccc;
rom[114203] = 12'hbbb;
rom[114204] = 12'hbbb;
rom[114205] = 12'hbbb;
rom[114206] = 12'haaa;
rom[114207] = 12'haaa;
rom[114208] = 12'haaa;
rom[114209] = 12'h999;
rom[114210] = 12'h999;
rom[114211] = 12'h888;
rom[114212] = 12'h888;
rom[114213] = 12'h777;
rom[114214] = 12'h777;
rom[114215] = 12'h888;
rom[114216] = 12'h777;
rom[114217] = 12'h777;
rom[114218] = 12'h666;
rom[114219] = 12'h555;
rom[114220] = 12'h555;
rom[114221] = 12'h666;
rom[114222] = 12'h888;
rom[114223] = 12'haaa;
rom[114224] = 12'h888;
rom[114225] = 12'h666;
rom[114226] = 12'h444;
rom[114227] = 12'h222;
rom[114228] = 12'h222;
rom[114229] = 12'h222;
rom[114230] = 12'h222;
rom[114231] = 12'h222;
rom[114232] = 12'h444;
rom[114233] = 12'h444;
rom[114234] = 12'h444;
rom[114235] = 12'h333;
rom[114236] = 12'h222;
rom[114237] = 12'h111;
rom[114238] = 12'h222;
rom[114239] = 12'h222;
rom[114240] = 12'h333;
rom[114241] = 12'h555;
rom[114242] = 12'h999;
rom[114243] = 12'hccc;
rom[114244] = 12'hbbb;
rom[114245] = 12'h666;
rom[114246] = 12'h333;
rom[114247] = 12'h111;
rom[114248] = 12'h111;
rom[114249] = 12'h111;
rom[114250] = 12'h  0;
rom[114251] = 12'h  0;
rom[114252] = 12'h  0;
rom[114253] = 12'h  0;
rom[114254] = 12'h  0;
rom[114255] = 12'h  0;
rom[114256] = 12'h  0;
rom[114257] = 12'h  0;
rom[114258] = 12'h  0;
rom[114259] = 12'h111;
rom[114260] = 12'h222;
rom[114261] = 12'h111;
rom[114262] = 12'h111;
rom[114263] = 12'h444;
rom[114264] = 12'hccc;
rom[114265] = 12'heee;
rom[114266] = 12'hbbb;
rom[114267] = 12'h666;
rom[114268] = 12'h333;
rom[114269] = 12'h222;
rom[114270] = 12'h111;
rom[114271] = 12'h111;
rom[114272] = 12'h111;
rom[114273] = 12'h111;
rom[114274] = 12'h555;
rom[114275] = 12'hbbb;
rom[114276] = 12'heee;
rom[114277] = 12'h888;
rom[114278] = 12'h222;
rom[114279] = 12'h  0;
rom[114280] = 12'h111;
rom[114281] = 12'h111;
rom[114282] = 12'h  0;
rom[114283] = 12'h  0;
rom[114284] = 12'h  0;
rom[114285] = 12'h111;
rom[114286] = 12'h  0;
rom[114287] = 12'h111;
rom[114288] = 12'h333;
rom[114289] = 12'h888;
rom[114290] = 12'h999;
rom[114291] = 12'h888;
rom[114292] = 12'hccc;
rom[114293] = 12'hbbb;
rom[114294] = 12'h666;
rom[114295] = 12'h222;
rom[114296] = 12'h111;
rom[114297] = 12'h111;
rom[114298] = 12'h111;
rom[114299] = 12'h111;
rom[114300] = 12'h111;
rom[114301] = 12'h111;
rom[114302] = 12'h111;
rom[114303] = 12'h  0;
rom[114304] = 12'h111;
rom[114305] = 12'h111;
rom[114306] = 12'h222;
rom[114307] = 12'h222;
rom[114308] = 12'h222;
rom[114309] = 12'h444;
rom[114310] = 12'h666;
rom[114311] = 12'h888;
rom[114312] = 12'haaa;
rom[114313] = 12'hbbb;
rom[114314] = 12'hbbb;
rom[114315] = 12'haaa;
rom[114316] = 12'h777;
rom[114317] = 12'h444;
rom[114318] = 12'h222;
rom[114319] = 12'h222;
rom[114320] = 12'h222;
rom[114321] = 12'h222;
rom[114322] = 12'h111;
rom[114323] = 12'h111;
rom[114324] = 12'h111;
rom[114325] = 12'h  0;
rom[114326] = 12'h  0;
rom[114327] = 12'h  0;
rom[114328] = 12'h  0;
rom[114329] = 12'h  0;
rom[114330] = 12'h  0;
rom[114331] = 12'h  0;
rom[114332] = 12'h  0;
rom[114333] = 12'h  0;
rom[114334] = 12'h  0;
rom[114335] = 12'h  0;
rom[114336] = 12'h  0;
rom[114337] = 12'h  0;
rom[114338] = 12'h  0;
rom[114339] = 12'h  0;
rom[114340] = 12'h  0;
rom[114341] = 12'h  0;
rom[114342] = 12'h  0;
rom[114343] = 12'h  0;
rom[114344] = 12'h  0;
rom[114345] = 12'h  0;
rom[114346] = 12'h  0;
rom[114347] = 12'h  0;
rom[114348] = 12'h  0;
rom[114349] = 12'h  0;
rom[114350] = 12'h  0;
rom[114351] = 12'h  0;
rom[114352] = 12'h  0;
rom[114353] = 12'h  0;
rom[114354] = 12'h  0;
rom[114355] = 12'h  0;
rom[114356] = 12'h  0;
rom[114357] = 12'h  0;
rom[114358] = 12'h  0;
rom[114359] = 12'h  0;
rom[114360] = 12'h  0;
rom[114361] = 12'h  0;
rom[114362] = 12'h  0;
rom[114363] = 12'h  0;
rom[114364] = 12'h111;
rom[114365] = 12'h111;
rom[114366] = 12'h333;
rom[114367] = 12'h555;
rom[114368] = 12'h999;
rom[114369] = 12'hbbb;
rom[114370] = 12'haaa;
rom[114371] = 12'h777;
rom[114372] = 12'h444;
rom[114373] = 12'h222;
rom[114374] = 12'h222;
rom[114375] = 12'h111;
rom[114376] = 12'h111;
rom[114377] = 12'h111;
rom[114378] = 12'h  0;
rom[114379] = 12'h  0;
rom[114380] = 12'h  0;
rom[114381] = 12'h  0;
rom[114382] = 12'h  0;
rom[114383] = 12'h  0;
rom[114384] = 12'h  0;
rom[114385] = 12'h  0;
rom[114386] = 12'h  0;
rom[114387] = 12'h  0;
rom[114388] = 12'h  0;
rom[114389] = 12'h  0;
rom[114390] = 12'h  0;
rom[114391] = 12'h  0;
rom[114392] = 12'h  0;
rom[114393] = 12'h  0;
rom[114394] = 12'h  0;
rom[114395] = 12'h  0;
rom[114396] = 12'h  0;
rom[114397] = 12'h  0;
rom[114398] = 12'h  0;
rom[114399] = 12'h  0;
rom[114400] = 12'hfff;
rom[114401] = 12'hfff;
rom[114402] = 12'hfff;
rom[114403] = 12'hfff;
rom[114404] = 12'hfff;
rom[114405] = 12'hfff;
rom[114406] = 12'hfff;
rom[114407] = 12'hfff;
rom[114408] = 12'hfff;
rom[114409] = 12'hfff;
rom[114410] = 12'hfff;
rom[114411] = 12'hfff;
rom[114412] = 12'hfff;
rom[114413] = 12'hfff;
rom[114414] = 12'hfff;
rom[114415] = 12'hfff;
rom[114416] = 12'hfff;
rom[114417] = 12'hfff;
rom[114418] = 12'hfff;
rom[114419] = 12'hfff;
rom[114420] = 12'hfff;
rom[114421] = 12'hfff;
rom[114422] = 12'hfff;
rom[114423] = 12'heee;
rom[114424] = 12'heee;
rom[114425] = 12'heee;
rom[114426] = 12'heee;
rom[114427] = 12'heee;
rom[114428] = 12'heee;
rom[114429] = 12'heee;
rom[114430] = 12'heee;
rom[114431] = 12'heee;
rom[114432] = 12'heee;
rom[114433] = 12'heee;
rom[114434] = 12'heee;
rom[114435] = 12'heee;
rom[114436] = 12'heee;
rom[114437] = 12'heee;
rom[114438] = 12'heee;
rom[114439] = 12'heee;
rom[114440] = 12'heee;
rom[114441] = 12'heee;
rom[114442] = 12'heee;
rom[114443] = 12'heee;
rom[114444] = 12'hddd;
rom[114445] = 12'hddd;
rom[114446] = 12'hddd;
rom[114447] = 12'hddd;
rom[114448] = 12'hddd;
rom[114449] = 12'hddd;
rom[114450] = 12'hddd;
rom[114451] = 12'hddd;
rom[114452] = 12'hddd;
rom[114453] = 12'hccc;
rom[114454] = 12'hccc;
rom[114455] = 12'hccc;
rom[114456] = 12'hccc;
rom[114457] = 12'hccc;
rom[114458] = 12'hccc;
rom[114459] = 12'hccc;
rom[114460] = 12'hccc;
rom[114461] = 12'hccc;
rom[114462] = 12'hccc;
rom[114463] = 12'hccc;
rom[114464] = 12'hddd;
rom[114465] = 12'hccc;
rom[114466] = 12'hccc;
rom[114467] = 12'hbbb;
rom[114468] = 12'hbbb;
rom[114469] = 12'hbbb;
rom[114470] = 12'hbbb;
rom[114471] = 12'hbbb;
rom[114472] = 12'hbbb;
rom[114473] = 12'hbbb;
rom[114474] = 12'hbbb;
rom[114475] = 12'hbbb;
rom[114476] = 12'hbbb;
rom[114477] = 12'hbbb;
rom[114478] = 12'hbbb;
rom[114479] = 12'hccc;
rom[114480] = 12'heee;
rom[114481] = 12'heee;
rom[114482] = 12'hfff;
rom[114483] = 12'hfff;
rom[114484] = 12'heee;
rom[114485] = 12'hccc;
rom[114486] = 12'hbbb;
rom[114487] = 12'haaa;
rom[114488] = 12'haaa;
rom[114489] = 12'haaa;
rom[114490] = 12'haaa;
rom[114491] = 12'haaa;
rom[114492] = 12'haaa;
rom[114493] = 12'haaa;
rom[114494] = 12'haaa;
rom[114495] = 12'haaa;
rom[114496] = 12'haaa;
rom[114497] = 12'h999;
rom[114498] = 12'h999;
rom[114499] = 12'haaa;
rom[114500] = 12'hbbb;
rom[114501] = 12'hccc;
rom[114502] = 12'hccc;
rom[114503] = 12'hbbb;
rom[114504] = 12'haaa;
rom[114505] = 12'haaa;
rom[114506] = 12'h999;
rom[114507] = 12'h888;
rom[114508] = 12'h888;
rom[114509] = 12'h888;
rom[114510] = 12'h888;
rom[114511] = 12'h888;
rom[114512] = 12'h777;
rom[114513] = 12'h777;
rom[114514] = 12'h777;
rom[114515] = 12'h777;
rom[114516] = 12'h777;
rom[114517] = 12'h777;
rom[114518] = 12'h777;
rom[114519] = 12'h777;
rom[114520] = 12'h777;
rom[114521] = 12'h777;
rom[114522] = 12'h888;
rom[114523] = 12'h888;
rom[114524] = 12'h777;
rom[114525] = 12'h666;
rom[114526] = 12'h555;
rom[114527] = 12'h666;
rom[114528] = 12'h666;
rom[114529] = 12'h666;
rom[114530] = 12'h777;
rom[114531] = 12'h777;
rom[114532] = 12'h666;
rom[114533] = 12'h555;
rom[114534] = 12'h555;
rom[114535] = 12'h666;
rom[114536] = 12'h666;
rom[114537] = 12'h666;
rom[114538] = 12'h666;
rom[114539] = 12'h777;
rom[114540] = 12'h666;
rom[114541] = 12'h555;
rom[114542] = 12'h555;
rom[114543] = 12'h555;
rom[114544] = 12'h555;
rom[114545] = 12'h555;
rom[114546] = 12'h555;
rom[114547] = 12'h555;
rom[114548] = 12'h555;
rom[114549] = 12'h555;
rom[114550] = 12'h555;
rom[114551] = 12'h555;
rom[114552] = 12'h555;
rom[114553] = 12'h555;
rom[114554] = 12'h555;
rom[114555] = 12'h555;
rom[114556] = 12'h666;
rom[114557] = 12'h666;
rom[114558] = 12'h777;
rom[114559] = 12'h777;
rom[114560] = 12'h888;
rom[114561] = 12'h888;
rom[114562] = 12'h888;
rom[114563] = 12'h888;
rom[114564] = 12'h888;
rom[114565] = 12'h888;
rom[114566] = 12'h888;
rom[114567] = 12'h888;
rom[114568] = 12'h888;
rom[114569] = 12'h888;
rom[114570] = 12'h888;
rom[114571] = 12'h888;
rom[114572] = 12'h999;
rom[114573] = 12'h999;
rom[114574] = 12'h999;
rom[114575] = 12'h999;
rom[114576] = 12'h999;
rom[114577] = 12'h999;
rom[114578] = 12'h999;
rom[114579] = 12'h999;
rom[114580] = 12'h999;
rom[114581] = 12'haaa;
rom[114582] = 12'haaa;
rom[114583] = 12'haaa;
rom[114584] = 12'haaa;
rom[114585] = 12'haaa;
rom[114586] = 12'haaa;
rom[114587] = 12'haaa;
rom[114588] = 12'hbbb;
rom[114589] = 12'hbbb;
rom[114590] = 12'hbbb;
rom[114591] = 12'hbbb;
rom[114592] = 12'hbbb;
rom[114593] = 12'hbbb;
rom[114594] = 12'hbbb;
rom[114595] = 12'hbbb;
rom[114596] = 12'hbbb;
rom[114597] = 12'hbbb;
rom[114598] = 12'hbbb;
rom[114599] = 12'hbbb;
rom[114600] = 12'haaa;
rom[114601] = 12'haaa;
rom[114602] = 12'haaa;
rom[114603] = 12'haaa;
rom[114604] = 12'h999;
rom[114605] = 12'h999;
rom[114606] = 12'h999;
rom[114607] = 12'h999;
rom[114608] = 12'h999;
rom[114609] = 12'h888;
rom[114610] = 12'h888;
rom[114611] = 12'h888;
rom[114612] = 12'h777;
rom[114613] = 12'h777;
rom[114614] = 12'h777;
rom[114615] = 12'h777;
rom[114616] = 12'h777;
rom[114617] = 12'h666;
rom[114618] = 12'h555;
rom[114619] = 12'h444;
rom[114620] = 12'h444;
rom[114621] = 12'h444;
rom[114622] = 12'h666;
rom[114623] = 12'h999;
rom[114624] = 12'haaa;
rom[114625] = 12'h777;
rom[114626] = 12'h444;
rom[114627] = 12'h222;
rom[114628] = 12'h222;
rom[114629] = 12'h222;
rom[114630] = 12'h111;
rom[114631] = 12'h111;
rom[114632] = 12'h222;
rom[114633] = 12'h333;
rom[114634] = 12'h444;
rom[114635] = 12'h333;
rom[114636] = 12'h222;
rom[114637] = 12'h111;
rom[114638] = 12'h111;
rom[114639] = 12'h222;
rom[114640] = 12'h333;
rom[114641] = 12'h666;
rom[114642] = 12'haaa;
rom[114643] = 12'hccc;
rom[114644] = 12'h999;
rom[114645] = 12'h444;
rom[114646] = 12'h111;
rom[114647] = 12'h111;
rom[114648] = 12'h111;
rom[114649] = 12'h111;
rom[114650] = 12'h  0;
rom[114651] = 12'h  0;
rom[114652] = 12'h  0;
rom[114653] = 12'h  0;
rom[114654] = 12'h  0;
rom[114655] = 12'h  0;
rom[114656] = 12'h  0;
rom[114657] = 12'h  0;
rom[114658] = 12'h  0;
rom[114659] = 12'h111;
rom[114660] = 12'h111;
rom[114661] = 12'h111;
rom[114662] = 12'h111;
rom[114663] = 12'h444;
rom[114664] = 12'hccc;
rom[114665] = 12'heee;
rom[114666] = 12'hbbb;
rom[114667] = 12'h666;
rom[114668] = 12'h333;
rom[114669] = 12'h222;
rom[114670] = 12'h111;
rom[114671] = 12'h111;
rom[114672] = 12'h111;
rom[114673] = 12'h111;
rom[114674] = 12'h444;
rom[114675] = 12'h999;
rom[114676] = 12'heee;
rom[114677] = 12'h999;
rom[114678] = 12'h333;
rom[114679] = 12'h  0;
rom[114680] = 12'h  0;
rom[114681] = 12'h111;
rom[114682] = 12'h  0;
rom[114683] = 12'h  0;
rom[114684] = 12'h  0;
rom[114685] = 12'h111;
rom[114686] = 12'h  0;
rom[114687] = 12'h  0;
rom[114688] = 12'h111;
rom[114689] = 12'h666;
rom[114690] = 12'h888;
rom[114691] = 12'h888;
rom[114692] = 12'h888;
rom[114693] = 12'hbbb;
rom[114694] = 12'h999;
rom[114695] = 12'h444;
rom[114696] = 12'h111;
rom[114697] = 12'h111;
rom[114698] = 12'h111;
rom[114699] = 12'h111;
rom[114700] = 12'h111;
rom[114701] = 12'h111;
rom[114702] = 12'h111;
rom[114703] = 12'h111;
rom[114704] = 12'h111;
rom[114705] = 12'h111;
rom[114706] = 12'h111;
rom[114707] = 12'h222;
rom[114708] = 12'h222;
rom[114709] = 12'h222;
rom[114710] = 12'h444;
rom[114711] = 12'h666;
rom[114712] = 12'h888;
rom[114713] = 12'h999;
rom[114714] = 12'hbbb;
rom[114715] = 12'hbbb;
rom[114716] = 12'h999;
rom[114717] = 12'h555;
rom[114718] = 12'h333;
rom[114719] = 12'h222;
rom[114720] = 12'h222;
rom[114721] = 12'h222;
rom[114722] = 12'h111;
rom[114723] = 12'h111;
rom[114724] = 12'h111;
rom[114725] = 12'h  0;
rom[114726] = 12'h  0;
rom[114727] = 12'h  0;
rom[114728] = 12'h  0;
rom[114729] = 12'h  0;
rom[114730] = 12'h  0;
rom[114731] = 12'h  0;
rom[114732] = 12'h  0;
rom[114733] = 12'h  0;
rom[114734] = 12'h  0;
rom[114735] = 12'h  0;
rom[114736] = 12'h  0;
rom[114737] = 12'h  0;
rom[114738] = 12'h  0;
rom[114739] = 12'h  0;
rom[114740] = 12'h  0;
rom[114741] = 12'h  0;
rom[114742] = 12'h  0;
rom[114743] = 12'h  0;
rom[114744] = 12'h  0;
rom[114745] = 12'h  0;
rom[114746] = 12'h  0;
rom[114747] = 12'h  0;
rom[114748] = 12'h  0;
rom[114749] = 12'h  0;
rom[114750] = 12'h  0;
rom[114751] = 12'h  0;
rom[114752] = 12'h  0;
rom[114753] = 12'h  0;
rom[114754] = 12'h  0;
rom[114755] = 12'h  0;
rom[114756] = 12'h  0;
rom[114757] = 12'h  0;
rom[114758] = 12'h  0;
rom[114759] = 12'h  0;
rom[114760] = 12'h  0;
rom[114761] = 12'h  0;
rom[114762] = 12'h  0;
rom[114763] = 12'h  0;
rom[114764] = 12'h  0;
rom[114765] = 12'h  0;
rom[114766] = 12'h222;
rom[114767] = 12'h333;
rom[114768] = 12'h777;
rom[114769] = 12'haaa;
rom[114770] = 12'hbbb;
rom[114771] = 12'h999;
rom[114772] = 12'h555;
rom[114773] = 12'h333;
rom[114774] = 12'h222;
rom[114775] = 12'h111;
rom[114776] = 12'h111;
rom[114777] = 12'h111;
rom[114778] = 12'h  0;
rom[114779] = 12'h  0;
rom[114780] = 12'h  0;
rom[114781] = 12'h  0;
rom[114782] = 12'h  0;
rom[114783] = 12'h  0;
rom[114784] = 12'h  0;
rom[114785] = 12'h  0;
rom[114786] = 12'h  0;
rom[114787] = 12'h  0;
rom[114788] = 12'h  0;
rom[114789] = 12'h  0;
rom[114790] = 12'h  0;
rom[114791] = 12'h  0;
rom[114792] = 12'h  0;
rom[114793] = 12'h  0;
rom[114794] = 12'h  0;
rom[114795] = 12'h  0;
rom[114796] = 12'h  0;
rom[114797] = 12'h  0;
rom[114798] = 12'h  0;
rom[114799] = 12'h  0;
rom[114800] = 12'hfff;
rom[114801] = 12'hfff;
rom[114802] = 12'hfff;
rom[114803] = 12'hfff;
rom[114804] = 12'hfff;
rom[114805] = 12'hfff;
rom[114806] = 12'hfff;
rom[114807] = 12'hfff;
rom[114808] = 12'hfff;
rom[114809] = 12'hfff;
rom[114810] = 12'hfff;
rom[114811] = 12'hfff;
rom[114812] = 12'hfff;
rom[114813] = 12'hfff;
rom[114814] = 12'hfff;
rom[114815] = 12'hfff;
rom[114816] = 12'hfff;
rom[114817] = 12'hfff;
rom[114818] = 12'hfff;
rom[114819] = 12'hfff;
rom[114820] = 12'hfff;
rom[114821] = 12'hfff;
rom[114822] = 12'heee;
rom[114823] = 12'heee;
rom[114824] = 12'heee;
rom[114825] = 12'heee;
rom[114826] = 12'heee;
rom[114827] = 12'heee;
rom[114828] = 12'heee;
rom[114829] = 12'heee;
rom[114830] = 12'heee;
rom[114831] = 12'heee;
rom[114832] = 12'heee;
rom[114833] = 12'heee;
rom[114834] = 12'heee;
rom[114835] = 12'heee;
rom[114836] = 12'heee;
rom[114837] = 12'heee;
rom[114838] = 12'heee;
rom[114839] = 12'heee;
rom[114840] = 12'heee;
rom[114841] = 12'heee;
rom[114842] = 12'heee;
rom[114843] = 12'heee;
rom[114844] = 12'hddd;
rom[114845] = 12'hddd;
rom[114846] = 12'hddd;
rom[114847] = 12'hddd;
rom[114848] = 12'hddd;
rom[114849] = 12'hddd;
rom[114850] = 12'hddd;
rom[114851] = 12'hddd;
rom[114852] = 12'hddd;
rom[114853] = 12'hccc;
rom[114854] = 12'hccc;
rom[114855] = 12'hccc;
rom[114856] = 12'hccc;
rom[114857] = 12'hccc;
rom[114858] = 12'hccc;
rom[114859] = 12'hccc;
rom[114860] = 12'hccc;
rom[114861] = 12'hccc;
rom[114862] = 12'hccc;
rom[114863] = 12'hccc;
rom[114864] = 12'hddd;
rom[114865] = 12'hccc;
rom[114866] = 12'hbbb;
rom[114867] = 12'hbbb;
rom[114868] = 12'hbbb;
rom[114869] = 12'hbbb;
rom[114870] = 12'hbbb;
rom[114871] = 12'hbbb;
rom[114872] = 12'hbbb;
rom[114873] = 12'hbbb;
rom[114874] = 12'hbbb;
rom[114875] = 12'hbbb;
rom[114876] = 12'hbbb;
rom[114877] = 12'hbbb;
rom[114878] = 12'hccc;
rom[114879] = 12'hddd;
rom[114880] = 12'heee;
rom[114881] = 12'heee;
rom[114882] = 12'hfff;
rom[114883] = 12'hfff;
rom[114884] = 12'hddd;
rom[114885] = 12'hbbb;
rom[114886] = 12'haaa;
rom[114887] = 12'haaa;
rom[114888] = 12'haaa;
rom[114889] = 12'haaa;
rom[114890] = 12'haaa;
rom[114891] = 12'hbbb;
rom[114892] = 12'haaa;
rom[114893] = 12'h999;
rom[114894] = 12'h999;
rom[114895] = 12'haaa;
rom[114896] = 12'haaa;
rom[114897] = 12'h999;
rom[114898] = 12'haaa;
rom[114899] = 12'haaa;
rom[114900] = 12'hccc;
rom[114901] = 12'hccc;
rom[114902] = 12'hbbb;
rom[114903] = 12'haaa;
rom[114904] = 12'haaa;
rom[114905] = 12'haaa;
rom[114906] = 12'h999;
rom[114907] = 12'h888;
rom[114908] = 12'h888;
rom[114909] = 12'h888;
rom[114910] = 12'h888;
rom[114911] = 12'h888;
rom[114912] = 12'h777;
rom[114913] = 12'h777;
rom[114914] = 12'h777;
rom[114915] = 12'h777;
rom[114916] = 12'h777;
rom[114917] = 12'h777;
rom[114918] = 12'h777;
rom[114919] = 12'h777;
rom[114920] = 12'h777;
rom[114921] = 12'h777;
rom[114922] = 12'h888;
rom[114923] = 12'h888;
rom[114924] = 12'h777;
rom[114925] = 12'h555;
rom[114926] = 12'h555;
rom[114927] = 12'h666;
rom[114928] = 12'h666;
rom[114929] = 12'h666;
rom[114930] = 12'h777;
rom[114931] = 12'h777;
rom[114932] = 12'h666;
rom[114933] = 12'h555;
rom[114934] = 12'h555;
rom[114935] = 12'h666;
rom[114936] = 12'h666;
rom[114937] = 12'h555;
rom[114938] = 12'h666;
rom[114939] = 12'h777;
rom[114940] = 12'h666;
rom[114941] = 12'h444;
rom[114942] = 12'h444;
rom[114943] = 12'h555;
rom[114944] = 12'h555;
rom[114945] = 12'h555;
rom[114946] = 12'h555;
rom[114947] = 12'h444;
rom[114948] = 12'h444;
rom[114949] = 12'h555;
rom[114950] = 12'h555;
rom[114951] = 12'h555;
rom[114952] = 12'h555;
rom[114953] = 12'h555;
rom[114954] = 12'h555;
rom[114955] = 12'h555;
rom[114956] = 12'h555;
rom[114957] = 12'h666;
rom[114958] = 12'h666;
rom[114959] = 12'h777;
rom[114960] = 12'h777;
rom[114961] = 12'h777;
rom[114962] = 12'h777;
rom[114963] = 12'h777;
rom[114964] = 12'h777;
rom[114965] = 12'h777;
rom[114966] = 12'h777;
rom[114967] = 12'h777;
rom[114968] = 12'h888;
rom[114969] = 12'h888;
rom[114970] = 12'h888;
rom[114971] = 12'h888;
rom[114972] = 12'h888;
rom[114973] = 12'h999;
rom[114974] = 12'h999;
rom[114975] = 12'h999;
rom[114976] = 12'h999;
rom[114977] = 12'h999;
rom[114978] = 12'h999;
rom[114979] = 12'h999;
rom[114980] = 12'h999;
rom[114981] = 12'h999;
rom[114982] = 12'h999;
rom[114983] = 12'h999;
rom[114984] = 12'h999;
rom[114985] = 12'h999;
rom[114986] = 12'h999;
rom[114987] = 12'h999;
rom[114988] = 12'haaa;
rom[114989] = 12'haaa;
rom[114990] = 12'haaa;
rom[114991] = 12'haaa;
rom[114992] = 12'haaa;
rom[114993] = 12'haaa;
rom[114994] = 12'haaa;
rom[114995] = 12'haaa;
rom[114996] = 12'haaa;
rom[114997] = 12'haaa;
rom[114998] = 12'h999;
rom[114999] = 12'h999;
rom[115000] = 12'h999;
rom[115001] = 12'h999;
rom[115002] = 12'h999;
rom[115003] = 12'h999;
rom[115004] = 12'h888;
rom[115005] = 12'h888;
rom[115006] = 12'h888;
rom[115007] = 12'h888;
rom[115008] = 12'h888;
rom[115009] = 12'h888;
rom[115010] = 12'h888;
rom[115011] = 12'h888;
rom[115012] = 12'h777;
rom[115013] = 12'h777;
rom[115014] = 12'h777;
rom[115015] = 12'h777;
rom[115016] = 12'h666;
rom[115017] = 12'h555;
rom[115018] = 12'h444;
rom[115019] = 12'h444;
rom[115020] = 12'h333;
rom[115021] = 12'h333;
rom[115022] = 12'h444;
rom[115023] = 12'h777;
rom[115024] = 12'hbbb;
rom[115025] = 12'h888;
rom[115026] = 12'h444;
rom[115027] = 12'h222;
rom[115028] = 12'h222;
rom[115029] = 12'h222;
rom[115030] = 12'h111;
rom[115031] = 12'h  0;
rom[115032] = 12'h111;
rom[115033] = 12'h222;
rom[115034] = 12'h444;
rom[115035] = 12'h333;
rom[115036] = 12'h222;
rom[115037] = 12'h111;
rom[115038] = 12'h111;
rom[115039] = 12'h222;
rom[115040] = 12'h333;
rom[115041] = 12'h666;
rom[115042] = 12'hbbb;
rom[115043] = 12'hccc;
rom[115044] = 12'h888;
rom[115045] = 12'h333;
rom[115046] = 12'h111;
rom[115047] = 12'h111;
rom[115048] = 12'h111;
rom[115049] = 12'h  0;
rom[115050] = 12'h  0;
rom[115051] = 12'h  0;
rom[115052] = 12'h  0;
rom[115053] = 12'h  0;
rom[115054] = 12'h  0;
rom[115055] = 12'h  0;
rom[115056] = 12'h  0;
rom[115057] = 12'h  0;
rom[115058] = 12'h  0;
rom[115059] = 12'h111;
rom[115060] = 12'h111;
rom[115061] = 12'h111;
rom[115062] = 12'h111;
rom[115063] = 12'h444;
rom[115064] = 12'hccc;
rom[115065] = 12'heee;
rom[115066] = 12'hbbb;
rom[115067] = 12'h666;
rom[115068] = 12'h333;
rom[115069] = 12'h222;
rom[115070] = 12'h111;
rom[115071] = 12'h111;
rom[115072] = 12'h111;
rom[115073] = 12'h111;
rom[115074] = 12'h333;
rom[115075] = 12'h888;
rom[115076] = 12'heee;
rom[115077] = 12'haaa;
rom[115078] = 12'h444;
rom[115079] = 12'h  0;
rom[115080] = 12'h  0;
rom[115081] = 12'h111;
rom[115082] = 12'h  0;
rom[115083] = 12'h  0;
rom[115084] = 12'h  0;
rom[115085] = 12'h111;
rom[115086] = 12'h  0;
rom[115087] = 12'h  0;
rom[115088] = 12'h111;
rom[115089] = 12'h444;
rom[115090] = 12'h888;
rom[115091] = 12'h888;
rom[115092] = 12'h555;
rom[115093] = 12'haaa;
rom[115094] = 12'hbbb;
rom[115095] = 12'h666;
rom[115096] = 12'h111;
rom[115097] = 12'h111;
rom[115098] = 12'h111;
rom[115099] = 12'h111;
rom[115100] = 12'h111;
rom[115101] = 12'h  0;
rom[115102] = 12'h111;
rom[115103] = 12'h111;
rom[115104] = 12'h111;
rom[115105] = 12'h111;
rom[115106] = 12'h111;
rom[115107] = 12'h222;
rom[115108] = 12'h111;
rom[115109] = 12'h111;
rom[115110] = 12'h333;
rom[115111] = 12'h555;
rom[115112] = 12'h777;
rom[115113] = 12'h888;
rom[115114] = 12'haaa;
rom[115115] = 12'hccc;
rom[115116] = 12'haaa;
rom[115117] = 12'h666;
rom[115118] = 12'h333;
rom[115119] = 12'h222;
rom[115120] = 12'h222;
rom[115121] = 12'h222;
rom[115122] = 12'h111;
rom[115123] = 12'h111;
rom[115124] = 12'h  0;
rom[115125] = 12'h  0;
rom[115126] = 12'h  0;
rom[115127] = 12'h  0;
rom[115128] = 12'h  0;
rom[115129] = 12'h  0;
rom[115130] = 12'h  0;
rom[115131] = 12'h  0;
rom[115132] = 12'h  0;
rom[115133] = 12'h  0;
rom[115134] = 12'h  0;
rom[115135] = 12'h  0;
rom[115136] = 12'h  0;
rom[115137] = 12'h  0;
rom[115138] = 12'h  0;
rom[115139] = 12'h  0;
rom[115140] = 12'h  0;
rom[115141] = 12'h  0;
rom[115142] = 12'h  0;
rom[115143] = 12'h  0;
rom[115144] = 12'h  0;
rom[115145] = 12'h  0;
rom[115146] = 12'h  0;
rom[115147] = 12'h  0;
rom[115148] = 12'h  0;
rom[115149] = 12'h  0;
rom[115150] = 12'h  0;
rom[115151] = 12'h  0;
rom[115152] = 12'h  0;
rom[115153] = 12'h  0;
rom[115154] = 12'h  0;
rom[115155] = 12'h  0;
rom[115156] = 12'h  0;
rom[115157] = 12'h  0;
rom[115158] = 12'h  0;
rom[115159] = 12'h  0;
rom[115160] = 12'h  0;
rom[115161] = 12'h  0;
rom[115162] = 12'h  0;
rom[115163] = 12'h  0;
rom[115164] = 12'h  0;
rom[115165] = 12'h  0;
rom[115166] = 12'h111;
rom[115167] = 12'h111;
rom[115168] = 12'h555;
rom[115169] = 12'h888;
rom[115170] = 12'hbbb;
rom[115171] = 12'haaa;
rom[115172] = 12'h777;
rom[115173] = 12'h444;
rom[115174] = 12'h222;
rom[115175] = 12'h222;
rom[115176] = 12'h111;
rom[115177] = 12'h111;
rom[115178] = 12'h  0;
rom[115179] = 12'h  0;
rom[115180] = 12'h  0;
rom[115181] = 12'h  0;
rom[115182] = 12'h  0;
rom[115183] = 12'h  0;
rom[115184] = 12'h  0;
rom[115185] = 12'h  0;
rom[115186] = 12'h  0;
rom[115187] = 12'h  0;
rom[115188] = 12'h  0;
rom[115189] = 12'h  0;
rom[115190] = 12'h  0;
rom[115191] = 12'h  0;
rom[115192] = 12'h  0;
rom[115193] = 12'h  0;
rom[115194] = 12'h  0;
rom[115195] = 12'h  0;
rom[115196] = 12'h  0;
rom[115197] = 12'h  0;
rom[115198] = 12'h  0;
rom[115199] = 12'h  0;
rom[115200] = 12'hfff;
rom[115201] = 12'hfff;
rom[115202] = 12'hfff;
rom[115203] = 12'hfff;
rom[115204] = 12'hfff;
rom[115205] = 12'hfff;
rom[115206] = 12'hfff;
rom[115207] = 12'hfff;
rom[115208] = 12'hfff;
rom[115209] = 12'hfff;
rom[115210] = 12'hfff;
rom[115211] = 12'hfff;
rom[115212] = 12'hfff;
rom[115213] = 12'hfff;
rom[115214] = 12'hfff;
rom[115215] = 12'hfff;
rom[115216] = 12'hfff;
rom[115217] = 12'hfff;
rom[115218] = 12'hfff;
rom[115219] = 12'heee;
rom[115220] = 12'heee;
rom[115221] = 12'heee;
rom[115222] = 12'heee;
rom[115223] = 12'heee;
rom[115224] = 12'heee;
rom[115225] = 12'heee;
rom[115226] = 12'heee;
rom[115227] = 12'heee;
rom[115228] = 12'heee;
rom[115229] = 12'heee;
rom[115230] = 12'heee;
rom[115231] = 12'heee;
rom[115232] = 12'heee;
rom[115233] = 12'heee;
rom[115234] = 12'heee;
rom[115235] = 12'heee;
rom[115236] = 12'heee;
rom[115237] = 12'heee;
rom[115238] = 12'heee;
rom[115239] = 12'heee;
rom[115240] = 12'heee;
rom[115241] = 12'hddd;
rom[115242] = 12'hddd;
rom[115243] = 12'hddd;
rom[115244] = 12'hddd;
rom[115245] = 12'hddd;
rom[115246] = 12'hddd;
rom[115247] = 12'hddd;
rom[115248] = 12'hddd;
rom[115249] = 12'hddd;
rom[115250] = 12'hddd;
rom[115251] = 12'hddd;
rom[115252] = 12'hddd;
rom[115253] = 12'hccc;
rom[115254] = 12'hccc;
rom[115255] = 12'hccc;
rom[115256] = 12'hccc;
rom[115257] = 12'hccc;
rom[115258] = 12'hccc;
rom[115259] = 12'hccc;
rom[115260] = 12'hccc;
rom[115261] = 12'hccc;
rom[115262] = 12'hccc;
rom[115263] = 12'hccc;
rom[115264] = 12'hbbb;
rom[115265] = 12'hbbb;
rom[115266] = 12'hbbb;
rom[115267] = 12'hbbb;
rom[115268] = 12'hbbb;
rom[115269] = 12'hbbb;
rom[115270] = 12'hbbb;
rom[115271] = 12'hbbb;
rom[115272] = 12'hbbb;
rom[115273] = 12'hbbb;
rom[115274] = 12'hbbb;
rom[115275] = 12'hbbb;
rom[115276] = 12'hbbb;
rom[115277] = 12'hccc;
rom[115278] = 12'hddd;
rom[115279] = 12'heee;
rom[115280] = 12'hfff;
rom[115281] = 12'hfff;
rom[115282] = 12'hfff;
rom[115283] = 12'hddd;
rom[115284] = 12'hbbb;
rom[115285] = 12'hbbb;
rom[115286] = 12'hbbb;
rom[115287] = 12'haaa;
rom[115288] = 12'haaa;
rom[115289] = 12'haaa;
rom[115290] = 12'haaa;
rom[115291] = 12'haaa;
rom[115292] = 12'h999;
rom[115293] = 12'haaa;
rom[115294] = 12'haaa;
rom[115295] = 12'h999;
rom[115296] = 12'h999;
rom[115297] = 12'haaa;
rom[115298] = 12'haaa;
rom[115299] = 12'hccc;
rom[115300] = 12'hccc;
rom[115301] = 12'haaa;
rom[115302] = 12'h999;
rom[115303] = 12'hbbb;
rom[115304] = 12'haaa;
rom[115305] = 12'h999;
rom[115306] = 12'h888;
rom[115307] = 12'h888;
rom[115308] = 12'h888;
rom[115309] = 12'h777;
rom[115310] = 12'h777;
rom[115311] = 12'h777;
rom[115312] = 12'h777;
rom[115313] = 12'h777;
rom[115314] = 12'h777;
rom[115315] = 12'h666;
rom[115316] = 12'h777;
rom[115317] = 12'h777;
rom[115318] = 12'h777;
rom[115319] = 12'h777;
rom[115320] = 12'h888;
rom[115321] = 12'h888;
rom[115322] = 12'h777;
rom[115323] = 12'h777;
rom[115324] = 12'h666;
rom[115325] = 12'h666;
rom[115326] = 12'h555;
rom[115327] = 12'h555;
rom[115328] = 12'h555;
rom[115329] = 12'h666;
rom[115330] = 12'h777;
rom[115331] = 12'h666;
rom[115332] = 12'h555;
rom[115333] = 12'h555;
rom[115334] = 12'h555;
rom[115335] = 12'h555;
rom[115336] = 12'h555;
rom[115337] = 12'h666;
rom[115338] = 12'h666;
rom[115339] = 12'h666;
rom[115340] = 12'h555;
rom[115341] = 12'h444;
rom[115342] = 12'h444;
rom[115343] = 12'h444;
rom[115344] = 12'h444;
rom[115345] = 12'h444;
rom[115346] = 12'h444;
rom[115347] = 12'h444;
rom[115348] = 12'h444;
rom[115349] = 12'h444;
rom[115350] = 12'h444;
rom[115351] = 12'h444;
rom[115352] = 12'h555;
rom[115353] = 12'h555;
rom[115354] = 12'h555;
rom[115355] = 12'h555;
rom[115356] = 12'h555;
rom[115357] = 12'h666;
rom[115358] = 12'h666;
rom[115359] = 12'h666;
rom[115360] = 12'h777;
rom[115361] = 12'h777;
rom[115362] = 12'h777;
rom[115363] = 12'h777;
rom[115364] = 12'h777;
rom[115365] = 12'h777;
rom[115366] = 12'h666;
rom[115367] = 12'h666;
rom[115368] = 12'h777;
rom[115369] = 12'h777;
rom[115370] = 12'h777;
rom[115371] = 12'h777;
rom[115372] = 12'h888;
rom[115373] = 12'h888;
rom[115374] = 12'h888;
rom[115375] = 12'h888;
rom[115376] = 12'h888;
rom[115377] = 12'h888;
rom[115378] = 12'h888;
rom[115379] = 12'h888;
rom[115380] = 12'h888;
rom[115381] = 12'h888;
rom[115382] = 12'h888;
rom[115383] = 12'h888;
rom[115384] = 12'h888;
rom[115385] = 12'h888;
rom[115386] = 12'h999;
rom[115387] = 12'h999;
rom[115388] = 12'h888;
rom[115389] = 12'h888;
rom[115390] = 12'h999;
rom[115391] = 12'h999;
rom[115392] = 12'h888;
rom[115393] = 12'h888;
rom[115394] = 12'h888;
rom[115395] = 12'h888;
rom[115396] = 12'h888;
rom[115397] = 12'h888;
rom[115398] = 12'h999;
rom[115399] = 12'h999;
rom[115400] = 12'h999;
rom[115401] = 12'h888;
rom[115402] = 12'h777;
rom[115403] = 12'h777;
rom[115404] = 12'h777;
rom[115405] = 12'h777;
rom[115406] = 12'h777;
rom[115407] = 12'h777;
rom[115408] = 12'h777;
rom[115409] = 12'h777;
rom[115410] = 12'h777;
rom[115411] = 12'h777;
rom[115412] = 12'h777;
rom[115413] = 12'h666;
rom[115414] = 12'h666;
rom[115415] = 12'h666;
rom[115416] = 12'h666;
rom[115417] = 12'h555;
rom[115418] = 12'h444;
rom[115419] = 12'h333;
rom[115420] = 12'h333;
rom[115421] = 12'h333;
rom[115422] = 12'h333;
rom[115423] = 12'h333;
rom[115424] = 12'h777;
rom[115425] = 12'haaa;
rom[115426] = 12'h888;
rom[115427] = 12'h333;
rom[115428] = 12'h111;
rom[115429] = 12'h111;
rom[115430] = 12'h111;
rom[115431] = 12'h111;
rom[115432] = 12'h  0;
rom[115433] = 12'h111;
rom[115434] = 12'h333;
rom[115435] = 12'h333;
rom[115436] = 12'h222;
rom[115437] = 12'h111;
rom[115438] = 12'h222;
rom[115439] = 12'h111;
rom[115440] = 12'h444;
rom[115441] = 12'h999;
rom[115442] = 12'hddd;
rom[115443] = 12'haaa;
rom[115444] = 12'h444;
rom[115445] = 12'h111;
rom[115446] = 12'h111;
rom[115447] = 12'h  0;
rom[115448] = 12'h  0;
rom[115449] = 12'h  0;
rom[115450] = 12'h  0;
rom[115451] = 12'h  0;
rom[115452] = 12'h  0;
rom[115453] = 12'h  0;
rom[115454] = 12'h  0;
rom[115455] = 12'h  0;
rom[115456] = 12'h  0;
rom[115457] = 12'h  0;
rom[115458] = 12'h111;
rom[115459] = 12'h  0;
rom[115460] = 12'h  0;
rom[115461] = 12'h111;
rom[115462] = 12'h111;
rom[115463] = 12'h444;
rom[115464] = 12'hbbb;
rom[115465] = 12'heee;
rom[115466] = 12'hccc;
rom[115467] = 12'h666;
rom[115468] = 12'h333;
rom[115469] = 12'h222;
rom[115470] = 12'h111;
rom[115471] = 12'h111;
rom[115472] = 12'h111;
rom[115473] = 12'h  0;
rom[115474] = 12'h222;
rom[115475] = 12'h666;
rom[115476] = 12'hddd;
rom[115477] = 12'hbbb;
rom[115478] = 12'h666;
rom[115479] = 12'h  0;
rom[115480] = 12'h  0;
rom[115481] = 12'h  0;
rom[115482] = 12'h  0;
rom[115483] = 12'h  0;
rom[115484] = 12'h  0;
rom[115485] = 12'h  0;
rom[115486] = 12'h111;
rom[115487] = 12'h  0;
rom[115488] = 12'h111;
rom[115489] = 12'h333;
rom[115490] = 12'h666;
rom[115491] = 12'h888;
rom[115492] = 12'h666;
rom[115493] = 12'h666;
rom[115494] = 12'h999;
rom[115495] = 12'haaa;
rom[115496] = 12'h444;
rom[115497] = 12'h111;
rom[115498] = 12'h  0;
rom[115499] = 12'h111;
rom[115500] = 12'h  0;
rom[115501] = 12'h  0;
rom[115502] = 12'h111;
rom[115503] = 12'h111;
rom[115504] = 12'h111;
rom[115505] = 12'h111;
rom[115506] = 12'h111;
rom[115507] = 12'h111;
rom[115508] = 12'h111;
rom[115509] = 12'h222;
rom[115510] = 12'h222;
rom[115511] = 12'h333;
rom[115512] = 12'h555;
rom[115513] = 12'h777;
rom[115514] = 12'h999;
rom[115515] = 12'haaa;
rom[115516] = 12'haaa;
rom[115517] = 12'h999;
rom[115518] = 12'h555;
rom[115519] = 12'h222;
rom[115520] = 12'h222;
rom[115521] = 12'h111;
rom[115522] = 12'h111;
rom[115523] = 12'h111;
rom[115524] = 12'h111;
rom[115525] = 12'h  0;
rom[115526] = 12'h  0;
rom[115527] = 12'h  0;
rom[115528] = 12'h  0;
rom[115529] = 12'h  0;
rom[115530] = 12'h  0;
rom[115531] = 12'h  0;
rom[115532] = 12'h  0;
rom[115533] = 12'h  0;
rom[115534] = 12'h  0;
rom[115535] = 12'h  0;
rom[115536] = 12'h  0;
rom[115537] = 12'h  0;
rom[115538] = 12'h  0;
rom[115539] = 12'h  0;
rom[115540] = 12'h  0;
rom[115541] = 12'h  0;
rom[115542] = 12'h  0;
rom[115543] = 12'h  0;
rom[115544] = 12'h  0;
rom[115545] = 12'h  0;
rom[115546] = 12'h  0;
rom[115547] = 12'h  0;
rom[115548] = 12'h  0;
rom[115549] = 12'h  0;
rom[115550] = 12'h  0;
rom[115551] = 12'h  0;
rom[115552] = 12'h  0;
rom[115553] = 12'h  0;
rom[115554] = 12'h  0;
rom[115555] = 12'h  0;
rom[115556] = 12'h  0;
rom[115557] = 12'h  0;
rom[115558] = 12'h  0;
rom[115559] = 12'h  0;
rom[115560] = 12'h  0;
rom[115561] = 12'h  0;
rom[115562] = 12'h  0;
rom[115563] = 12'h  0;
rom[115564] = 12'h  0;
rom[115565] = 12'h  0;
rom[115566] = 12'h111;
rom[115567] = 12'h111;
rom[115568] = 12'h333;
rom[115569] = 12'h666;
rom[115570] = 12'haaa;
rom[115571] = 12'hbbb;
rom[115572] = 12'haaa;
rom[115573] = 12'h666;
rom[115574] = 12'h333;
rom[115575] = 12'h111;
rom[115576] = 12'h111;
rom[115577] = 12'h111;
rom[115578] = 12'h  0;
rom[115579] = 12'h  0;
rom[115580] = 12'h  0;
rom[115581] = 12'h  0;
rom[115582] = 12'h  0;
rom[115583] = 12'h  0;
rom[115584] = 12'h  0;
rom[115585] = 12'h  0;
rom[115586] = 12'h  0;
rom[115587] = 12'h  0;
rom[115588] = 12'h  0;
rom[115589] = 12'h  0;
rom[115590] = 12'h  0;
rom[115591] = 12'h  0;
rom[115592] = 12'h  0;
rom[115593] = 12'h  0;
rom[115594] = 12'h  0;
rom[115595] = 12'h  0;
rom[115596] = 12'h  0;
rom[115597] = 12'h  0;
rom[115598] = 12'h  0;
rom[115599] = 12'h  0;
rom[115600] = 12'hfff;
rom[115601] = 12'hfff;
rom[115602] = 12'hfff;
rom[115603] = 12'hfff;
rom[115604] = 12'hfff;
rom[115605] = 12'hfff;
rom[115606] = 12'hfff;
rom[115607] = 12'hfff;
rom[115608] = 12'hfff;
rom[115609] = 12'hfff;
rom[115610] = 12'hfff;
rom[115611] = 12'hfff;
rom[115612] = 12'hfff;
rom[115613] = 12'hfff;
rom[115614] = 12'hfff;
rom[115615] = 12'hfff;
rom[115616] = 12'hfff;
rom[115617] = 12'hfff;
rom[115618] = 12'hfff;
rom[115619] = 12'heee;
rom[115620] = 12'heee;
rom[115621] = 12'heee;
rom[115622] = 12'heee;
rom[115623] = 12'heee;
rom[115624] = 12'heee;
rom[115625] = 12'heee;
rom[115626] = 12'heee;
rom[115627] = 12'heee;
rom[115628] = 12'heee;
rom[115629] = 12'heee;
rom[115630] = 12'heee;
rom[115631] = 12'heee;
rom[115632] = 12'heee;
rom[115633] = 12'heee;
rom[115634] = 12'heee;
rom[115635] = 12'heee;
rom[115636] = 12'heee;
rom[115637] = 12'heee;
rom[115638] = 12'heee;
rom[115639] = 12'heee;
rom[115640] = 12'heee;
rom[115641] = 12'hddd;
rom[115642] = 12'hddd;
rom[115643] = 12'hddd;
rom[115644] = 12'hddd;
rom[115645] = 12'hddd;
rom[115646] = 12'hddd;
rom[115647] = 12'hddd;
rom[115648] = 12'hddd;
rom[115649] = 12'hddd;
rom[115650] = 12'hddd;
rom[115651] = 12'hddd;
rom[115652] = 12'hddd;
rom[115653] = 12'hccc;
rom[115654] = 12'hccc;
rom[115655] = 12'hccc;
rom[115656] = 12'hccc;
rom[115657] = 12'hccc;
rom[115658] = 12'hccc;
rom[115659] = 12'hccc;
rom[115660] = 12'hccc;
rom[115661] = 12'hccc;
rom[115662] = 12'hccc;
rom[115663] = 12'hccc;
rom[115664] = 12'hbbb;
rom[115665] = 12'hbbb;
rom[115666] = 12'hbbb;
rom[115667] = 12'hbbb;
rom[115668] = 12'hbbb;
rom[115669] = 12'hbbb;
rom[115670] = 12'hbbb;
rom[115671] = 12'hbbb;
rom[115672] = 12'hbbb;
rom[115673] = 12'hbbb;
rom[115674] = 12'hbbb;
rom[115675] = 12'hbbb;
rom[115676] = 12'hccc;
rom[115677] = 12'hddd;
rom[115678] = 12'heee;
rom[115679] = 12'hfff;
rom[115680] = 12'hfff;
rom[115681] = 12'hfff;
rom[115682] = 12'heee;
rom[115683] = 12'hccc;
rom[115684] = 12'hbbb;
rom[115685] = 12'haaa;
rom[115686] = 12'haaa;
rom[115687] = 12'haaa;
rom[115688] = 12'haaa;
rom[115689] = 12'haaa;
rom[115690] = 12'haaa;
rom[115691] = 12'haaa;
rom[115692] = 12'haaa;
rom[115693] = 12'haaa;
rom[115694] = 12'h999;
rom[115695] = 12'h999;
rom[115696] = 12'h999;
rom[115697] = 12'haaa;
rom[115698] = 12'hbbb;
rom[115699] = 12'hccc;
rom[115700] = 12'hbbb;
rom[115701] = 12'h999;
rom[115702] = 12'h999;
rom[115703] = 12'hbbb;
rom[115704] = 12'haaa;
rom[115705] = 12'h888;
rom[115706] = 12'h777;
rom[115707] = 12'h888;
rom[115708] = 12'h888;
rom[115709] = 12'h777;
rom[115710] = 12'h777;
rom[115711] = 12'h777;
rom[115712] = 12'h666;
rom[115713] = 12'h666;
rom[115714] = 12'h666;
rom[115715] = 12'h666;
rom[115716] = 12'h666;
rom[115717] = 12'h666;
rom[115718] = 12'h777;
rom[115719] = 12'h777;
rom[115720] = 12'h777;
rom[115721] = 12'h777;
rom[115722] = 12'h777;
rom[115723] = 12'h777;
rom[115724] = 12'h666;
rom[115725] = 12'h555;
rom[115726] = 12'h555;
rom[115727] = 12'h555;
rom[115728] = 12'h666;
rom[115729] = 12'h666;
rom[115730] = 12'h777;
rom[115731] = 12'h666;
rom[115732] = 12'h555;
rom[115733] = 12'h555;
rom[115734] = 12'h555;
rom[115735] = 12'h555;
rom[115736] = 12'h555;
rom[115737] = 12'h666;
rom[115738] = 12'h666;
rom[115739] = 12'h666;
rom[115740] = 12'h555;
rom[115741] = 12'h444;
rom[115742] = 12'h444;
rom[115743] = 12'h444;
rom[115744] = 12'h444;
rom[115745] = 12'h444;
rom[115746] = 12'h444;
rom[115747] = 12'h444;
rom[115748] = 12'h444;
rom[115749] = 12'h444;
rom[115750] = 12'h444;
rom[115751] = 12'h444;
rom[115752] = 12'h444;
rom[115753] = 12'h444;
rom[115754] = 12'h444;
rom[115755] = 12'h555;
rom[115756] = 12'h555;
rom[115757] = 12'h555;
rom[115758] = 12'h666;
rom[115759] = 12'h666;
rom[115760] = 12'h777;
rom[115761] = 12'h777;
rom[115762] = 12'h777;
rom[115763] = 12'h666;
rom[115764] = 12'h666;
rom[115765] = 12'h666;
rom[115766] = 12'h666;
rom[115767] = 12'h666;
rom[115768] = 12'h666;
rom[115769] = 12'h666;
rom[115770] = 12'h666;
rom[115771] = 12'h777;
rom[115772] = 12'h777;
rom[115773] = 12'h777;
rom[115774] = 12'h777;
rom[115775] = 12'h777;
rom[115776] = 12'h777;
rom[115777] = 12'h888;
rom[115778] = 12'h888;
rom[115779] = 12'h777;
rom[115780] = 12'h777;
rom[115781] = 12'h777;
rom[115782] = 12'h888;
rom[115783] = 12'h777;
rom[115784] = 12'h777;
rom[115785] = 12'h888;
rom[115786] = 12'h888;
rom[115787] = 12'h777;
rom[115788] = 12'h777;
rom[115789] = 12'h888;
rom[115790] = 12'h888;
rom[115791] = 12'h888;
rom[115792] = 12'h888;
rom[115793] = 12'h777;
rom[115794] = 12'h777;
rom[115795] = 12'h888;
rom[115796] = 12'h888;
rom[115797] = 12'h888;
rom[115798] = 12'h888;
rom[115799] = 12'h888;
rom[115800] = 12'h888;
rom[115801] = 12'h777;
rom[115802] = 12'h777;
rom[115803] = 12'h777;
rom[115804] = 12'h777;
rom[115805] = 12'h666;
rom[115806] = 12'h666;
rom[115807] = 12'h666;
rom[115808] = 12'h666;
rom[115809] = 12'h666;
rom[115810] = 12'h666;
rom[115811] = 12'h777;
rom[115812] = 12'h777;
rom[115813] = 12'h666;
rom[115814] = 12'h555;
rom[115815] = 12'h555;
rom[115816] = 12'h666;
rom[115817] = 12'h555;
rom[115818] = 12'h444;
rom[115819] = 12'h333;
rom[115820] = 12'h222;
rom[115821] = 12'h333;
rom[115822] = 12'h333;
rom[115823] = 12'h333;
rom[115824] = 12'h555;
rom[115825] = 12'h888;
rom[115826] = 12'h999;
rom[115827] = 12'h555;
rom[115828] = 12'h111;
rom[115829] = 12'h111;
rom[115830] = 12'h111;
rom[115831] = 12'h111;
rom[115832] = 12'h  0;
rom[115833] = 12'h111;
rom[115834] = 12'h333;
rom[115835] = 12'h333;
rom[115836] = 12'h222;
rom[115837] = 12'h222;
rom[115838] = 12'h222;
rom[115839] = 12'h222;
rom[115840] = 12'h666;
rom[115841] = 12'haaa;
rom[115842] = 12'hccc;
rom[115843] = 12'h888;
rom[115844] = 12'h333;
rom[115845] = 12'h  0;
rom[115846] = 12'h  0;
rom[115847] = 12'h  0;
rom[115848] = 12'h  0;
rom[115849] = 12'h  0;
rom[115850] = 12'h  0;
rom[115851] = 12'h  0;
rom[115852] = 12'h  0;
rom[115853] = 12'h  0;
rom[115854] = 12'h  0;
rom[115855] = 12'h  0;
rom[115856] = 12'h  0;
rom[115857] = 12'h  0;
rom[115858] = 12'h  0;
rom[115859] = 12'h  0;
rom[115860] = 12'h  0;
rom[115861] = 12'h111;
rom[115862] = 12'h111;
rom[115863] = 12'h444;
rom[115864] = 12'hbbb;
rom[115865] = 12'heee;
rom[115866] = 12'hccc;
rom[115867] = 12'h666;
rom[115868] = 12'h333;
rom[115869] = 12'h222;
rom[115870] = 12'h111;
rom[115871] = 12'h111;
rom[115872] = 12'h111;
rom[115873] = 12'h  0;
rom[115874] = 12'h222;
rom[115875] = 12'h555;
rom[115876] = 12'hbbb;
rom[115877] = 12'hccc;
rom[115878] = 12'h777;
rom[115879] = 12'h111;
rom[115880] = 12'h111;
rom[115881] = 12'h  0;
rom[115882] = 12'h  0;
rom[115883] = 12'h  0;
rom[115884] = 12'h  0;
rom[115885] = 12'h  0;
rom[115886] = 12'h  0;
rom[115887] = 12'h  0;
rom[115888] = 12'h  0;
rom[115889] = 12'h222;
rom[115890] = 12'h666;
rom[115891] = 12'h888;
rom[115892] = 12'h666;
rom[115893] = 12'h555;
rom[115894] = 12'h888;
rom[115895] = 12'haaa;
rom[115896] = 12'h555;
rom[115897] = 12'h222;
rom[115898] = 12'h  0;
rom[115899] = 12'h111;
rom[115900] = 12'h111;
rom[115901] = 12'h111;
rom[115902] = 12'h111;
rom[115903] = 12'h111;
rom[115904] = 12'h111;
rom[115905] = 12'h111;
rom[115906] = 12'h111;
rom[115907] = 12'h111;
rom[115908] = 12'h111;
rom[115909] = 12'h222;
rom[115910] = 12'h222;
rom[115911] = 12'h222;
rom[115912] = 12'h444;
rom[115913] = 12'h666;
rom[115914] = 12'h888;
rom[115915] = 12'haaa;
rom[115916] = 12'haaa;
rom[115917] = 12'h999;
rom[115918] = 12'h666;
rom[115919] = 12'h333;
rom[115920] = 12'h222;
rom[115921] = 12'h111;
rom[115922] = 12'h111;
rom[115923] = 12'h111;
rom[115924] = 12'h111;
rom[115925] = 12'h  0;
rom[115926] = 12'h  0;
rom[115927] = 12'h  0;
rom[115928] = 12'h  0;
rom[115929] = 12'h  0;
rom[115930] = 12'h  0;
rom[115931] = 12'h  0;
rom[115932] = 12'h  0;
rom[115933] = 12'h  0;
rom[115934] = 12'h  0;
rom[115935] = 12'h  0;
rom[115936] = 12'h  0;
rom[115937] = 12'h  0;
rom[115938] = 12'h  0;
rom[115939] = 12'h  0;
rom[115940] = 12'h  0;
rom[115941] = 12'h  0;
rom[115942] = 12'h  0;
rom[115943] = 12'h  0;
rom[115944] = 12'h  0;
rom[115945] = 12'h  0;
rom[115946] = 12'h  0;
rom[115947] = 12'h  0;
rom[115948] = 12'h  0;
rom[115949] = 12'h  0;
rom[115950] = 12'h  0;
rom[115951] = 12'h  0;
rom[115952] = 12'h  0;
rom[115953] = 12'h  0;
rom[115954] = 12'h  0;
rom[115955] = 12'h  0;
rom[115956] = 12'h  0;
rom[115957] = 12'h  0;
rom[115958] = 12'h  0;
rom[115959] = 12'h  0;
rom[115960] = 12'h  0;
rom[115961] = 12'h  0;
rom[115962] = 12'h  0;
rom[115963] = 12'h  0;
rom[115964] = 12'h  0;
rom[115965] = 12'h  0;
rom[115966] = 12'h  0;
rom[115967] = 12'h111;
rom[115968] = 12'h222;
rom[115969] = 12'h444;
rom[115970] = 12'h888;
rom[115971] = 12'haaa;
rom[115972] = 12'haaa;
rom[115973] = 12'h777;
rom[115974] = 12'h444;
rom[115975] = 12'h222;
rom[115976] = 12'h111;
rom[115977] = 12'h111;
rom[115978] = 12'h  0;
rom[115979] = 12'h  0;
rom[115980] = 12'h  0;
rom[115981] = 12'h  0;
rom[115982] = 12'h  0;
rom[115983] = 12'h  0;
rom[115984] = 12'h  0;
rom[115985] = 12'h  0;
rom[115986] = 12'h  0;
rom[115987] = 12'h  0;
rom[115988] = 12'h  0;
rom[115989] = 12'h  0;
rom[115990] = 12'h  0;
rom[115991] = 12'h  0;
rom[115992] = 12'h  0;
rom[115993] = 12'h  0;
rom[115994] = 12'h  0;
rom[115995] = 12'h  0;
rom[115996] = 12'h  0;
rom[115997] = 12'h  0;
rom[115998] = 12'h  0;
rom[115999] = 12'h  0;
rom[116000] = 12'hfff;
rom[116001] = 12'hfff;
rom[116002] = 12'hfff;
rom[116003] = 12'hfff;
rom[116004] = 12'hfff;
rom[116005] = 12'hfff;
rom[116006] = 12'hfff;
rom[116007] = 12'hfff;
rom[116008] = 12'hfff;
rom[116009] = 12'hfff;
rom[116010] = 12'hfff;
rom[116011] = 12'hfff;
rom[116012] = 12'hfff;
rom[116013] = 12'hfff;
rom[116014] = 12'hfff;
rom[116015] = 12'hfff;
rom[116016] = 12'hfff;
rom[116017] = 12'hfff;
rom[116018] = 12'heee;
rom[116019] = 12'heee;
rom[116020] = 12'heee;
rom[116021] = 12'heee;
rom[116022] = 12'heee;
rom[116023] = 12'heee;
rom[116024] = 12'heee;
rom[116025] = 12'heee;
rom[116026] = 12'heee;
rom[116027] = 12'heee;
rom[116028] = 12'heee;
rom[116029] = 12'heee;
rom[116030] = 12'heee;
rom[116031] = 12'heee;
rom[116032] = 12'heee;
rom[116033] = 12'heee;
rom[116034] = 12'heee;
rom[116035] = 12'heee;
rom[116036] = 12'hddd;
rom[116037] = 12'hddd;
rom[116038] = 12'heee;
rom[116039] = 12'heee;
rom[116040] = 12'hddd;
rom[116041] = 12'hddd;
rom[116042] = 12'hddd;
rom[116043] = 12'hddd;
rom[116044] = 12'hddd;
rom[116045] = 12'hddd;
rom[116046] = 12'hddd;
rom[116047] = 12'hddd;
rom[116048] = 12'hddd;
rom[116049] = 12'hddd;
rom[116050] = 12'hddd;
rom[116051] = 12'hddd;
rom[116052] = 12'hccc;
rom[116053] = 12'hccc;
rom[116054] = 12'hccc;
rom[116055] = 12'hccc;
rom[116056] = 12'hccc;
rom[116057] = 12'hccc;
rom[116058] = 12'hccc;
rom[116059] = 12'hbbb;
rom[116060] = 12'hbbb;
rom[116061] = 12'hccc;
rom[116062] = 12'hccc;
rom[116063] = 12'hccc;
rom[116064] = 12'hbbb;
rom[116065] = 12'hbbb;
rom[116066] = 12'hbbb;
rom[116067] = 12'hbbb;
rom[116068] = 12'hbbb;
rom[116069] = 12'hbbb;
rom[116070] = 12'hbbb;
rom[116071] = 12'hbbb;
rom[116072] = 12'hbbb;
rom[116073] = 12'hbbb;
rom[116074] = 12'hbbb;
rom[116075] = 12'hbbb;
rom[116076] = 12'hccc;
rom[116077] = 12'heee;
rom[116078] = 12'hfff;
rom[116079] = 12'hfff;
rom[116080] = 12'hfff;
rom[116081] = 12'heee;
rom[116082] = 12'hccc;
rom[116083] = 12'hbbb;
rom[116084] = 12'haaa;
rom[116085] = 12'haaa;
rom[116086] = 12'haaa;
rom[116087] = 12'haaa;
rom[116088] = 12'haaa;
rom[116089] = 12'haaa;
rom[116090] = 12'haaa;
rom[116091] = 12'haaa;
rom[116092] = 12'haaa;
rom[116093] = 12'h999;
rom[116094] = 12'h999;
rom[116095] = 12'h888;
rom[116096] = 12'h999;
rom[116097] = 12'hbbb;
rom[116098] = 12'hbbb;
rom[116099] = 12'hbbb;
rom[116100] = 12'haaa;
rom[116101] = 12'h999;
rom[116102] = 12'h999;
rom[116103] = 12'hbbb;
rom[116104] = 12'h999;
rom[116105] = 12'h888;
rom[116106] = 12'h777;
rom[116107] = 12'h777;
rom[116108] = 12'h777;
rom[116109] = 12'h777;
rom[116110] = 12'h666;
rom[116111] = 12'h666;
rom[116112] = 12'h666;
rom[116113] = 12'h666;
rom[116114] = 12'h666;
rom[116115] = 12'h666;
rom[116116] = 12'h666;
rom[116117] = 12'h666;
rom[116118] = 12'h666;
rom[116119] = 12'h666;
rom[116120] = 12'h777;
rom[116121] = 12'h777;
rom[116122] = 12'h777;
rom[116123] = 12'h777;
rom[116124] = 12'h666;
rom[116125] = 12'h555;
rom[116126] = 12'h555;
rom[116127] = 12'h555;
rom[116128] = 12'h666;
rom[116129] = 12'h666;
rom[116130] = 12'h666;
rom[116131] = 12'h555;
rom[116132] = 12'h555;
rom[116133] = 12'h555;
rom[116134] = 12'h555;
rom[116135] = 12'h555;
rom[116136] = 12'h666;
rom[116137] = 12'h666;
rom[116138] = 12'h666;
rom[116139] = 12'h555;
rom[116140] = 12'h555;
rom[116141] = 12'h444;
rom[116142] = 12'h444;
rom[116143] = 12'h444;
rom[116144] = 12'h444;
rom[116145] = 12'h444;
rom[116146] = 12'h444;
rom[116147] = 12'h444;
rom[116148] = 12'h444;
rom[116149] = 12'h444;
rom[116150] = 12'h444;
rom[116151] = 12'h444;
rom[116152] = 12'h444;
rom[116153] = 12'h444;
rom[116154] = 12'h444;
rom[116155] = 12'h444;
rom[116156] = 12'h555;
rom[116157] = 12'h555;
rom[116158] = 12'h666;
rom[116159] = 12'h666;
rom[116160] = 12'h666;
rom[116161] = 12'h666;
rom[116162] = 12'h666;
rom[116163] = 12'h666;
rom[116164] = 12'h666;
rom[116165] = 12'h666;
rom[116166] = 12'h666;
rom[116167] = 12'h666;
rom[116168] = 12'h666;
rom[116169] = 12'h666;
rom[116170] = 12'h666;
rom[116171] = 12'h666;
rom[116172] = 12'h777;
rom[116173] = 12'h777;
rom[116174] = 12'h666;
rom[116175] = 12'h666;
rom[116176] = 12'h777;
rom[116177] = 12'h777;
rom[116178] = 12'h777;
rom[116179] = 12'h777;
rom[116180] = 12'h666;
rom[116181] = 12'h777;
rom[116182] = 12'h777;
rom[116183] = 12'h666;
rom[116184] = 12'h666;
rom[116185] = 12'h666;
rom[116186] = 12'h666;
rom[116187] = 12'h666;
rom[116188] = 12'h666;
rom[116189] = 12'h666;
rom[116190] = 12'h777;
rom[116191] = 12'h888;
rom[116192] = 12'h888;
rom[116193] = 12'h777;
rom[116194] = 12'h666;
rom[116195] = 12'h777;
rom[116196] = 12'h888;
rom[116197] = 12'h888;
rom[116198] = 12'h777;
rom[116199] = 12'h777;
rom[116200] = 12'h777;
rom[116201] = 12'h666;
rom[116202] = 12'h666;
rom[116203] = 12'h666;
rom[116204] = 12'h666;
rom[116205] = 12'h666;
rom[116206] = 12'h666;
rom[116207] = 12'h555;
rom[116208] = 12'h555;
rom[116209] = 12'h555;
rom[116210] = 12'h666;
rom[116211] = 12'h666;
rom[116212] = 12'h666;
rom[116213] = 12'h666;
rom[116214] = 12'h555;
rom[116215] = 12'h444;
rom[116216] = 12'h555;
rom[116217] = 12'h555;
rom[116218] = 12'h444;
rom[116219] = 12'h333;
rom[116220] = 12'h222;
rom[116221] = 12'h222;
rom[116222] = 12'h222;
rom[116223] = 12'h222;
rom[116224] = 12'h222;
rom[116225] = 12'h555;
rom[116226] = 12'h999;
rom[116227] = 12'h888;
rom[116228] = 12'h222;
rom[116229] = 12'h111;
rom[116230] = 12'h111;
rom[116231] = 12'h111;
rom[116232] = 12'h  0;
rom[116233] = 12'h111;
rom[116234] = 12'h111;
rom[116235] = 12'h222;
rom[116236] = 12'h222;
rom[116237] = 12'h222;
rom[116238] = 12'h222;
rom[116239] = 12'h333;
rom[116240] = 12'h888;
rom[116241] = 12'hbbb;
rom[116242] = 12'haaa;
rom[116243] = 12'h555;
rom[116244] = 12'h111;
rom[116245] = 12'h  0;
rom[116246] = 12'h  0;
rom[116247] = 12'h  0;
rom[116248] = 12'h  0;
rom[116249] = 12'h  0;
rom[116250] = 12'h  0;
rom[116251] = 12'h  0;
rom[116252] = 12'h  0;
rom[116253] = 12'h  0;
rom[116254] = 12'h  0;
rom[116255] = 12'h  0;
rom[116256] = 12'h  0;
rom[116257] = 12'h  0;
rom[116258] = 12'h  0;
rom[116259] = 12'h  0;
rom[116260] = 12'h  0;
rom[116261] = 12'h111;
rom[116262] = 12'h111;
rom[116263] = 12'h333;
rom[116264] = 12'haaa;
rom[116265] = 12'heee;
rom[116266] = 12'hccc;
rom[116267] = 12'h666;
rom[116268] = 12'h333;
rom[116269] = 12'h222;
rom[116270] = 12'h111;
rom[116271] = 12'h111;
rom[116272] = 12'h111;
rom[116273] = 12'h  0;
rom[116274] = 12'h111;
rom[116275] = 12'h444;
rom[116276] = 12'haaa;
rom[116277] = 12'hccc;
rom[116278] = 12'h888;
rom[116279] = 12'h222;
rom[116280] = 12'h111;
rom[116281] = 12'h  0;
rom[116282] = 12'h  0;
rom[116283] = 12'h111;
rom[116284] = 12'h  0;
rom[116285] = 12'h  0;
rom[116286] = 12'h  0;
rom[116287] = 12'h  0;
rom[116288] = 12'h  0;
rom[116289] = 12'h111;
rom[116290] = 12'h444;
rom[116291] = 12'h777;
rom[116292] = 12'h666;
rom[116293] = 12'h444;
rom[116294] = 12'h666;
rom[116295] = 12'h999;
rom[116296] = 12'h777;
rom[116297] = 12'h333;
rom[116298] = 12'h111;
rom[116299] = 12'h111;
rom[116300] = 12'h  0;
rom[116301] = 12'h111;
rom[116302] = 12'h111;
rom[116303] = 12'h111;
rom[116304] = 12'h111;
rom[116305] = 12'h111;
rom[116306] = 12'h111;
rom[116307] = 12'h111;
rom[116308] = 12'h111;
rom[116309] = 12'h111;
rom[116310] = 12'h111;
rom[116311] = 12'h111;
rom[116312] = 12'h333;
rom[116313] = 12'h555;
rom[116314] = 12'h777;
rom[116315] = 12'h999;
rom[116316] = 12'haaa;
rom[116317] = 12'haaa;
rom[116318] = 12'h777;
rom[116319] = 12'h444;
rom[116320] = 12'h222;
rom[116321] = 12'h111;
rom[116322] = 12'h111;
rom[116323] = 12'h111;
rom[116324] = 12'h111;
rom[116325] = 12'h  0;
rom[116326] = 12'h  0;
rom[116327] = 12'h  0;
rom[116328] = 12'h  0;
rom[116329] = 12'h  0;
rom[116330] = 12'h  0;
rom[116331] = 12'h  0;
rom[116332] = 12'h  0;
rom[116333] = 12'h  0;
rom[116334] = 12'h  0;
rom[116335] = 12'h  0;
rom[116336] = 12'h  0;
rom[116337] = 12'h  0;
rom[116338] = 12'h  0;
rom[116339] = 12'h  0;
rom[116340] = 12'h  0;
rom[116341] = 12'h  0;
rom[116342] = 12'h  0;
rom[116343] = 12'h  0;
rom[116344] = 12'h  0;
rom[116345] = 12'h  0;
rom[116346] = 12'h  0;
rom[116347] = 12'h  0;
rom[116348] = 12'h  0;
rom[116349] = 12'h  0;
rom[116350] = 12'h  0;
rom[116351] = 12'h  0;
rom[116352] = 12'h  0;
rom[116353] = 12'h  0;
rom[116354] = 12'h  0;
rom[116355] = 12'h  0;
rom[116356] = 12'h  0;
rom[116357] = 12'h  0;
rom[116358] = 12'h  0;
rom[116359] = 12'h  0;
rom[116360] = 12'h  0;
rom[116361] = 12'h  0;
rom[116362] = 12'h  0;
rom[116363] = 12'h  0;
rom[116364] = 12'h  0;
rom[116365] = 12'h  0;
rom[116366] = 12'h  0;
rom[116367] = 12'h  0;
rom[116368] = 12'h  0;
rom[116369] = 12'h222;
rom[116370] = 12'h555;
rom[116371] = 12'h999;
rom[116372] = 12'haaa;
rom[116373] = 12'h999;
rom[116374] = 12'h666;
rom[116375] = 12'h333;
rom[116376] = 12'h111;
rom[116377] = 12'h111;
rom[116378] = 12'h111;
rom[116379] = 12'h  0;
rom[116380] = 12'h  0;
rom[116381] = 12'h  0;
rom[116382] = 12'h  0;
rom[116383] = 12'h  0;
rom[116384] = 12'h  0;
rom[116385] = 12'h  0;
rom[116386] = 12'h  0;
rom[116387] = 12'h  0;
rom[116388] = 12'h  0;
rom[116389] = 12'h  0;
rom[116390] = 12'h  0;
rom[116391] = 12'h  0;
rom[116392] = 12'h  0;
rom[116393] = 12'h  0;
rom[116394] = 12'h  0;
rom[116395] = 12'h  0;
rom[116396] = 12'h  0;
rom[116397] = 12'h  0;
rom[116398] = 12'h  0;
rom[116399] = 12'h  0;
rom[116400] = 12'hfff;
rom[116401] = 12'hfff;
rom[116402] = 12'hfff;
rom[116403] = 12'hfff;
rom[116404] = 12'hfff;
rom[116405] = 12'hfff;
rom[116406] = 12'hfff;
rom[116407] = 12'hfff;
rom[116408] = 12'hfff;
rom[116409] = 12'hfff;
rom[116410] = 12'hfff;
rom[116411] = 12'hfff;
rom[116412] = 12'heee;
rom[116413] = 12'hfff;
rom[116414] = 12'hfff;
rom[116415] = 12'hfff;
rom[116416] = 12'hfff;
rom[116417] = 12'heee;
rom[116418] = 12'heee;
rom[116419] = 12'heee;
rom[116420] = 12'heee;
rom[116421] = 12'heee;
rom[116422] = 12'heee;
rom[116423] = 12'heee;
rom[116424] = 12'heee;
rom[116425] = 12'heee;
rom[116426] = 12'heee;
rom[116427] = 12'heee;
rom[116428] = 12'heee;
rom[116429] = 12'heee;
rom[116430] = 12'heee;
rom[116431] = 12'heee;
rom[116432] = 12'heee;
rom[116433] = 12'heee;
rom[116434] = 12'hddd;
rom[116435] = 12'hddd;
rom[116436] = 12'hddd;
rom[116437] = 12'hddd;
rom[116438] = 12'hddd;
rom[116439] = 12'hddd;
rom[116440] = 12'hddd;
rom[116441] = 12'hddd;
rom[116442] = 12'hddd;
rom[116443] = 12'hddd;
rom[116444] = 12'hddd;
rom[116445] = 12'hddd;
rom[116446] = 12'hddd;
rom[116447] = 12'hddd;
rom[116448] = 12'hddd;
rom[116449] = 12'hddd;
rom[116450] = 12'hddd;
rom[116451] = 12'hddd;
rom[116452] = 12'hccc;
rom[116453] = 12'hccc;
rom[116454] = 12'hccc;
rom[116455] = 12'hccc;
rom[116456] = 12'hccc;
rom[116457] = 12'hccc;
rom[116458] = 12'hccc;
rom[116459] = 12'hbbb;
rom[116460] = 12'hbbb;
rom[116461] = 12'hbbb;
rom[116462] = 12'hbbb;
rom[116463] = 12'hbbb;
rom[116464] = 12'hbbb;
rom[116465] = 12'hbbb;
rom[116466] = 12'hbbb;
rom[116467] = 12'hbbb;
rom[116468] = 12'hbbb;
rom[116469] = 12'hbbb;
rom[116470] = 12'hbbb;
rom[116471] = 12'hbbb;
rom[116472] = 12'hccc;
rom[116473] = 12'hbbb;
rom[116474] = 12'hbbb;
rom[116475] = 12'hccc;
rom[116476] = 12'hddd;
rom[116477] = 12'heee;
rom[116478] = 12'hfff;
rom[116479] = 12'hfff;
rom[116480] = 12'heee;
rom[116481] = 12'hddd;
rom[116482] = 12'hbbb;
rom[116483] = 12'hbbb;
rom[116484] = 12'hbbb;
rom[116485] = 12'haaa;
rom[116486] = 12'haaa;
rom[116487] = 12'haaa;
rom[116488] = 12'haaa;
rom[116489] = 12'h999;
rom[116490] = 12'h999;
rom[116491] = 12'haaa;
rom[116492] = 12'haaa;
rom[116493] = 12'h999;
rom[116494] = 12'h888;
rom[116495] = 12'h888;
rom[116496] = 12'hbbb;
rom[116497] = 12'hbbb;
rom[116498] = 12'hbbb;
rom[116499] = 12'hbbb;
rom[116500] = 12'h999;
rom[116501] = 12'h888;
rom[116502] = 12'h999;
rom[116503] = 12'haaa;
rom[116504] = 12'h999;
rom[116505] = 12'h888;
rom[116506] = 12'h777;
rom[116507] = 12'h777;
rom[116508] = 12'h777;
rom[116509] = 12'h666;
rom[116510] = 12'h666;
rom[116511] = 12'h666;
rom[116512] = 12'h666;
rom[116513] = 12'h666;
rom[116514] = 12'h666;
rom[116515] = 12'h666;
rom[116516] = 12'h666;
rom[116517] = 12'h666;
rom[116518] = 12'h666;
rom[116519] = 12'h666;
rom[116520] = 12'h777;
rom[116521] = 12'h777;
rom[116522] = 12'h777;
rom[116523] = 12'h777;
rom[116524] = 12'h666;
rom[116525] = 12'h555;
rom[116526] = 12'h555;
rom[116527] = 12'h666;
rom[116528] = 12'h666;
rom[116529] = 12'h666;
rom[116530] = 12'h555;
rom[116531] = 12'h555;
rom[116532] = 12'h444;
rom[116533] = 12'h444;
rom[116534] = 12'h555;
rom[116535] = 12'h555;
rom[116536] = 12'h666;
rom[116537] = 12'h555;
rom[116538] = 12'h555;
rom[116539] = 12'h555;
rom[116540] = 12'h444;
rom[116541] = 12'h444;
rom[116542] = 12'h444;
rom[116543] = 12'h444;
rom[116544] = 12'h444;
rom[116545] = 12'h444;
rom[116546] = 12'h333;
rom[116547] = 12'h333;
rom[116548] = 12'h333;
rom[116549] = 12'h333;
rom[116550] = 12'h333;
rom[116551] = 12'h444;
rom[116552] = 12'h444;
rom[116553] = 12'h444;
rom[116554] = 12'h444;
rom[116555] = 12'h444;
rom[116556] = 12'h555;
rom[116557] = 12'h555;
rom[116558] = 12'h666;
rom[116559] = 12'h666;
rom[116560] = 12'h666;
rom[116561] = 12'h666;
rom[116562] = 12'h666;
rom[116563] = 12'h666;
rom[116564] = 12'h555;
rom[116565] = 12'h555;
rom[116566] = 12'h555;
rom[116567] = 12'h555;
rom[116568] = 12'h555;
rom[116569] = 12'h555;
rom[116570] = 12'h666;
rom[116571] = 12'h666;
rom[116572] = 12'h666;
rom[116573] = 12'h666;
rom[116574] = 12'h666;
rom[116575] = 12'h666;
rom[116576] = 12'h666;
rom[116577] = 12'h666;
rom[116578] = 12'h666;
rom[116579] = 12'h666;
rom[116580] = 12'h666;
rom[116581] = 12'h666;
rom[116582] = 12'h666;
rom[116583] = 12'h666;
rom[116584] = 12'h555;
rom[116585] = 12'h555;
rom[116586] = 12'h555;
rom[116587] = 12'h555;
rom[116588] = 12'h555;
rom[116589] = 12'h666;
rom[116590] = 12'h777;
rom[116591] = 12'h888;
rom[116592] = 12'h888;
rom[116593] = 12'h777;
rom[116594] = 12'h666;
rom[116595] = 12'h666;
rom[116596] = 12'h777;
rom[116597] = 12'h777;
rom[116598] = 12'h777;
rom[116599] = 12'h666;
rom[116600] = 12'h666;
rom[116601] = 12'h666;
rom[116602] = 12'h555;
rom[116603] = 12'h666;
rom[116604] = 12'h666;
rom[116605] = 12'h666;
rom[116606] = 12'h555;
rom[116607] = 12'h555;
rom[116608] = 12'h444;
rom[116609] = 12'h444;
rom[116610] = 12'h555;
rom[116611] = 12'h666;
rom[116612] = 12'h666;
rom[116613] = 12'h555;
rom[116614] = 12'h444;
rom[116615] = 12'h444;
rom[116616] = 12'h555;
rom[116617] = 12'h555;
rom[116618] = 12'h444;
rom[116619] = 12'h333;
rom[116620] = 12'h222;
rom[116621] = 12'h111;
rom[116622] = 12'h111;
rom[116623] = 12'h222;
rom[116624] = 12'h111;
rom[116625] = 12'h222;
rom[116626] = 12'h666;
rom[116627] = 12'h888;
rom[116628] = 12'h555;
rom[116629] = 12'h222;
rom[116630] = 12'h111;
rom[116631] = 12'h  0;
rom[116632] = 12'h  0;
rom[116633] = 12'h111;
rom[116634] = 12'h111;
rom[116635] = 12'h222;
rom[116636] = 12'h333;
rom[116637] = 12'h222;
rom[116638] = 12'h222;
rom[116639] = 12'h555;
rom[116640] = 12'h999;
rom[116641] = 12'hbbb;
rom[116642] = 12'h777;
rom[116643] = 12'h222;
rom[116644] = 12'h  0;
rom[116645] = 12'h  0;
rom[116646] = 12'h  0;
rom[116647] = 12'h  0;
rom[116648] = 12'h  0;
rom[116649] = 12'h  0;
rom[116650] = 12'h  0;
rom[116651] = 12'h  0;
rom[116652] = 12'h  0;
rom[116653] = 12'h  0;
rom[116654] = 12'h  0;
rom[116655] = 12'h  0;
rom[116656] = 12'h  0;
rom[116657] = 12'h  0;
rom[116658] = 12'h  0;
rom[116659] = 12'h  0;
rom[116660] = 12'h  0;
rom[116661] = 12'h  0;
rom[116662] = 12'h  0;
rom[116663] = 12'h333;
rom[116664] = 12'haaa;
rom[116665] = 12'heee;
rom[116666] = 12'hccc;
rom[116667] = 12'h666;
rom[116668] = 12'h333;
rom[116669] = 12'h111;
rom[116670] = 12'h  0;
rom[116671] = 12'h111;
rom[116672] = 12'h111;
rom[116673] = 12'h  0;
rom[116674] = 12'h  0;
rom[116675] = 12'h222;
rom[116676] = 12'h888;
rom[116677] = 12'hccc;
rom[116678] = 12'haaa;
rom[116679] = 12'h333;
rom[116680] = 12'h111;
rom[116681] = 12'h  0;
rom[116682] = 12'h  0;
rom[116683] = 12'h111;
rom[116684] = 12'h  0;
rom[116685] = 12'h  0;
rom[116686] = 12'h  0;
rom[116687] = 12'h  0;
rom[116688] = 12'h  0;
rom[116689] = 12'h111;
rom[116690] = 12'h333;
rom[116691] = 12'h777;
rom[116692] = 12'h666;
rom[116693] = 12'h333;
rom[116694] = 12'h444;
rom[116695] = 12'h888;
rom[116696] = 12'h888;
rom[116697] = 12'h555;
rom[116698] = 12'h222;
rom[116699] = 12'h111;
rom[116700] = 12'h  0;
rom[116701] = 12'h111;
rom[116702] = 12'h111;
rom[116703] = 12'h111;
rom[116704] = 12'h111;
rom[116705] = 12'h111;
rom[116706] = 12'h111;
rom[116707] = 12'h111;
rom[116708] = 12'h111;
rom[116709] = 12'h111;
rom[116710] = 12'h111;
rom[116711] = 12'h111;
rom[116712] = 12'h222;
rom[116713] = 12'h333;
rom[116714] = 12'h555;
rom[116715] = 12'h777;
rom[116716] = 12'h999;
rom[116717] = 12'haaa;
rom[116718] = 12'h888;
rom[116719] = 12'h666;
rom[116720] = 12'h333;
rom[116721] = 12'h222;
rom[116722] = 12'h111;
rom[116723] = 12'h111;
rom[116724] = 12'h111;
rom[116725] = 12'h  0;
rom[116726] = 12'h  0;
rom[116727] = 12'h  0;
rom[116728] = 12'h  0;
rom[116729] = 12'h  0;
rom[116730] = 12'h  0;
rom[116731] = 12'h  0;
rom[116732] = 12'h  0;
rom[116733] = 12'h  0;
rom[116734] = 12'h  0;
rom[116735] = 12'h  0;
rom[116736] = 12'h  0;
rom[116737] = 12'h  0;
rom[116738] = 12'h  0;
rom[116739] = 12'h  0;
rom[116740] = 12'h  0;
rom[116741] = 12'h  0;
rom[116742] = 12'h  0;
rom[116743] = 12'h  0;
rom[116744] = 12'h  0;
rom[116745] = 12'h  0;
rom[116746] = 12'h  0;
rom[116747] = 12'h  0;
rom[116748] = 12'h  0;
rom[116749] = 12'h  0;
rom[116750] = 12'h  0;
rom[116751] = 12'h  0;
rom[116752] = 12'h  0;
rom[116753] = 12'h  0;
rom[116754] = 12'h  0;
rom[116755] = 12'h  0;
rom[116756] = 12'h  0;
rom[116757] = 12'h  0;
rom[116758] = 12'h  0;
rom[116759] = 12'h  0;
rom[116760] = 12'h  0;
rom[116761] = 12'h  0;
rom[116762] = 12'h  0;
rom[116763] = 12'h  0;
rom[116764] = 12'h  0;
rom[116765] = 12'h  0;
rom[116766] = 12'h  0;
rom[116767] = 12'h  0;
rom[116768] = 12'h  0;
rom[116769] = 12'h111;
rom[116770] = 12'h333;
rom[116771] = 12'h666;
rom[116772] = 12'haaa;
rom[116773] = 12'haaa;
rom[116774] = 12'h777;
rom[116775] = 12'h444;
rom[116776] = 12'h222;
rom[116777] = 12'h111;
rom[116778] = 12'h  0;
rom[116779] = 12'h  0;
rom[116780] = 12'h  0;
rom[116781] = 12'h  0;
rom[116782] = 12'h  0;
rom[116783] = 12'h  0;
rom[116784] = 12'h  0;
rom[116785] = 12'h  0;
rom[116786] = 12'h  0;
rom[116787] = 12'h  0;
rom[116788] = 12'h  0;
rom[116789] = 12'h  0;
rom[116790] = 12'h  0;
rom[116791] = 12'h  0;
rom[116792] = 12'h  0;
rom[116793] = 12'h  0;
rom[116794] = 12'h  0;
rom[116795] = 12'h  0;
rom[116796] = 12'h  0;
rom[116797] = 12'h  0;
rom[116798] = 12'h  0;
rom[116799] = 12'h  0;
rom[116800] = 12'hfff;
rom[116801] = 12'hfff;
rom[116802] = 12'hfff;
rom[116803] = 12'hfff;
rom[116804] = 12'hfff;
rom[116805] = 12'hfff;
rom[116806] = 12'hfff;
rom[116807] = 12'hfff;
rom[116808] = 12'hfff;
rom[116809] = 12'heee;
rom[116810] = 12'heee;
rom[116811] = 12'heee;
rom[116812] = 12'heee;
rom[116813] = 12'heee;
rom[116814] = 12'heee;
rom[116815] = 12'heee;
rom[116816] = 12'heee;
rom[116817] = 12'heee;
rom[116818] = 12'heee;
rom[116819] = 12'heee;
rom[116820] = 12'heee;
rom[116821] = 12'heee;
rom[116822] = 12'heee;
rom[116823] = 12'heee;
rom[116824] = 12'heee;
rom[116825] = 12'heee;
rom[116826] = 12'heee;
rom[116827] = 12'heee;
rom[116828] = 12'heee;
rom[116829] = 12'heee;
rom[116830] = 12'heee;
rom[116831] = 12'heee;
rom[116832] = 12'hddd;
rom[116833] = 12'hddd;
rom[116834] = 12'hddd;
rom[116835] = 12'hddd;
rom[116836] = 12'hddd;
rom[116837] = 12'hddd;
rom[116838] = 12'hddd;
rom[116839] = 12'hddd;
rom[116840] = 12'hddd;
rom[116841] = 12'hddd;
rom[116842] = 12'hddd;
rom[116843] = 12'hddd;
rom[116844] = 12'hddd;
rom[116845] = 12'hddd;
rom[116846] = 12'hddd;
rom[116847] = 12'hccc;
rom[116848] = 12'hccc;
rom[116849] = 12'hccc;
rom[116850] = 12'hccc;
rom[116851] = 12'hccc;
rom[116852] = 12'hccc;
rom[116853] = 12'hccc;
rom[116854] = 12'hccc;
rom[116855] = 12'hccc;
rom[116856] = 12'hccc;
rom[116857] = 12'hccc;
rom[116858] = 12'hccc;
rom[116859] = 12'hbbb;
rom[116860] = 12'hbbb;
rom[116861] = 12'hbbb;
rom[116862] = 12'hbbb;
rom[116863] = 12'hbbb;
rom[116864] = 12'hbbb;
rom[116865] = 12'hbbb;
rom[116866] = 12'hbbb;
rom[116867] = 12'hbbb;
rom[116868] = 12'hbbb;
rom[116869] = 12'hbbb;
rom[116870] = 12'hbbb;
rom[116871] = 12'hbbb;
rom[116872] = 12'hbbb;
rom[116873] = 12'hbbb;
rom[116874] = 12'hccc;
rom[116875] = 12'hddd;
rom[116876] = 12'heee;
rom[116877] = 12'hfff;
rom[116878] = 12'hfff;
rom[116879] = 12'hfff;
rom[116880] = 12'heee;
rom[116881] = 12'hccc;
rom[116882] = 12'hbbb;
rom[116883] = 12'hbbb;
rom[116884] = 12'hbbb;
rom[116885] = 12'haaa;
rom[116886] = 12'haaa;
rom[116887] = 12'haaa;
rom[116888] = 12'h999;
rom[116889] = 12'h999;
rom[116890] = 12'h999;
rom[116891] = 12'haaa;
rom[116892] = 12'h999;
rom[116893] = 12'h888;
rom[116894] = 12'h888;
rom[116895] = 12'haaa;
rom[116896] = 12'hccc;
rom[116897] = 12'hbbb;
rom[116898] = 12'hbbb;
rom[116899] = 12'h999;
rom[116900] = 12'h888;
rom[116901] = 12'h888;
rom[116902] = 12'h999;
rom[116903] = 12'haaa;
rom[116904] = 12'h888;
rom[116905] = 12'h888;
rom[116906] = 12'h777;
rom[116907] = 12'h777;
rom[116908] = 12'h777;
rom[116909] = 12'h666;
rom[116910] = 12'h666;
rom[116911] = 12'h666;
rom[116912] = 12'h666;
rom[116913] = 12'h666;
rom[116914] = 12'h666;
rom[116915] = 12'h666;
rom[116916] = 12'h666;
rom[116917] = 12'h666;
rom[116918] = 12'h666;
rom[116919] = 12'h666;
rom[116920] = 12'h666;
rom[116921] = 12'h777;
rom[116922] = 12'h777;
rom[116923] = 12'h777;
rom[116924] = 12'h666;
rom[116925] = 12'h555;
rom[116926] = 12'h555;
rom[116927] = 12'h666;
rom[116928] = 12'h777;
rom[116929] = 12'h666;
rom[116930] = 12'h555;
rom[116931] = 12'h444;
rom[116932] = 12'h444;
rom[116933] = 12'h444;
rom[116934] = 12'h555;
rom[116935] = 12'h555;
rom[116936] = 12'h555;
rom[116937] = 12'h555;
rom[116938] = 12'h444;
rom[116939] = 12'h444;
rom[116940] = 12'h444;
rom[116941] = 12'h444;
rom[116942] = 12'h444;
rom[116943] = 12'h444;
rom[116944] = 12'h444;
rom[116945] = 12'h333;
rom[116946] = 12'h333;
rom[116947] = 12'h333;
rom[116948] = 12'h333;
rom[116949] = 12'h333;
rom[116950] = 12'h333;
rom[116951] = 12'h333;
rom[116952] = 12'h333;
rom[116953] = 12'h333;
rom[116954] = 12'h444;
rom[116955] = 12'h444;
rom[116956] = 12'h555;
rom[116957] = 12'h555;
rom[116958] = 12'h555;
rom[116959] = 12'h555;
rom[116960] = 12'h666;
rom[116961] = 12'h555;
rom[116962] = 12'h555;
rom[116963] = 12'h555;
rom[116964] = 12'h555;
rom[116965] = 12'h555;
rom[116966] = 12'h555;
rom[116967] = 12'h555;
rom[116968] = 12'h555;
rom[116969] = 12'h555;
rom[116970] = 12'h666;
rom[116971] = 12'h666;
rom[116972] = 12'h666;
rom[116973] = 12'h666;
rom[116974] = 12'h666;
rom[116975] = 12'h555;
rom[116976] = 12'h666;
rom[116977] = 12'h666;
rom[116978] = 12'h666;
rom[116979] = 12'h666;
rom[116980] = 12'h666;
rom[116981] = 12'h555;
rom[116982] = 12'h555;
rom[116983] = 12'h555;
rom[116984] = 12'h555;
rom[116985] = 12'h555;
rom[116986] = 12'h555;
rom[116987] = 12'h444;
rom[116988] = 12'h444;
rom[116989] = 12'h555;
rom[116990] = 12'h666;
rom[116991] = 12'h777;
rom[116992] = 12'h777;
rom[116993] = 12'h666;
rom[116994] = 12'h666;
rom[116995] = 12'h666;
rom[116996] = 12'h777;
rom[116997] = 12'h777;
rom[116998] = 12'h666;
rom[116999] = 12'h555;
rom[117000] = 12'h555;
rom[117001] = 12'h555;
rom[117002] = 12'h555;
rom[117003] = 12'h555;
rom[117004] = 12'h555;
rom[117005] = 12'h555;
rom[117006] = 12'h555;
rom[117007] = 12'h444;
rom[117008] = 12'h333;
rom[117009] = 12'h444;
rom[117010] = 12'h444;
rom[117011] = 12'h555;
rom[117012] = 12'h555;
rom[117013] = 12'h555;
rom[117014] = 12'h444;
rom[117015] = 12'h333;
rom[117016] = 12'h444;
rom[117017] = 12'h444;
rom[117018] = 12'h444;
rom[117019] = 12'h333;
rom[117020] = 12'h222;
rom[117021] = 12'h111;
rom[117022] = 12'h111;
rom[117023] = 12'h111;
rom[117024] = 12'h111;
rom[117025] = 12'h111;
rom[117026] = 12'h333;
rom[117027] = 12'h666;
rom[117028] = 12'h888;
rom[117029] = 12'h444;
rom[117030] = 12'h  0;
rom[117031] = 12'h  0;
rom[117032] = 12'h  0;
rom[117033] = 12'h  0;
rom[117034] = 12'h  0;
rom[117035] = 12'h111;
rom[117036] = 12'h222;
rom[117037] = 12'h222;
rom[117038] = 12'h333;
rom[117039] = 12'h666;
rom[117040] = 12'haaa;
rom[117041] = 12'haaa;
rom[117042] = 12'h555;
rom[117043] = 12'h111;
rom[117044] = 12'h  0;
rom[117045] = 12'h  0;
rom[117046] = 12'h  0;
rom[117047] = 12'h  0;
rom[117048] = 12'h  0;
rom[117049] = 12'h  0;
rom[117050] = 12'h  0;
rom[117051] = 12'h  0;
rom[117052] = 12'h  0;
rom[117053] = 12'h  0;
rom[117054] = 12'h  0;
rom[117055] = 12'h  0;
rom[117056] = 12'h  0;
rom[117057] = 12'h  0;
rom[117058] = 12'h  0;
rom[117059] = 12'h  0;
rom[117060] = 12'h  0;
rom[117061] = 12'h  0;
rom[117062] = 12'h  0;
rom[117063] = 12'h333;
rom[117064] = 12'haaa;
rom[117065] = 12'heee;
rom[117066] = 12'hccc;
rom[117067] = 12'h555;
rom[117068] = 12'h222;
rom[117069] = 12'h111;
rom[117070] = 12'h  0;
rom[117071] = 12'h111;
rom[117072] = 12'h111;
rom[117073] = 12'h  0;
rom[117074] = 12'h  0;
rom[117075] = 12'h222;
rom[117076] = 12'h666;
rom[117077] = 12'hccc;
rom[117078] = 12'hbbb;
rom[117079] = 12'h555;
rom[117080] = 12'h111;
rom[117081] = 12'h  0;
rom[117082] = 12'h  0;
rom[117083] = 12'h111;
rom[117084] = 12'h  0;
rom[117085] = 12'h  0;
rom[117086] = 12'h  0;
rom[117087] = 12'h  0;
rom[117088] = 12'h111;
rom[117089] = 12'h111;
rom[117090] = 12'h333;
rom[117091] = 12'h666;
rom[117092] = 12'h666;
rom[117093] = 12'h333;
rom[117094] = 12'h333;
rom[117095] = 12'h666;
rom[117096] = 12'h999;
rom[117097] = 12'h777;
rom[117098] = 12'h333;
rom[117099] = 12'h111;
rom[117100] = 12'h  0;
rom[117101] = 12'h111;
rom[117102] = 12'h111;
rom[117103] = 12'h111;
rom[117104] = 12'h111;
rom[117105] = 12'h111;
rom[117106] = 12'h111;
rom[117107] = 12'h111;
rom[117108] = 12'h111;
rom[117109] = 12'h111;
rom[117110] = 12'h111;
rom[117111] = 12'h111;
rom[117112] = 12'h111;
rom[117113] = 12'h222;
rom[117114] = 12'h444;
rom[117115] = 12'h666;
rom[117116] = 12'h888;
rom[117117] = 12'h999;
rom[117118] = 12'h999;
rom[117119] = 12'h777;
rom[117120] = 12'h444;
rom[117121] = 12'h222;
rom[117122] = 12'h111;
rom[117123] = 12'h  0;
rom[117124] = 12'h  0;
rom[117125] = 12'h  0;
rom[117126] = 12'h  0;
rom[117127] = 12'h  0;
rom[117128] = 12'h  0;
rom[117129] = 12'h  0;
rom[117130] = 12'h  0;
rom[117131] = 12'h  0;
rom[117132] = 12'h  0;
rom[117133] = 12'h  0;
rom[117134] = 12'h  0;
rom[117135] = 12'h  0;
rom[117136] = 12'h  0;
rom[117137] = 12'h  0;
rom[117138] = 12'h  0;
rom[117139] = 12'h  0;
rom[117140] = 12'h  0;
rom[117141] = 12'h  0;
rom[117142] = 12'h  0;
rom[117143] = 12'h  0;
rom[117144] = 12'h  0;
rom[117145] = 12'h  0;
rom[117146] = 12'h  0;
rom[117147] = 12'h  0;
rom[117148] = 12'h  0;
rom[117149] = 12'h  0;
rom[117150] = 12'h  0;
rom[117151] = 12'h  0;
rom[117152] = 12'h  0;
rom[117153] = 12'h  0;
rom[117154] = 12'h  0;
rom[117155] = 12'h  0;
rom[117156] = 12'h  0;
rom[117157] = 12'h  0;
rom[117158] = 12'h  0;
rom[117159] = 12'h  0;
rom[117160] = 12'h  0;
rom[117161] = 12'h  0;
rom[117162] = 12'h  0;
rom[117163] = 12'h  0;
rom[117164] = 12'h  0;
rom[117165] = 12'h  0;
rom[117166] = 12'h  0;
rom[117167] = 12'h  0;
rom[117168] = 12'h111;
rom[117169] = 12'h111;
rom[117170] = 12'h222;
rom[117171] = 12'h444;
rom[117172] = 12'h888;
rom[117173] = 12'haaa;
rom[117174] = 12'h888;
rom[117175] = 12'h555;
rom[117176] = 12'h222;
rom[117177] = 12'h111;
rom[117178] = 12'h  0;
rom[117179] = 12'h  0;
rom[117180] = 12'h  0;
rom[117181] = 12'h  0;
rom[117182] = 12'h  0;
rom[117183] = 12'h  0;
rom[117184] = 12'h  0;
rom[117185] = 12'h  0;
rom[117186] = 12'h  0;
rom[117187] = 12'h  0;
rom[117188] = 12'h  0;
rom[117189] = 12'h  0;
rom[117190] = 12'h  0;
rom[117191] = 12'h  0;
rom[117192] = 12'h  0;
rom[117193] = 12'h  0;
rom[117194] = 12'h  0;
rom[117195] = 12'h  0;
rom[117196] = 12'h  0;
rom[117197] = 12'h  0;
rom[117198] = 12'h  0;
rom[117199] = 12'h  0;
rom[117200] = 12'hfff;
rom[117201] = 12'hfff;
rom[117202] = 12'hfff;
rom[117203] = 12'hfff;
rom[117204] = 12'hfff;
rom[117205] = 12'hfff;
rom[117206] = 12'heee;
rom[117207] = 12'heee;
rom[117208] = 12'heee;
rom[117209] = 12'heee;
rom[117210] = 12'heee;
rom[117211] = 12'heee;
rom[117212] = 12'heee;
rom[117213] = 12'heee;
rom[117214] = 12'heee;
rom[117215] = 12'heee;
rom[117216] = 12'heee;
rom[117217] = 12'heee;
rom[117218] = 12'heee;
rom[117219] = 12'heee;
rom[117220] = 12'heee;
rom[117221] = 12'heee;
rom[117222] = 12'heee;
rom[117223] = 12'heee;
rom[117224] = 12'heee;
rom[117225] = 12'heee;
rom[117226] = 12'heee;
rom[117227] = 12'heee;
rom[117228] = 12'heee;
rom[117229] = 12'heee;
rom[117230] = 12'hddd;
rom[117231] = 12'hddd;
rom[117232] = 12'hddd;
rom[117233] = 12'hddd;
rom[117234] = 12'hddd;
rom[117235] = 12'hddd;
rom[117236] = 12'hddd;
rom[117237] = 12'hddd;
rom[117238] = 12'hddd;
rom[117239] = 12'hddd;
rom[117240] = 12'hddd;
rom[117241] = 12'hddd;
rom[117242] = 12'hccc;
rom[117243] = 12'hccc;
rom[117244] = 12'hccc;
rom[117245] = 12'hccc;
rom[117246] = 12'hccc;
rom[117247] = 12'hccc;
rom[117248] = 12'hccc;
rom[117249] = 12'hccc;
rom[117250] = 12'hccc;
rom[117251] = 12'hccc;
rom[117252] = 12'hccc;
rom[117253] = 12'hccc;
rom[117254] = 12'hccc;
rom[117255] = 12'hccc;
rom[117256] = 12'hccc;
rom[117257] = 12'hccc;
rom[117258] = 12'hccc;
rom[117259] = 12'hbbb;
rom[117260] = 12'hbbb;
rom[117261] = 12'hbbb;
rom[117262] = 12'hbbb;
rom[117263] = 12'hbbb;
rom[117264] = 12'hbbb;
rom[117265] = 12'hbbb;
rom[117266] = 12'hbbb;
rom[117267] = 12'hbbb;
rom[117268] = 12'hbbb;
rom[117269] = 12'hbbb;
rom[117270] = 12'hbbb;
rom[117271] = 12'hbbb;
rom[117272] = 12'hbbb;
rom[117273] = 12'hbbb;
rom[117274] = 12'hccc;
rom[117275] = 12'heee;
rom[117276] = 12'hfff;
rom[117277] = 12'hfff;
rom[117278] = 12'hfff;
rom[117279] = 12'heee;
rom[117280] = 12'hccc;
rom[117281] = 12'hbbb;
rom[117282] = 12'haaa;
rom[117283] = 12'haaa;
rom[117284] = 12'haaa;
rom[117285] = 12'haaa;
rom[117286] = 12'h999;
rom[117287] = 12'h999;
rom[117288] = 12'h999;
rom[117289] = 12'h999;
rom[117290] = 12'h999;
rom[117291] = 12'h999;
rom[117292] = 12'h888;
rom[117293] = 12'h777;
rom[117294] = 12'h999;
rom[117295] = 12'hbbb;
rom[117296] = 12'hccc;
rom[117297] = 12'hbbb;
rom[117298] = 12'h999;
rom[117299] = 12'h888;
rom[117300] = 12'h888;
rom[117301] = 12'h888;
rom[117302] = 12'h999;
rom[117303] = 12'h999;
rom[117304] = 12'h777;
rom[117305] = 12'h777;
rom[117306] = 12'h777;
rom[117307] = 12'h777;
rom[117308] = 12'h777;
rom[117309] = 12'h666;
rom[117310] = 12'h666;
rom[117311] = 12'h666;
rom[117312] = 12'h555;
rom[117313] = 12'h555;
rom[117314] = 12'h555;
rom[117315] = 12'h555;
rom[117316] = 12'h555;
rom[117317] = 12'h666;
rom[117318] = 12'h666;
rom[117319] = 12'h666;
rom[117320] = 12'h666;
rom[117321] = 12'h777;
rom[117322] = 12'h777;
rom[117323] = 12'h777;
rom[117324] = 12'h666;
rom[117325] = 12'h555;
rom[117326] = 12'h666;
rom[117327] = 12'h666;
rom[117328] = 12'h666;
rom[117329] = 12'h555;
rom[117330] = 12'h444;
rom[117331] = 12'h444;
rom[117332] = 12'h444;
rom[117333] = 12'h444;
rom[117334] = 12'h555;
rom[117335] = 12'h555;
rom[117336] = 12'h555;
rom[117337] = 12'h555;
rom[117338] = 12'h444;
rom[117339] = 12'h444;
rom[117340] = 12'h444;
rom[117341] = 12'h444;
rom[117342] = 12'h444;
rom[117343] = 12'h444;
rom[117344] = 12'h333;
rom[117345] = 12'h333;
rom[117346] = 12'h333;
rom[117347] = 12'h333;
rom[117348] = 12'h333;
rom[117349] = 12'h333;
rom[117350] = 12'h333;
rom[117351] = 12'h333;
rom[117352] = 12'h333;
rom[117353] = 12'h333;
rom[117354] = 12'h444;
rom[117355] = 12'h444;
rom[117356] = 12'h444;
rom[117357] = 12'h555;
rom[117358] = 12'h555;
rom[117359] = 12'h555;
rom[117360] = 12'h555;
rom[117361] = 12'h555;
rom[117362] = 12'h555;
rom[117363] = 12'h555;
rom[117364] = 12'h555;
rom[117365] = 12'h555;
rom[117366] = 12'h555;
rom[117367] = 12'h555;
rom[117368] = 12'h555;
rom[117369] = 12'h555;
rom[117370] = 12'h555;
rom[117371] = 12'h666;
rom[117372] = 12'h666;
rom[117373] = 12'h666;
rom[117374] = 12'h555;
rom[117375] = 12'h555;
rom[117376] = 12'h555;
rom[117377] = 12'h555;
rom[117378] = 12'h555;
rom[117379] = 12'h666;
rom[117380] = 12'h555;
rom[117381] = 12'h555;
rom[117382] = 12'h444;
rom[117383] = 12'h555;
rom[117384] = 12'h555;
rom[117385] = 12'h444;
rom[117386] = 12'h444;
rom[117387] = 12'h444;
rom[117388] = 12'h444;
rom[117389] = 12'h555;
rom[117390] = 12'h666;
rom[117391] = 12'h666;
rom[117392] = 12'h777;
rom[117393] = 12'h666;
rom[117394] = 12'h555;
rom[117395] = 12'h666;
rom[117396] = 12'h666;
rom[117397] = 12'h666;
rom[117398] = 12'h555;
rom[117399] = 12'h555;
rom[117400] = 12'h444;
rom[117401] = 12'h444;
rom[117402] = 12'h444;
rom[117403] = 12'h444;
rom[117404] = 12'h444;
rom[117405] = 12'h555;
rom[117406] = 12'h444;
rom[117407] = 12'h444;
rom[117408] = 12'h333;
rom[117409] = 12'h333;
rom[117410] = 12'h333;
rom[117411] = 12'h444;
rom[117412] = 12'h555;
rom[117413] = 12'h555;
rom[117414] = 12'h444;
rom[117415] = 12'h333;
rom[117416] = 12'h333;
rom[117417] = 12'h333;
rom[117418] = 12'h444;
rom[117419] = 12'h333;
rom[117420] = 12'h222;
rom[117421] = 12'h111;
rom[117422] = 12'h  0;
rom[117423] = 12'h111;
rom[117424] = 12'h111;
rom[117425] = 12'h111;
rom[117426] = 12'h  0;
rom[117427] = 12'h444;
rom[117428] = 12'h888;
rom[117429] = 12'h666;
rom[117430] = 12'h111;
rom[117431] = 12'h111;
rom[117432] = 12'h  0;
rom[117433] = 12'h  0;
rom[117434] = 12'h  0;
rom[117435] = 12'h111;
rom[117436] = 12'h222;
rom[117437] = 12'h222;
rom[117438] = 12'h444;
rom[117439] = 12'h777;
rom[117440] = 12'haaa;
rom[117441] = 12'h888;
rom[117442] = 12'h444;
rom[117443] = 12'h  0;
rom[117444] = 12'h  0;
rom[117445] = 12'h  0;
rom[117446] = 12'h  0;
rom[117447] = 12'h  0;
rom[117448] = 12'h  0;
rom[117449] = 12'h  0;
rom[117450] = 12'h  0;
rom[117451] = 12'h  0;
rom[117452] = 12'h  0;
rom[117453] = 12'h  0;
rom[117454] = 12'h  0;
rom[117455] = 12'h  0;
rom[117456] = 12'h  0;
rom[117457] = 12'h  0;
rom[117458] = 12'h  0;
rom[117459] = 12'h  0;
rom[117460] = 12'h  0;
rom[117461] = 12'h  0;
rom[117462] = 12'h  0;
rom[117463] = 12'h333;
rom[117464] = 12'hbbb;
rom[117465] = 12'heee;
rom[117466] = 12'hbbb;
rom[117467] = 12'h555;
rom[117468] = 12'h222;
rom[117469] = 12'h111;
rom[117470] = 12'h  0;
rom[117471] = 12'h111;
rom[117472] = 12'h  0;
rom[117473] = 12'h  0;
rom[117474] = 12'h  0;
rom[117475] = 12'h111;
rom[117476] = 12'h555;
rom[117477] = 12'hbbb;
rom[117478] = 12'hbbb;
rom[117479] = 12'h666;
rom[117480] = 12'h111;
rom[117481] = 12'h  0;
rom[117482] = 12'h  0;
rom[117483] = 12'h111;
rom[117484] = 12'h  0;
rom[117485] = 12'h  0;
rom[117486] = 12'h  0;
rom[117487] = 12'h  0;
rom[117488] = 12'h  0;
rom[117489] = 12'h111;
rom[117490] = 12'h222;
rom[117491] = 12'h555;
rom[117492] = 12'h666;
rom[117493] = 12'h333;
rom[117494] = 12'h222;
rom[117495] = 12'h444;
rom[117496] = 12'h777;
rom[117497] = 12'h777;
rom[117498] = 12'h555;
rom[117499] = 12'h222;
rom[117500] = 12'h  0;
rom[117501] = 12'h111;
rom[117502] = 12'h111;
rom[117503] = 12'h111;
rom[117504] = 12'h111;
rom[117505] = 12'h111;
rom[117506] = 12'h111;
rom[117507] = 12'h111;
rom[117508] = 12'h111;
rom[117509] = 12'h111;
rom[117510] = 12'h111;
rom[117511] = 12'h111;
rom[117512] = 12'h111;
rom[117513] = 12'h222;
rom[117514] = 12'h333;
rom[117515] = 12'h555;
rom[117516] = 12'h777;
rom[117517] = 12'h888;
rom[117518] = 12'h888;
rom[117519] = 12'h888;
rom[117520] = 12'h555;
rom[117521] = 12'h333;
rom[117522] = 12'h111;
rom[117523] = 12'h  0;
rom[117524] = 12'h  0;
rom[117525] = 12'h  0;
rom[117526] = 12'h  0;
rom[117527] = 12'h  0;
rom[117528] = 12'h  0;
rom[117529] = 12'h  0;
rom[117530] = 12'h  0;
rom[117531] = 12'h  0;
rom[117532] = 12'h  0;
rom[117533] = 12'h  0;
rom[117534] = 12'h  0;
rom[117535] = 12'h  0;
rom[117536] = 12'h  0;
rom[117537] = 12'h  0;
rom[117538] = 12'h  0;
rom[117539] = 12'h  0;
rom[117540] = 12'h  0;
rom[117541] = 12'h  0;
rom[117542] = 12'h  0;
rom[117543] = 12'h  0;
rom[117544] = 12'h  0;
rom[117545] = 12'h  0;
rom[117546] = 12'h  0;
rom[117547] = 12'h  0;
rom[117548] = 12'h  0;
rom[117549] = 12'h  0;
rom[117550] = 12'h  0;
rom[117551] = 12'h  0;
rom[117552] = 12'h  0;
rom[117553] = 12'h  0;
rom[117554] = 12'h  0;
rom[117555] = 12'h  0;
rom[117556] = 12'h  0;
rom[117557] = 12'h  0;
rom[117558] = 12'h  0;
rom[117559] = 12'h  0;
rom[117560] = 12'h  0;
rom[117561] = 12'h  0;
rom[117562] = 12'h  0;
rom[117563] = 12'h  0;
rom[117564] = 12'h  0;
rom[117565] = 12'h  0;
rom[117566] = 12'h  0;
rom[117567] = 12'h  0;
rom[117568] = 12'h111;
rom[117569] = 12'h111;
rom[117570] = 12'h111;
rom[117571] = 12'h333;
rom[117572] = 12'h666;
rom[117573] = 12'haaa;
rom[117574] = 12'h999;
rom[117575] = 12'h777;
rom[117576] = 12'h444;
rom[117577] = 12'h222;
rom[117578] = 12'h  0;
rom[117579] = 12'h  0;
rom[117580] = 12'h  0;
rom[117581] = 12'h  0;
rom[117582] = 12'h  0;
rom[117583] = 12'h  0;
rom[117584] = 12'h  0;
rom[117585] = 12'h  0;
rom[117586] = 12'h  0;
rom[117587] = 12'h  0;
rom[117588] = 12'h  0;
rom[117589] = 12'h  0;
rom[117590] = 12'h  0;
rom[117591] = 12'h  0;
rom[117592] = 12'h  0;
rom[117593] = 12'h  0;
rom[117594] = 12'h  0;
rom[117595] = 12'h  0;
rom[117596] = 12'h  0;
rom[117597] = 12'h  0;
rom[117598] = 12'h  0;
rom[117599] = 12'h  0;
rom[117600] = 12'hfff;
rom[117601] = 12'hfff;
rom[117602] = 12'hfff;
rom[117603] = 12'hfff;
rom[117604] = 12'hfff;
rom[117605] = 12'heee;
rom[117606] = 12'heee;
rom[117607] = 12'heee;
rom[117608] = 12'heee;
rom[117609] = 12'heee;
rom[117610] = 12'heee;
rom[117611] = 12'heee;
rom[117612] = 12'heee;
rom[117613] = 12'heee;
rom[117614] = 12'heee;
rom[117615] = 12'heee;
rom[117616] = 12'heee;
rom[117617] = 12'heee;
rom[117618] = 12'heee;
rom[117619] = 12'heee;
rom[117620] = 12'heee;
rom[117621] = 12'heee;
rom[117622] = 12'heee;
rom[117623] = 12'heee;
rom[117624] = 12'heee;
rom[117625] = 12'heee;
rom[117626] = 12'hddd;
rom[117627] = 12'hddd;
rom[117628] = 12'hddd;
rom[117629] = 12'hddd;
rom[117630] = 12'hddd;
rom[117631] = 12'hddd;
rom[117632] = 12'hddd;
rom[117633] = 12'hddd;
rom[117634] = 12'hddd;
rom[117635] = 12'hddd;
rom[117636] = 12'hddd;
rom[117637] = 12'hddd;
rom[117638] = 12'hddd;
rom[117639] = 12'hddd;
rom[117640] = 12'hccc;
rom[117641] = 12'hccc;
rom[117642] = 12'hccc;
rom[117643] = 12'hccc;
rom[117644] = 12'hccc;
rom[117645] = 12'hccc;
rom[117646] = 12'hccc;
rom[117647] = 12'hccc;
rom[117648] = 12'hccc;
rom[117649] = 12'hccc;
rom[117650] = 12'hccc;
rom[117651] = 12'hccc;
rom[117652] = 12'hccc;
rom[117653] = 12'hccc;
rom[117654] = 12'hccc;
rom[117655] = 12'hccc;
rom[117656] = 12'hccc;
rom[117657] = 12'hccc;
rom[117658] = 12'hccc;
rom[117659] = 12'hbbb;
rom[117660] = 12'hbbb;
rom[117661] = 12'hbbb;
rom[117662] = 12'hbbb;
rom[117663] = 12'hbbb;
rom[117664] = 12'hbbb;
rom[117665] = 12'hbbb;
rom[117666] = 12'hbbb;
rom[117667] = 12'hbbb;
rom[117668] = 12'hbbb;
rom[117669] = 12'hbbb;
rom[117670] = 12'hbbb;
rom[117671] = 12'hbbb;
rom[117672] = 12'hbbb;
rom[117673] = 12'hccc;
rom[117674] = 12'hddd;
rom[117675] = 12'heee;
rom[117676] = 12'hfff;
rom[117677] = 12'hfff;
rom[117678] = 12'heee;
rom[117679] = 12'hddd;
rom[117680] = 12'hbbb;
rom[117681] = 12'hbbb;
rom[117682] = 12'haaa;
rom[117683] = 12'haaa;
rom[117684] = 12'haaa;
rom[117685] = 12'h999;
rom[117686] = 12'h999;
rom[117687] = 12'h999;
rom[117688] = 12'h999;
rom[117689] = 12'h999;
rom[117690] = 12'h999;
rom[117691] = 12'h888;
rom[117692] = 12'h888;
rom[117693] = 12'h888;
rom[117694] = 12'haaa;
rom[117695] = 12'hccc;
rom[117696] = 12'hbbb;
rom[117697] = 12'haaa;
rom[117698] = 12'h999;
rom[117699] = 12'h888;
rom[117700] = 12'h777;
rom[117701] = 12'h888;
rom[117702] = 12'h999;
rom[117703] = 12'h888;
rom[117704] = 12'h777;
rom[117705] = 12'h777;
rom[117706] = 12'h777;
rom[117707] = 12'h777;
rom[117708] = 12'h666;
rom[117709] = 12'h666;
rom[117710] = 12'h666;
rom[117711] = 12'h555;
rom[117712] = 12'h555;
rom[117713] = 12'h555;
rom[117714] = 12'h555;
rom[117715] = 12'h555;
rom[117716] = 12'h555;
rom[117717] = 12'h555;
rom[117718] = 12'h555;
rom[117719] = 12'h555;
rom[117720] = 12'h666;
rom[117721] = 12'h666;
rom[117722] = 12'h777;
rom[117723] = 12'h666;
rom[117724] = 12'h666;
rom[117725] = 12'h666;
rom[117726] = 12'h666;
rom[117727] = 12'h666;
rom[117728] = 12'h666;
rom[117729] = 12'h555;
rom[117730] = 12'h444;
rom[117731] = 12'h444;
rom[117732] = 12'h444;
rom[117733] = 12'h555;
rom[117734] = 12'h555;
rom[117735] = 12'h555;
rom[117736] = 12'h555;
rom[117737] = 12'h444;
rom[117738] = 12'h333;
rom[117739] = 12'h333;
rom[117740] = 12'h333;
rom[117741] = 12'h444;
rom[117742] = 12'h444;
rom[117743] = 12'h444;
rom[117744] = 12'h444;
rom[117745] = 12'h333;
rom[117746] = 12'h333;
rom[117747] = 12'h333;
rom[117748] = 12'h333;
rom[117749] = 12'h333;
rom[117750] = 12'h333;
rom[117751] = 12'h333;
rom[117752] = 12'h333;
rom[117753] = 12'h333;
rom[117754] = 12'h444;
rom[117755] = 12'h444;
rom[117756] = 12'h444;
rom[117757] = 12'h555;
rom[117758] = 12'h555;
rom[117759] = 12'h555;
rom[117760] = 12'h555;
rom[117761] = 12'h555;
rom[117762] = 12'h444;
rom[117763] = 12'h444;
rom[117764] = 12'h444;
rom[117765] = 12'h444;
rom[117766] = 12'h444;
rom[117767] = 12'h444;
rom[117768] = 12'h555;
rom[117769] = 12'h555;
rom[117770] = 12'h555;
rom[117771] = 12'h555;
rom[117772] = 12'h555;
rom[117773] = 12'h555;
rom[117774] = 12'h555;
rom[117775] = 12'h444;
rom[117776] = 12'h555;
rom[117777] = 12'h555;
rom[117778] = 12'h555;
rom[117779] = 12'h555;
rom[117780] = 12'h555;
rom[117781] = 12'h444;
rom[117782] = 12'h444;
rom[117783] = 12'h444;
rom[117784] = 12'h444;
rom[117785] = 12'h444;
rom[117786] = 12'h444;
rom[117787] = 12'h333;
rom[117788] = 12'h333;
rom[117789] = 12'h444;
rom[117790] = 12'h555;
rom[117791] = 12'h555;
rom[117792] = 12'h777;
rom[117793] = 12'h666;
rom[117794] = 12'h555;
rom[117795] = 12'h555;
rom[117796] = 12'h666;
rom[117797] = 12'h555;
rom[117798] = 12'h444;
rom[117799] = 12'h444;
rom[117800] = 12'h333;
rom[117801] = 12'h333;
rom[117802] = 12'h333;
rom[117803] = 12'h333;
rom[117804] = 12'h444;
rom[117805] = 12'h444;
rom[117806] = 12'h444;
rom[117807] = 12'h444;
rom[117808] = 12'h333;
rom[117809] = 12'h333;
rom[117810] = 12'h333;
rom[117811] = 12'h333;
rom[117812] = 12'h444;
rom[117813] = 12'h444;
rom[117814] = 12'h444;
rom[117815] = 12'h333;
rom[117816] = 12'h222;
rom[117817] = 12'h333;
rom[117818] = 12'h333;
rom[117819] = 12'h333;
rom[117820] = 12'h222;
rom[117821] = 12'h  0;
rom[117822] = 12'h  0;
rom[117823] = 12'h  0;
rom[117824] = 12'h111;
rom[117825] = 12'h  0;
rom[117826] = 12'h  0;
rom[117827] = 12'h222;
rom[117828] = 12'h555;
rom[117829] = 12'h666;
rom[117830] = 12'h444;
rom[117831] = 12'h222;
rom[117832] = 12'h111;
rom[117833] = 12'h  0;
rom[117834] = 12'h  0;
rom[117835] = 12'h111;
rom[117836] = 12'h111;
rom[117837] = 12'h333;
rom[117838] = 12'h666;
rom[117839] = 12'h888;
rom[117840] = 12'h999;
rom[117841] = 12'h666;
rom[117842] = 12'h222;
rom[117843] = 12'h  0;
rom[117844] = 12'h  0;
rom[117845] = 12'h  0;
rom[117846] = 12'h  0;
rom[117847] = 12'h  0;
rom[117848] = 12'h  0;
rom[117849] = 12'h  0;
rom[117850] = 12'h  0;
rom[117851] = 12'h  0;
rom[117852] = 12'h  0;
rom[117853] = 12'h  0;
rom[117854] = 12'h  0;
rom[117855] = 12'h  0;
rom[117856] = 12'h  0;
rom[117857] = 12'h  0;
rom[117858] = 12'h  0;
rom[117859] = 12'h  0;
rom[117860] = 12'h  0;
rom[117861] = 12'h  0;
rom[117862] = 12'h  0;
rom[117863] = 12'h333;
rom[117864] = 12'hbbb;
rom[117865] = 12'heee;
rom[117866] = 12'hbbb;
rom[117867] = 12'h555;
rom[117868] = 12'h222;
rom[117869] = 12'h111;
rom[117870] = 12'h111;
rom[117871] = 12'h111;
rom[117872] = 12'h  0;
rom[117873] = 12'h  0;
rom[117874] = 12'h  0;
rom[117875] = 12'h111;
rom[117876] = 12'h333;
rom[117877] = 12'haaa;
rom[117878] = 12'hbbb;
rom[117879] = 12'h777;
rom[117880] = 12'h222;
rom[117881] = 12'h  0;
rom[117882] = 12'h  0;
rom[117883] = 12'h111;
rom[117884] = 12'h  0;
rom[117885] = 12'h  0;
rom[117886] = 12'h  0;
rom[117887] = 12'h  0;
rom[117888] = 12'h  0;
rom[117889] = 12'h111;
rom[117890] = 12'h222;
rom[117891] = 12'h444;
rom[117892] = 12'h555;
rom[117893] = 12'h444;
rom[117894] = 12'h222;
rom[117895] = 12'h222;
rom[117896] = 12'h666;
rom[117897] = 12'h777;
rom[117898] = 12'h666;
rom[117899] = 12'h333;
rom[117900] = 12'h111;
rom[117901] = 12'h111;
rom[117902] = 12'h111;
rom[117903] = 12'h111;
rom[117904] = 12'h111;
rom[117905] = 12'h111;
rom[117906] = 12'h  0;
rom[117907] = 12'h  0;
rom[117908] = 12'h  0;
rom[117909] = 12'h111;
rom[117910] = 12'h  0;
rom[117911] = 12'h  0;
rom[117912] = 12'h111;
rom[117913] = 12'h111;
rom[117914] = 12'h222;
rom[117915] = 12'h444;
rom[117916] = 12'h666;
rom[117917] = 12'h777;
rom[117918] = 12'h888;
rom[117919] = 12'h888;
rom[117920] = 12'h666;
rom[117921] = 12'h333;
rom[117922] = 12'h111;
rom[117923] = 12'h111;
rom[117924] = 12'h  0;
rom[117925] = 12'h  0;
rom[117926] = 12'h  0;
rom[117927] = 12'h  0;
rom[117928] = 12'h  0;
rom[117929] = 12'h  0;
rom[117930] = 12'h  0;
rom[117931] = 12'h  0;
rom[117932] = 12'h  0;
rom[117933] = 12'h  0;
rom[117934] = 12'h  0;
rom[117935] = 12'h  0;
rom[117936] = 12'h  0;
rom[117937] = 12'h  0;
rom[117938] = 12'h  0;
rom[117939] = 12'h  0;
rom[117940] = 12'h  0;
rom[117941] = 12'h  0;
rom[117942] = 12'h  0;
rom[117943] = 12'h  0;
rom[117944] = 12'h  0;
rom[117945] = 12'h  0;
rom[117946] = 12'h  0;
rom[117947] = 12'h  0;
rom[117948] = 12'h  0;
rom[117949] = 12'h  0;
rom[117950] = 12'h  0;
rom[117951] = 12'h  0;
rom[117952] = 12'h  0;
rom[117953] = 12'h  0;
rom[117954] = 12'h  0;
rom[117955] = 12'h  0;
rom[117956] = 12'h  0;
rom[117957] = 12'h  0;
rom[117958] = 12'h  0;
rom[117959] = 12'h  0;
rom[117960] = 12'h  0;
rom[117961] = 12'h  0;
rom[117962] = 12'h  0;
rom[117963] = 12'h  0;
rom[117964] = 12'h  0;
rom[117965] = 12'h  0;
rom[117966] = 12'h  0;
rom[117967] = 12'h  0;
rom[117968] = 12'h  0;
rom[117969] = 12'h111;
rom[117970] = 12'h111;
rom[117971] = 12'h222;
rom[117972] = 12'h444;
rom[117973] = 12'h888;
rom[117974] = 12'h999;
rom[117975] = 12'h888;
rom[117976] = 12'h555;
rom[117977] = 12'h333;
rom[117978] = 12'h111;
rom[117979] = 12'h  0;
rom[117980] = 12'h  0;
rom[117981] = 12'h  0;
rom[117982] = 12'h  0;
rom[117983] = 12'h  0;
rom[117984] = 12'h  0;
rom[117985] = 12'h  0;
rom[117986] = 12'h  0;
rom[117987] = 12'h  0;
rom[117988] = 12'h  0;
rom[117989] = 12'h  0;
rom[117990] = 12'h  0;
rom[117991] = 12'h  0;
rom[117992] = 12'h  0;
rom[117993] = 12'h  0;
rom[117994] = 12'h  0;
rom[117995] = 12'h  0;
rom[117996] = 12'h  0;
rom[117997] = 12'h  0;
rom[117998] = 12'h  0;
rom[117999] = 12'h  0;
rom[118000] = 12'hfff;
rom[118001] = 12'hfff;
rom[118002] = 12'hfff;
rom[118003] = 12'hfff;
rom[118004] = 12'heee;
rom[118005] = 12'heee;
rom[118006] = 12'heee;
rom[118007] = 12'heee;
rom[118008] = 12'heee;
rom[118009] = 12'heee;
rom[118010] = 12'heee;
rom[118011] = 12'heee;
rom[118012] = 12'heee;
rom[118013] = 12'heee;
rom[118014] = 12'heee;
rom[118015] = 12'heee;
rom[118016] = 12'heee;
rom[118017] = 12'heee;
rom[118018] = 12'heee;
rom[118019] = 12'heee;
rom[118020] = 12'heee;
rom[118021] = 12'heee;
rom[118022] = 12'hddd;
rom[118023] = 12'hddd;
rom[118024] = 12'hddd;
rom[118025] = 12'hddd;
rom[118026] = 12'hddd;
rom[118027] = 12'hddd;
rom[118028] = 12'hddd;
rom[118029] = 12'hddd;
rom[118030] = 12'hddd;
rom[118031] = 12'hddd;
rom[118032] = 12'hddd;
rom[118033] = 12'hddd;
rom[118034] = 12'hddd;
rom[118035] = 12'hddd;
rom[118036] = 12'hccc;
rom[118037] = 12'hccc;
rom[118038] = 12'hccc;
rom[118039] = 12'hccc;
rom[118040] = 12'hccc;
rom[118041] = 12'hccc;
rom[118042] = 12'hccc;
rom[118043] = 12'hccc;
rom[118044] = 12'hccc;
rom[118045] = 12'hccc;
rom[118046] = 12'hccc;
rom[118047] = 12'hccc;
rom[118048] = 12'hccc;
rom[118049] = 12'hccc;
rom[118050] = 12'hccc;
rom[118051] = 12'hccc;
rom[118052] = 12'hccc;
rom[118053] = 12'hccc;
rom[118054] = 12'hccc;
rom[118055] = 12'hccc;
rom[118056] = 12'hccc;
rom[118057] = 12'hccc;
rom[118058] = 12'hccc;
rom[118059] = 12'hbbb;
rom[118060] = 12'hbbb;
rom[118061] = 12'hbbb;
rom[118062] = 12'hbbb;
rom[118063] = 12'hbbb;
rom[118064] = 12'hbbb;
rom[118065] = 12'hbbb;
rom[118066] = 12'hbbb;
rom[118067] = 12'hbbb;
rom[118068] = 12'hbbb;
rom[118069] = 12'hbbb;
rom[118070] = 12'hbbb;
rom[118071] = 12'hbbb;
rom[118072] = 12'hccc;
rom[118073] = 12'hccc;
rom[118074] = 12'heee;
rom[118075] = 12'hfff;
rom[118076] = 12'hfff;
rom[118077] = 12'hfff;
rom[118078] = 12'hddd;
rom[118079] = 12'hbbb;
rom[118080] = 12'haaa;
rom[118081] = 12'hbbb;
rom[118082] = 12'haaa;
rom[118083] = 12'haaa;
rom[118084] = 12'h999;
rom[118085] = 12'h999;
rom[118086] = 12'h999;
rom[118087] = 12'h999;
rom[118088] = 12'h999;
rom[118089] = 12'h999;
rom[118090] = 12'h999;
rom[118091] = 12'h888;
rom[118092] = 12'h888;
rom[118093] = 12'h999;
rom[118094] = 12'hbbb;
rom[118095] = 12'hddd;
rom[118096] = 12'hbbb;
rom[118097] = 12'h999;
rom[118098] = 12'h888;
rom[118099] = 12'h888;
rom[118100] = 12'h777;
rom[118101] = 12'h888;
rom[118102] = 12'h999;
rom[118103] = 12'h777;
rom[118104] = 12'h666;
rom[118105] = 12'h777;
rom[118106] = 12'h777;
rom[118107] = 12'h777;
rom[118108] = 12'h666;
rom[118109] = 12'h666;
rom[118110] = 12'h666;
rom[118111] = 12'h555;
rom[118112] = 12'h555;
rom[118113] = 12'h555;
rom[118114] = 12'h555;
rom[118115] = 12'h555;
rom[118116] = 12'h555;
rom[118117] = 12'h555;
rom[118118] = 12'h555;
rom[118119] = 12'h555;
rom[118120] = 12'h666;
rom[118121] = 12'h666;
rom[118122] = 12'h666;
rom[118123] = 12'h666;
rom[118124] = 12'h666;
rom[118125] = 12'h666;
rom[118126] = 12'h666;
rom[118127] = 12'h666;
rom[118128] = 12'h666;
rom[118129] = 12'h555;
rom[118130] = 12'h444;
rom[118131] = 12'h444;
rom[118132] = 12'h555;
rom[118133] = 12'h555;
rom[118134] = 12'h555;
rom[118135] = 12'h555;
rom[118136] = 12'h555;
rom[118137] = 12'h444;
rom[118138] = 12'h333;
rom[118139] = 12'h333;
rom[118140] = 12'h333;
rom[118141] = 12'h444;
rom[118142] = 12'h444;
rom[118143] = 12'h444;
rom[118144] = 12'h444;
rom[118145] = 12'h333;
rom[118146] = 12'h333;
rom[118147] = 12'h333;
rom[118148] = 12'h333;
rom[118149] = 12'h333;
rom[118150] = 12'h333;
rom[118151] = 12'h333;
rom[118152] = 12'h333;
rom[118153] = 12'h444;
rom[118154] = 12'h444;
rom[118155] = 12'h444;
rom[118156] = 12'h444;
rom[118157] = 12'h555;
rom[118158] = 12'h555;
rom[118159] = 12'h555;
rom[118160] = 12'h444;
rom[118161] = 12'h444;
rom[118162] = 12'h444;
rom[118163] = 12'h444;
rom[118164] = 12'h444;
rom[118165] = 12'h444;
rom[118166] = 12'h444;
rom[118167] = 12'h444;
rom[118168] = 12'h444;
rom[118169] = 12'h555;
rom[118170] = 12'h555;
rom[118171] = 12'h555;
rom[118172] = 12'h555;
rom[118173] = 12'h444;
rom[118174] = 12'h444;
rom[118175] = 12'h444;
rom[118176] = 12'h444;
rom[118177] = 12'h444;
rom[118178] = 12'h444;
rom[118179] = 12'h555;
rom[118180] = 12'h555;
rom[118181] = 12'h444;
rom[118182] = 12'h333;
rom[118183] = 12'h444;
rom[118184] = 12'h444;
rom[118185] = 12'h444;
rom[118186] = 12'h333;
rom[118187] = 12'h333;
rom[118188] = 12'h333;
rom[118189] = 12'h333;
rom[118190] = 12'h444;
rom[118191] = 12'h555;
rom[118192] = 12'h666;
rom[118193] = 12'h555;
rom[118194] = 12'h555;
rom[118195] = 12'h555;
rom[118196] = 12'h555;
rom[118197] = 12'h555;
rom[118198] = 12'h444;
rom[118199] = 12'h333;
rom[118200] = 12'h333;
rom[118201] = 12'h333;
rom[118202] = 12'h333;
rom[118203] = 12'h333;
rom[118204] = 12'h333;
rom[118205] = 12'h444;
rom[118206] = 12'h444;
rom[118207] = 12'h333;
rom[118208] = 12'h333;
rom[118209] = 12'h222;
rom[118210] = 12'h222;
rom[118211] = 12'h222;
rom[118212] = 12'h333;
rom[118213] = 12'h444;
rom[118214] = 12'h444;
rom[118215] = 12'h333;
rom[118216] = 12'h222;
rom[118217] = 12'h222;
rom[118218] = 12'h333;
rom[118219] = 12'h333;
rom[118220] = 12'h222;
rom[118221] = 12'h  0;
rom[118222] = 12'h  0;
rom[118223] = 12'h  0;
rom[118224] = 12'h111;
rom[118225] = 12'h  0;
rom[118226] = 12'h  0;
rom[118227] = 12'h111;
rom[118228] = 12'h333;
rom[118229] = 12'h666;
rom[118230] = 12'h666;
rom[118231] = 12'h222;
rom[118232] = 12'h111;
rom[118233] = 12'h  0;
rom[118234] = 12'h  0;
rom[118235] = 12'h111;
rom[118236] = 12'h111;
rom[118237] = 12'h444;
rom[118238] = 12'h777;
rom[118239] = 12'h888;
rom[118240] = 12'h888;
rom[118241] = 12'h444;
rom[118242] = 12'h111;
rom[118243] = 12'h  0;
rom[118244] = 12'h  0;
rom[118245] = 12'h  0;
rom[118246] = 12'h  0;
rom[118247] = 12'h  0;
rom[118248] = 12'h  0;
rom[118249] = 12'h  0;
rom[118250] = 12'h  0;
rom[118251] = 12'h  0;
rom[118252] = 12'h  0;
rom[118253] = 12'h  0;
rom[118254] = 12'h  0;
rom[118255] = 12'h  0;
rom[118256] = 12'h  0;
rom[118257] = 12'h  0;
rom[118258] = 12'h  0;
rom[118259] = 12'h  0;
rom[118260] = 12'h  0;
rom[118261] = 12'h  0;
rom[118262] = 12'h111;
rom[118263] = 12'h444;
rom[118264] = 12'hccc;
rom[118265] = 12'heee;
rom[118266] = 12'hbbb;
rom[118267] = 12'h444;
rom[118268] = 12'h222;
rom[118269] = 12'h111;
rom[118270] = 12'h111;
rom[118271] = 12'h111;
rom[118272] = 12'h111;
rom[118273] = 12'h  0;
rom[118274] = 12'h  0;
rom[118275] = 12'h111;
rom[118276] = 12'h222;
rom[118277] = 12'h999;
rom[118278] = 12'hbbb;
rom[118279] = 12'h888;
rom[118280] = 12'h222;
rom[118281] = 12'h  0;
rom[118282] = 12'h  0;
rom[118283] = 12'h111;
rom[118284] = 12'h  0;
rom[118285] = 12'h  0;
rom[118286] = 12'h  0;
rom[118287] = 12'h  0;
rom[118288] = 12'h  0;
rom[118289] = 12'h111;
rom[118290] = 12'h222;
rom[118291] = 12'h333;
rom[118292] = 12'h555;
rom[118293] = 12'h444;
rom[118294] = 12'h222;
rom[118295] = 12'h222;
rom[118296] = 12'h444;
rom[118297] = 12'h777;
rom[118298] = 12'h666;
rom[118299] = 12'h333;
rom[118300] = 12'h222;
rom[118301] = 12'h111;
rom[118302] = 12'h  0;
rom[118303] = 12'h111;
rom[118304] = 12'h111;
rom[118305] = 12'h111;
rom[118306] = 12'h  0;
rom[118307] = 12'h  0;
rom[118308] = 12'h  0;
rom[118309] = 12'h  0;
rom[118310] = 12'h  0;
rom[118311] = 12'h  0;
rom[118312] = 12'h  0;
rom[118313] = 12'h111;
rom[118314] = 12'h222;
rom[118315] = 12'h333;
rom[118316] = 12'h555;
rom[118317] = 12'h777;
rom[118318] = 12'h888;
rom[118319] = 12'h888;
rom[118320] = 12'h666;
rom[118321] = 12'h444;
rom[118322] = 12'h222;
rom[118323] = 12'h111;
rom[118324] = 12'h  0;
rom[118325] = 12'h  0;
rom[118326] = 12'h  0;
rom[118327] = 12'h  0;
rom[118328] = 12'h  0;
rom[118329] = 12'h  0;
rom[118330] = 12'h  0;
rom[118331] = 12'h  0;
rom[118332] = 12'h  0;
rom[118333] = 12'h  0;
rom[118334] = 12'h  0;
rom[118335] = 12'h  0;
rom[118336] = 12'h  0;
rom[118337] = 12'h  0;
rom[118338] = 12'h  0;
rom[118339] = 12'h  0;
rom[118340] = 12'h  0;
rom[118341] = 12'h  0;
rom[118342] = 12'h  0;
rom[118343] = 12'h  0;
rom[118344] = 12'h  0;
rom[118345] = 12'h  0;
rom[118346] = 12'h  0;
rom[118347] = 12'h  0;
rom[118348] = 12'h  0;
rom[118349] = 12'h  0;
rom[118350] = 12'h  0;
rom[118351] = 12'h  0;
rom[118352] = 12'h  0;
rom[118353] = 12'h  0;
rom[118354] = 12'h  0;
rom[118355] = 12'h  0;
rom[118356] = 12'h  0;
rom[118357] = 12'h  0;
rom[118358] = 12'h  0;
rom[118359] = 12'h  0;
rom[118360] = 12'h  0;
rom[118361] = 12'h  0;
rom[118362] = 12'h  0;
rom[118363] = 12'h  0;
rom[118364] = 12'h  0;
rom[118365] = 12'h  0;
rom[118366] = 12'h  0;
rom[118367] = 12'h  0;
rom[118368] = 12'h  0;
rom[118369] = 12'h111;
rom[118370] = 12'h111;
rom[118371] = 12'h111;
rom[118372] = 12'h333;
rom[118373] = 12'h777;
rom[118374] = 12'h888;
rom[118375] = 12'h888;
rom[118376] = 12'h666;
rom[118377] = 12'h444;
rom[118378] = 12'h111;
rom[118379] = 12'h  0;
rom[118380] = 12'h  0;
rom[118381] = 12'h  0;
rom[118382] = 12'h  0;
rom[118383] = 12'h  0;
rom[118384] = 12'h  0;
rom[118385] = 12'h  0;
rom[118386] = 12'h  0;
rom[118387] = 12'h  0;
rom[118388] = 12'h  0;
rom[118389] = 12'h  0;
rom[118390] = 12'h  0;
rom[118391] = 12'h  0;
rom[118392] = 12'h  0;
rom[118393] = 12'h  0;
rom[118394] = 12'h  0;
rom[118395] = 12'h  0;
rom[118396] = 12'h  0;
rom[118397] = 12'h  0;
rom[118398] = 12'h  0;
rom[118399] = 12'h  0;
rom[118400] = 12'hfff;
rom[118401] = 12'hfff;
rom[118402] = 12'heee;
rom[118403] = 12'heee;
rom[118404] = 12'heee;
rom[118405] = 12'heee;
rom[118406] = 12'heee;
rom[118407] = 12'heee;
rom[118408] = 12'heee;
rom[118409] = 12'heee;
rom[118410] = 12'heee;
rom[118411] = 12'heee;
rom[118412] = 12'heee;
rom[118413] = 12'heee;
rom[118414] = 12'heee;
rom[118415] = 12'heee;
rom[118416] = 12'heee;
rom[118417] = 12'heee;
rom[118418] = 12'heee;
rom[118419] = 12'heee;
rom[118420] = 12'heee;
rom[118421] = 12'heee;
rom[118422] = 12'hddd;
rom[118423] = 12'hddd;
rom[118424] = 12'hddd;
rom[118425] = 12'hddd;
rom[118426] = 12'hddd;
rom[118427] = 12'hddd;
rom[118428] = 12'hddd;
rom[118429] = 12'hddd;
rom[118430] = 12'hddd;
rom[118431] = 12'hddd;
rom[118432] = 12'hddd;
rom[118433] = 12'hddd;
rom[118434] = 12'hddd;
rom[118435] = 12'hccc;
rom[118436] = 12'hccc;
rom[118437] = 12'hccc;
rom[118438] = 12'hccc;
rom[118439] = 12'hccc;
rom[118440] = 12'hccc;
rom[118441] = 12'hccc;
rom[118442] = 12'hccc;
rom[118443] = 12'hccc;
rom[118444] = 12'hccc;
rom[118445] = 12'hccc;
rom[118446] = 12'hccc;
rom[118447] = 12'hccc;
rom[118448] = 12'hccc;
rom[118449] = 12'hbbb;
rom[118450] = 12'hbbb;
rom[118451] = 12'hbbb;
rom[118452] = 12'hbbb;
rom[118453] = 12'hbbb;
rom[118454] = 12'hbbb;
rom[118455] = 12'hbbb;
rom[118456] = 12'hbbb;
rom[118457] = 12'hbbb;
rom[118458] = 12'hbbb;
rom[118459] = 12'hbbb;
rom[118460] = 12'hbbb;
rom[118461] = 12'hbbb;
rom[118462] = 12'hbbb;
rom[118463] = 12'hbbb;
rom[118464] = 12'hccc;
rom[118465] = 12'hbbb;
rom[118466] = 12'hbbb;
rom[118467] = 12'hbbb;
rom[118468] = 12'hbbb;
rom[118469] = 12'hbbb;
rom[118470] = 12'hbbb;
rom[118471] = 12'hbbb;
rom[118472] = 12'hccc;
rom[118473] = 12'heee;
rom[118474] = 12'hfff;
rom[118475] = 12'hfff;
rom[118476] = 12'hfff;
rom[118477] = 12'hddd;
rom[118478] = 12'hccc;
rom[118479] = 12'hbbb;
rom[118480] = 12'h999;
rom[118481] = 12'h999;
rom[118482] = 12'h999;
rom[118483] = 12'h999;
rom[118484] = 12'h999;
rom[118485] = 12'h999;
rom[118486] = 12'h888;
rom[118487] = 12'h888;
rom[118488] = 12'h888;
rom[118489] = 12'h888;
rom[118490] = 12'h888;
rom[118491] = 12'h888;
rom[118492] = 12'h999;
rom[118493] = 12'hbbb;
rom[118494] = 12'hbbb;
rom[118495] = 12'hbbb;
rom[118496] = 12'h999;
rom[118497] = 12'h888;
rom[118498] = 12'h888;
rom[118499] = 12'h888;
rom[118500] = 12'h777;
rom[118501] = 12'h888;
rom[118502] = 12'h888;
rom[118503] = 12'h777;
rom[118504] = 12'h666;
rom[118505] = 12'h777;
rom[118506] = 12'h777;
rom[118507] = 12'h777;
rom[118508] = 12'h666;
rom[118509] = 12'h666;
rom[118510] = 12'h555;
rom[118511] = 12'h555;
rom[118512] = 12'h555;
rom[118513] = 12'h555;
rom[118514] = 12'h555;
rom[118515] = 12'h555;
rom[118516] = 12'h555;
rom[118517] = 12'h555;
rom[118518] = 12'h555;
rom[118519] = 12'h666;
rom[118520] = 12'h666;
rom[118521] = 12'h666;
rom[118522] = 12'h666;
rom[118523] = 12'h666;
rom[118524] = 12'h666;
rom[118525] = 12'h666;
rom[118526] = 12'h666;
rom[118527] = 12'h666;
rom[118528] = 12'h555;
rom[118529] = 12'h555;
rom[118530] = 12'h444;
rom[118531] = 12'h444;
rom[118532] = 12'h444;
rom[118533] = 12'h555;
rom[118534] = 12'h555;
rom[118535] = 12'h444;
rom[118536] = 12'h444;
rom[118537] = 12'h444;
rom[118538] = 12'h444;
rom[118539] = 12'h333;
rom[118540] = 12'h333;
rom[118541] = 12'h333;
rom[118542] = 12'h333;
rom[118543] = 12'h333;
rom[118544] = 12'h444;
rom[118545] = 12'h444;
rom[118546] = 12'h444;
rom[118547] = 12'h333;
rom[118548] = 12'h333;
rom[118549] = 12'h333;
rom[118550] = 12'h333;
rom[118551] = 12'h333;
rom[118552] = 12'h444;
rom[118553] = 12'h444;
rom[118554] = 12'h444;
rom[118555] = 12'h444;
rom[118556] = 12'h444;
rom[118557] = 12'h444;
rom[118558] = 12'h444;
rom[118559] = 12'h444;
rom[118560] = 12'h444;
rom[118561] = 12'h444;
rom[118562] = 12'h444;
rom[118563] = 12'h333;
rom[118564] = 12'h333;
rom[118565] = 12'h444;
rom[118566] = 12'h444;
rom[118567] = 12'h444;
rom[118568] = 12'h555;
rom[118569] = 12'h555;
rom[118570] = 12'h444;
rom[118571] = 12'h444;
rom[118572] = 12'h444;
rom[118573] = 12'h444;
rom[118574] = 12'h444;
rom[118575] = 12'h333;
rom[118576] = 12'h333;
rom[118577] = 12'h333;
rom[118578] = 12'h333;
rom[118579] = 12'h444;
rom[118580] = 12'h555;
rom[118581] = 12'h444;
rom[118582] = 12'h333;
rom[118583] = 12'h333;
rom[118584] = 12'h333;
rom[118585] = 12'h333;
rom[118586] = 12'h333;
rom[118587] = 12'h333;
rom[118588] = 12'h222;
rom[118589] = 12'h333;
rom[118590] = 12'h333;
rom[118591] = 12'h444;
rom[118592] = 12'h666;
rom[118593] = 12'h555;
rom[118594] = 12'h555;
rom[118595] = 12'h444;
rom[118596] = 12'h444;
rom[118597] = 12'h444;
rom[118598] = 12'h333;
rom[118599] = 12'h222;
rom[118600] = 12'h333;
rom[118601] = 12'h222;
rom[118602] = 12'h222;
rom[118603] = 12'h222;
rom[118604] = 12'h333;
rom[118605] = 12'h333;
rom[118606] = 12'h333;
rom[118607] = 12'h333;
rom[118608] = 12'h333;
rom[118609] = 12'h222;
rom[118610] = 12'h222;
rom[118611] = 12'h222;
rom[118612] = 12'h222;
rom[118613] = 12'h333;
rom[118614] = 12'h333;
rom[118615] = 12'h333;
rom[118616] = 12'h222;
rom[118617] = 12'h111;
rom[118618] = 12'h222;
rom[118619] = 12'h222;
rom[118620] = 12'h222;
rom[118621] = 12'h111;
rom[118622] = 12'h  0;
rom[118623] = 12'h  0;
rom[118624] = 12'h  0;
rom[118625] = 12'h  0;
rom[118626] = 12'h  0;
rom[118627] = 12'h  0;
rom[118628] = 12'h111;
rom[118629] = 12'h444;
rom[118630] = 12'h555;
rom[118631] = 12'h555;
rom[118632] = 12'h222;
rom[118633] = 12'h  0;
rom[118634] = 12'h  0;
rom[118635] = 12'h111;
rom[118636] = 12'h333;
rom[118637] = 12'h555;
rom[118638] = 12'h666;
rom[118639] = 12'h888;
rom[118640] = 12'h666;
rom[118641] = 12'h333;
rom[118642] = 12'h  0;
rom[118643] = 12'h  0;
rom[118644] = 12'h  0;
rom[118645] = 12'h  0;
rom[118646] = 12'h  0;
rom[118647] = 12'h  0;
rom[118648] = 12'h  0;
rom[118649] = 12'h  0;
rom[118650] = 12'h  0;
rom[118651] = 12'h  0;
rom[118652] = 12'h  0;
rom[118653] = 12'h  0;
rom[118654] = 12'h  0;
rom[118655] = 12'h  0;
rom[118656] = 12'h  0;
rom[118657] = 12'h  0;
rom[118658] = 12'h  0;
rom[118659] = 12'h  0;
rom[118660] = 12'h  0;
rom[118661] = 12'h  0;
rom[118662] = 12'h  0;
rom[118663] = 12'h444;
rom[118664] = 12'hccc;
rom[118665] = 12'heee;
rom[118666] = 12'hbbb;
rom[118667] = 12'h444;
rom[118668] = 12'h111;
rom[118669] = 12'h111;
rom[118670] = 12'h111;
rom[118671] = 12'h111;
rom[118672] = 12'h  0;
rom[118673] = 12'h  0;
rom[118674] = 12'h  0;
rom[118675] = 12'h  0;
rom[118676] = 12'h222;
rom[118677] = 12'h777;
rom[118678] = 12'haaa;
rom[118679] = 12'haaa;
rom[118680] = 12'h333;
rom[118681] = 12'h111;
rom[118682] = 12'h  0;
rom[118683] = 12'h  0;
rom[118684] = 12'h  0;
rom[118685] = 12'h111;
rom[118686] = 12'h111;
rom[118687] = 12'h  0;
rom[118688] = 12'h111;
rom[118689] = 12'h  0;
rom[118690] = 12'h111;
rom[118691] = 12'h333;
rom[118692] = 12'h555;
rom[118693] = 12'h444;
rom[118694] = 12'h222;
rom[118695] = 12'h  0;
rom[118696] = 12'h333;
rom[118697] = 12'h555;
rom[118698] = 12'h666;
rom[118699] = 12'h555;
rom[118700] = 12'h222;
rom[118701] = 12'h  0;
rom[118702] = 12'h  0;
rom[118703] = 12'h111;
rom[118704] = 12'h111;
rom[118705] = 12'h  0;
rom[118706] = 12'h  0;
rom[118707] = 12'h  0;
rom[118708] = 12'h  0;
rom[118709] = 12'h  0;
rom[118710] = 12'h  0;
rom[118711] = 12'h  0;
rom[118712] = 12'h111;
rom[118713] = 12'h111;
rom[118714] = 12'h111;
rom[118715] = 12'h222;
rom[118716] = 12'h444;
rom[118717] = 12'h555;
rom[118718] = 12'h777;
rom[118719] = 12'h888;
rom[118720] = 12'h777;
rom[118721] = 12'h555;
rom[118722] = 12'h333;
rom[118723] = 12'h111;
rom[118724] = 12'h  0;
rom[118725] = 12'h  0;
rom[118726] = 12'h  0;
rom[118727] = 12'h  0;
rom[118728] = 12'h  0;
rom[118729] = 12'h  0;
rom[118730] = 12'h  0;
rom[118731] = 12'h  0;
rom[118732] = 12'h  0;
rom[118733] = 12'h  0;
rom[118734] = 12'h  0;
rom[118735] = 12'h  0;
rom[118736] = 12'h  0;
rom[118737] = 12'h  0;
rom[118738] = 12'h  0;
rom[118739] = 12'h  0;
rom[118740] = 12'h  0;
rom[118741] = 12'h  0;
rom[118742] = 12'h  0;
rom[118743] = 12'h  0;
rom[118744] = 12'h  0;
rom[118745] = 12'h  0;
rom[118746] = 12'h  0;
rom[118747] = 12'h  0;
rom[118748] = 12'h  0;
rom[118749] = 12'h  0;
rom[118750] = 12'h  0;
rom[118751] = 12'h  0;
rom[118752] = 12'h  0;
rom[118753] = 12'h  0;
rom[118754] = 12'h  0;
rom[118755] = 12'h  0;
rom[118756] = 12'h  0;
rom[118757] = 12'h  0;
rom[118758] = 12'h  0;
rom[118759] = 12'h  0;
rom[118760] = 12'h  0;
rom[118761] = 12'h  0;
rom[118762] = 12'h  0;
rom[118763] = 12'h  0;
rom[118764] = 12'h  0;
rom[118765] = 12'h  0;
rom[118766] = 12'h  0;
rom[118767] = 12'h  0;
rom[118768] = 12'h  0;
rom[118769] = 12'h  0;
rom[118770] = 12'h  0;
rom[118771] = 12'h111;
rom[118772] = 12'h222;
rom[118773] = 12'h444;
rom[118774] = 12'h777;
rom[118775] = 12'h999;
rom[118776] = 12'h888;
rom[118777] = 12'h555;
rom[118778] = 12'h222;
rom[118779] = 12'h111;
rom[118780] = 12'h111;
rom[118781] = 12'h  0;
rom[118782] = 12'h  0;
rom[118783] = 12'h  0;
rom[118784] = 12'h  0;
rom[118785] = 12'h  0;
rom[118786] = 12'h  0;
rom[118787] = 12'h  0;
rom[118788] = 12'h  0;
rom[118789] = 12'h  0;
rom[118790] = 12'h  0;
rom[118791] = 12'h  0;
rom[118792] = 12'h  0;
rom[118793] = 12'h  0;
rom[118794] = 12'h  0;
rom[118795] = 12'h  0;
rom[118796] = 12'h  0;
rom[118797] = 12'h  0;
rom[118798] = 12'h  0;
rom[118799] = 12'h  0;
rom[118800] = 12'hfff;
rom[118801] = 12'hfff;
rom[118802] = 12'heee;
rom[118803] = 12'heee;
rom[118804] = 12'heee;
rom[118805] = 12'heee;
rom[118806] = 12'heee;
rom[118807] = 12'heee;
rom[118808] = 12'heee;
rom[118809] = 12'heee;
rom[118810] = 12'heee;
rom[118811] = 12'heee;
rom[118812] = 12'heee;
rom[118813] = 12'heee;
rom[118814] = 12'heee;
rom[118815] = 12'heee;
rom[118816] = 12'heee;
rom[118817] = 12'heee;
rom[118818] = 12'hddd;
rom[118819] = 12'hddd;
rom[118820] = 12'hddd;
rom[118821] = 12'hddd;
rom[118822] = 12'hddd;
rom[118823] = 12'hddd;
rom[118824] = 12'hddd;
rom[118825] = 12'hddd;
rom[118826] = 12'hddd;
rom[118827] = 12'hddd;
rom[118828] = 12'hddd;
rom[118829] = 12'hddd;
rom[118830] = 12'hddd;
rom[118831] = 12'hddd;
rom[118832] = 12'hddd;
rom[118833] = 12'hddd;
rom[118834] = 12'hccc;
rom[118835] = 12'hccc;
rom[118836] = 12'hccc;
rom[118837] = 12'hccc;
rom[118838] = 12'hccc;
rom[118839] = 12'hccc;
rom[118840] = 12'hccc;
rom[118841] = 12'hccc;
rom[118842] = 12'hccc;
rom[118843] = 12'hccc;
rom[118844] = 12'hccc;
rom[118845] = 12'hccc;
rom[118846] = 12'hccc;
rom[118847] = 12'hccc;
rom[118848] = 12'hbbb;
rom[118849] = 12'hbbb;
rom[118850] = 12'hbbb;
rom[118851] = 12'hbbb;
rom[118852] = 12'hbbb;
rom[118853] = 12'hbbb;
rom[118854] = 12'hbbb;
rom[118855] = 12'hbbb;
rom[118856] = 12'hbbb;
rom[118857] = 12'hbbb;
rom[118858] = 12'hbbb;
rom[118859] = 12'hbbb;
rom[118860] = 12'hbbb;
rom[118861] = 12'hbbb;
rom[118862] = 12'hbbb;
rom[118863] = 12'hbbb;
rom[118864] = 12'hbbb;
rom[118865] = 12'hbbb;
rom[118866] = 12'hbbb;
rom[118867] = 12'hbbb;
rom[118868] = 12'hbbb;
rom[118869] = 12'hbbb;
rom[118870] = 12'hbbb;
rom[118871] = 12'hbbb;
rom[118872] = 12'hddd;
rom[118873] = 12'heee;
rom[118874] = 12'hfff;
rom[118875] = 12'hfff;
rom[118876] = 12'heee;
rom[118877] = 12'hccc;
rom[118878] = 12'hbbb;
rom[118879] = 12'haaa;
rom[118880] = 12'h999;
rom[118881] = 12'h999;
rom[118882] = 12'h999;
rom[118883] = 12'h999;
rom[118884] = 12'h888;
rom[118885] = 12'h888;
rom[118886] = 12'h888;
rom[118887] = 12'h888;
rom[118888] = 12'h888;
rom[118889] = 12'h777;
rom[118890] = 12'h777;
rom[118891] = 12'h888;
rom[118892] = 12'haaa;
rom[118893] = 12'hbbb;
rom[118894] = 12'hbbb;
rom[118895] = 12'haaa;
rom[118896] = 12'h888;
rom[118897] = 12'h777;
rom[118898] = 12'h888;
rom[118899] = 12'h888;
rom[118900] = 12'h777;
rom[118901] = 12'h777;
rom[118902] = 12'h888;
rom[118903] = 12'h777;
rom[118904] = 12'h666;
rom[118905] = 12'h666;
rom[118906] = 12'h777;
rom[118907] = 12'h777;
rom[118908] = 12'h666;
rom[118909] = 12'h666;
rom[118910] = 12'h555;
rom[118911] = 12'h555;
rom[118912] = 12'h555;
rom[118913] = 12'h555;
rom[118914] = 12'h555;
rom[118915] = 12'h555;
rom[118916] = 12'h555;
rom[118917] = 12'h555;
rom[118918] = 12'h555;
rom[118919] = 12'h666;
rom[118920] = 12'h666;
rom[118921] = 12'h666;
rom[118922] = 12'h666;
rom[118923] = 12'h666;
rom[118924] = 12'h666;
rom[118925] = 12'h666;
rom[118926] = 12'h666;
rom[118927] = 12'h666;
rom[118928] = 12'h555;
rom[118929] = 12'h444;
rom[118930] = 12'h444;
rom[118931] = 12'h444;
rom[118932] = 12'h444;
rom[118933] = 12'h555;
rom[118934] = 12'h555;
rom[118935] = 12'h444;
rom[118936] = 12'h444;
rom[118937] = 12'h444;
rom[118938] = 12'h333;
rom[118939] = 12'h333;
rom[118940] = 12'h333;
rom[118941] = 12'h333;
rom[118942] = 12'h333;
rom[118943] = 12'h333;
rom[118944] = 12'h333;
rom[118945] = 12'h444;
rom[118946] = 12'h444;
rom[118947] = 12'h333;
rom[118948] = 12'h333;
rom[118949] = 12'h333;
rom[118950] = 12'h333;
rom[118951] = 12'h333;
rom[118952] = 12'h333;
rom[118953] = 12'h444;
rom[118954] = 12'h444;
rom[118955] = 12'h444;
rom[118956] = 12'h444;
rom[118957] = 12'h444;
rom[118958] = 12'h444;
rom[118959] = 12'h444;
rom[118960] = 12'h444;
rom[118961] = 12'h444;
rom[118962] = 12'h333;
rom[118963] = 12'h333;
rom[118964] = 12'h333;
rom[118965] = 12'h333;
rom[118966] = 12'h444;
rom[118967] = 12'h444;
rom[118968] = 12'h444;
rom[118969] = 12'h444;
rom[118970] = 12'h444;
rom[118971] = 12'h444;
rom[118972] = 12'h444;
rom[118973] = 12'h444;
rom[118974] = 12'h333;
rom[118975] = 12'h333;
rom[118976] = 12'h333;
rom[118977] = 12'h333;
rom[118978] = 12'h333;
rom[118979] = 12'h444;
rom[118980] = 12'h444;
rom[118981] = 12'h444;
rom[118982] = 12'h333;
rom[118983] = 12'h333;
rom[118984] = 12'h333;
rom[118985] = 12'h333;
rom[118986] = 12'h333;
rom[118987] = 12'h222;
rom[118988] = 12'h222;
rom[118989] = 12'h222;
rom[118990] = 12'h333;
rom[118991] = 12'h333;
rom[118992] = 12'h555;
rom[118993] = 12'h555;
rom[118994] = 12'h555;
rom[118995] = 12'h444;
rom[118996] = 12'h444;
rom[118997] = 12'h333;
rom[118998] = 12'h333;
rom[118999] = 12'h222;
rom[119000] = 12'h222;
rom[119001] = 12'h222;
rom[119002] = 12'h222;
rom[119003] = 12'h222;
rom[119004] = 12'h222;
rom[119005] = 12'h222;
rom[119006] = 12'h222;
rom[119007] = 12'h222;
rom[119008] = 12'h222;
rom[119009] = 12'h222;
rom[119010] = 12'h111;
rom[119011] = 12'h111;
rom[119012] = 12'h222;
rom[119013] = 12'h222;
rom[119014] = 12'h333;
rom[119015] = 12'h333;
rom[119016] = 12'h222;
rom[119017] = 12'h111;
rom[119018] = 12'h111;
rom[119019] = 12'h222;
rom[119020] = 12'h222;
rom[119021] = 12'h111;
rom[119022] = 12'h  0;
rom[119023] = 12'h  0;
rom[119024] = 12'h  0;
rom[119025] = 12'h  0;
rom[119026] = 12'h  0;
rom[119027] = 12'h  0;
rom[119028] = 12'h  0;
rom[119029] = 12'h222;
rom[119030] = 12'h444;
rom[119031] = 12'h555;
rom[119032] = 12'h333;
rom[119033] = 12'h111;
rom[119034] = 12'h111;
rom[119035] = 12'h111;
rom[119036] = 12'h333;
rom[119037] = 12'h555;
rom[119038] = 12'h666;
rom[119039] = 12'h777;
rom[119040] = 12'h444;
rom[119041] = 12'h222;
rom[119042] = 12'h  0;
rom[119043] = 12'h  0;
rom[119044] = 12'h  0;
rom[119045] = 12'h  0;
rom[119046] = 12'h  0;
rom[119047] = 12'h  0;
rom[119048] = 12'h  0;
rom[119049] = 12'h  0;
rom[119050] = 12'h  0;
rom[119051] = 12'h  0;
rom[119052] = 12'h  0;
rom[119053] = 12'h  0;
rom[119054] = 12'h  0;
rom[119055] = 12'h  0;
rom[119056] = 12'h  0;
rom[119057] = 12'h  0;
rom[119058] = 12'h  0;
rom[119059] = 12'h  0;
rom[119060] = 12'h  0;
rom[119061] = 12'h  0;
rom[119062] = 12'h  0;
rom[119063] = 12'h444;
rom[119064] = 12'hccc;
rom[119065] = 12'heee;
rom[119066] = 12'hbbb;
rom[119067] = 12'h444;
rom[119068] = 12'h111;
rom[119069] = 12'h111;
rom[119070] = 12'h111;
rom[119071] = 12'h111;
rom[119072] = 12'h  0;
rom[119073] = 12'h  0;
rom[119074] = 12'h  0;
rom[119075] = 12'h  0;
rom[119076] = 12'h222;
rom[119077] = 12'h777;
rom[119078] = 12'haaa;
rom[119079] = 12'haaa;
rom[119080] = 12'h444;
rom[119081] = 12'h111;
rom[119082] = 12'h  0;
rom[119083] = 12'h  0;
rom[119084] = 12'h  0;
rom[119085] = 12'h  0;
rom[119086] = 12'h  0;
rom[119087] = 12'h  0;
rom[119088] = 12'h111;
rom[119089] = 12'h  0;
rom[119090] = 12'h111;
rom[119091] = 12'h333;
rom[119092] = 12'h444;
rom[119093] = 12'h444;
rom[119094] = 12'h222;
rom[119095] = 12'h  0;
rom[119096] = 12'h111;
rom[119097] = 12'h333;
rom[119098] = 12'h555;
rom[119099] = 12'h555;
rom[119100] = 12'h444;
rom[119101] = 12'h111;
rom[119102] = 12'h  0;
rom[119103] = 12'h  0;
rom[119104] = 12'h  0;
rom[119105] = 12'h  0;
rom[119106] = 12'h  0;
rom[119107] = 12'h  0;
rom[119108] = 12'h  0;
rom[119109] = 12'h  0;
rom[119110] = 12'h  0;
rom[119111] = 12'h  0;
rom[119112] = 12'h  0;
rom[119113] = 12'h  0;
rom[119114] = 12'h111;
rom[119115] = 12'h222;
rom[119116] = 12'h333;
rom[119117] = 12'h444;
rom[119118] = 12'h666;
rom[119119] = 12'h888;
rom[119120] = 12'h777;
rom[119121] = 12'h555;
rom[119122] = 12'h333;
rom[119123] = 12'h111;
rom[119124] = 12'h  0;
rom[119125] = 12'h  0;
rom[119126] = 12'h  0;
rom[119127] = 12'h  0;
rom[119128] = 12'h  0;
rom[119129] = 12'h  0;
rom[119130] = 12'h  0;
rom[119131] = 12'h  0;
rom[119132] = 12'h  0;
rom[119133] = 12'h  0;
rom[119134] = 12'h  0;
rom[119135] = 12'h  0;
rom[119136] = 12'h  0;
rom[119137] = 12'h  0;
rom[119138] = 12'h  0;
rom[119139] = 12'h  0;
rom[119140] = 12'h  0;
rom[119141] = 12'h  0;
rom[119142] = 12'h  0;
rom[119143] = 12'h  0;
rom[119144] = 12'h  0;
rom[119145] = 12'h  0;
rom[119146] = 12'h  0;
rom[119147] = 12'h  0;
rom[119148] = 12'h  0;
rom[119149] = 12'h  0;
rom[119150] = 12'h  0;
rom[119151] = 12'h  0;
rom[119152] = 12'h  0;
rom[119153] = 12'h  0;
rom[119154] = 12'h  0;
rom[119155] = 12'h  0;
rom[119156] = 12'h  0;
rom[119157] = 12'h  0;
rom[119158] = 12'h  0;
rom[119159] = 12'h  0;
rom[119160] = 12'h  0;
rom[119161] = 12'h  0;
rom[119162] = 12'h  0;
rom[119163] = 12'h  0;
rom[119164] = 12'h  0;
rom[119165] = 12'h  0;
rom[119166] = 12'h  0;
rom[119167] = 12'h  0;
rom[119168] = 12'h  0;
rom[119169] = 12'h  0;
rom[119170] = 12'h  0;
rom[119171] = 12'h111;
rom[119172] = 12'h222;
rom[119173] = 12'h333;
rom[119174] = 12'h666;
rom[119175] = 12'h888;
rom[119176] = 12'h888;
rom[119177] = 12'h555;
rom[119178] = 12'h222;
rom[119179] = 12'h111;
rom[119180] = 12'h111;
rom[119181] = 12'h  0;
rom[119182] = 12'h  0;
rom[119183] = 12'h  0;
rom[119184] = 12'h  0;
rom[119185] = 12'h  0;
rom[119186] = 12'h  0;
rom[119187] = 12'h  0;
rom[119188] = 12'h  0;
rom[119189] = 12'h  0;
rom[119190] = 12'h  0;
rom[119191] = 12'h  0;
rom[119192] = 12'h  0;
rom[119193] = 12'h  0;
rom[119194] = 12'h  0;
rom[119195] = 12'h  0;
rom[119196] = 12'h  0;
rom[119197] = 12'h  0;
rom[119198] = 12'h  0;
rom[119199] = 12'h  0;
rom[119200] = 12'hfff;
rom[119201] = 12'heee;
rom[119202] = 12'heee;
rom[119203] = 12'heee;
rom[119204] = 12'heee;
rom[119205] = 12'heee;
rom[119206] = 12'heee;
rom[119207] = 12'heee;
rom[119208] = 12'heee;
rom[119209] = 12'heee;
rom[119210] = 12'heee;
rom[119211] = 12'heee;
rom[119212] = 12'heee;
rom[119213] = 12'heee;
rom[119214] = 12'heee;
rom[119215] = 12'heee;
rom[119216] = 12'heee;
rom[119217] = 12'heee;
rom[119218] = 12'hddd;
rom[119219] = 12'hddd;
rom[119220] = 12'hddd;
rom[119221] = 12'hddd;
rom[119222] = 12'hddd;
rom[119223] = 12'hddd;
rom[119224] = 12'hddd;
rom[119225] = 12'hddd;
rom[119226] = 12'hddd;
rom[119227] = 12'hddd;
rom[119228] = 12'hddd;
rom[119229] = 12'hddd;
rom[119230] = 12'hddd;
rom[119231] = 12'hddd;
rom[119232] = 12'hccc;
rom[119233] = 12'hccc;
rom[119234] = 12'hccc;
rom[119235] = 12'hccc;
rom[119236] = 12'hccc;
rom[119237] = 12'hccc;
rom[119238] = 12'hccc;
rom[119239] = 12'hccc;
rom[119240] = 12'hccc;
rom[119241] = 12'hccc;
rom[119242] = 12'hccc;
rom[119243] = 12'hccc;
rom[119244] = 12'hccc;
rom[119245] = 12'hccc;
rom[119246] = 12'hccc;
rom[119247] = 12'hbbb;
rom[119248] = 12'hbbb;
rom[119249] = 12'hbbb;
rom[119250] = 12'hbbb;
rom[119251] = 12'hbbb;
rom[119252] = 12'hbbb;
rom[119253] = 12'hbbb;
rom[119254] = 12'hbbb;
rom[119255] = 12'hbbb;
rom[119256] = 12'hbbb;
rom[119257] = 12'hbbb;
rom[119258] = 12'hbbb;
rom[119259] = 12'hbbb;
rom[119260] = 12'hbbb;
rom[119261] = 12'hbbb;
rom[119262] = 12'hbbb;
rom[119263] = 12'hbbb;
rom[119264] = 12'hbbb;
rom[119265] = 12'hbbb;
rom[119266] = 12'hbbb;
rom[119267] = 12'hbbb;
rom[119268] = 12'hbbb;
rom[119269] = 12'haaa;
rom[119270] = 12'hbbb;
rom[119271] = 12'hccc;
rom[119272] = 12'heee;
rom[119273] = 12'hfff;
rom[119274] = 12'hfff;
rom[119275] = 12'heee;
rom[119276] = 12'hddd;
rom[119277] = 12'hbbb;
rom[119278] = 12'haaa;
rom[119279] = 12'h999;
rom[119280] = 12'h999;
rom[119281] = 12'h999;
rom[119282] = 12'h888;
rom[119283] = 12'h888;
rom[119284] = 12'h888;
rom[119285] = 12'h888;
rom[119286] = 12'h777;
rom[119287] = 12'h777;
rom[119288] = 12'h777;
rom[119289] = 12'h666;
rom[119290] = 12'h666;
rom[119291] = 12'h888;
rom[119292] = 12'hbbb;
rom[119293] = 12'hccc;
rom[119294] = 12'haaa;
rom[119295] = 12'h888;
rom[119296] = 12'h777;
rom[119297] = 12'h777;
rom[119298] = 12'h888;
rom[119299] = 12'h888;
rom[119300] = 12'h777;
rom[119301] = 12'h777;
rom[119302] = 12'h777;
rom[119303] = 12'h777;
rom[119304] = 12'h666;
rom[119305] = 12'h666;
rom[119306] = 12'h666;
rom[119307] = 12'h666;
rom[119308] = 12'h666;
rom[119309] = 12'h666;
rom[119310] = 12'h555;
rom[119311] = 12'h555;
rom[119312] = 12'h555;
rom[119313] = 12'h555;
rom[119314] = 12'h555;
rom[119315] = 12'h555;
rom[119316] = 12'h444;
rom[119317] = 12'h444;
rom[119318] = 12'h555;
rom[119319] = 12'h666;
rom[119320] = 12'h666;
rom[119321] = 12'h666;
rom[119322] = 12'h555;
rom[119323] = 12'h555;
rom[119324] = 12'h666;
rom[119325] = 12'h666;
rom[119326] = 12'h666;
rom[119327] = 12'h555;
rom[119328] = 12'h444;
rom[119329] = 12'h444;
rom[119330] = 12'h444;
rom[119331] = 12'h444;
rom[119332] = 12'h555;
rom[119333] = 12'h555;
rom[119334] = 12'h555;
rom[119335] = 12'h444;
rom[119336] = 12'h333;
rom[119337] = 12'h333;
rom[119338] = 12'h333;
rom[119339] = 12'h333;
rom[119340] = 12'h333;
rom[119341] = 12'h333;
rom[119342] = 12'h333;
rom[119343] = 12'h333;
rom[119344] = 12'h333;
rom[119345] = 12'h333;
rom[119346] = 12'h333;
rom[119347] = 12'h333;
rom[119348] = 12'h333;
rom[119349] = 12'h333;
rom[119350] = 12'h333;
rom[119351] = 12'h333;
rom[119352] = 12'h333;
rom[119353] = 12'h444;
rom[119354] = 12'h444;
rom[119355] = 12'h444;
rom[119356] = 12'h444;
rom[119357] = 12'h444;
rom[119358] = 12'h333;
rom[119359] = 12'h333;
rom[119360] = 12'h333;
rom[119361] = 12'h333;
rom[119362] = 12'h333;
rom[119363] = 12'h333;
rom[119364] = 12'h333;
rom[119365] = 12'h333;
rom[119366] = 12'h444;
rom[119367] = 12'h444;
rom[119368] = 12'h444;
rom[119369] = 12'h444;
rom[119370] = 12'h444;
rom[119371] = 12'h333;
rom[119372] = 12'h333;
rom[119373] = 12'h333;
rom[119374] = 12'h333;
rom[119375] = 12'h222;
rom[119376] = 12'h222;
rom[119377] = 12'h222;
rom[119378] = 12'h333;
rom[119379] = 12'h333;
rom[119380] = 12'h444;
rom[119381] = 12'h333;
rom[119382] = 12'h333;
rom[119383] = 12'h222;
rom[119384] = 12'h222;
rom[119385] = 12'h222;
rom[119386] = 12'h222;
rom[119387] = 12'h222;
rom[119388] = 12'h222;
rom[119389] = 12'h222;
rom[119390] = 12'h222;
rom[119391] = 12'h333;
rom[119392] = 12'h555;
rom[119393] = 12'h555;
rom[119394] = 12'h444;
rom[119395] = 12'h444;
rom[119396] = 12'h333;
rom[119397] = 12'h333;
rom[119398] = 12'h222;
rom[119399] = 12'h222;
rom[119400] = 12'h222;
rom[119401] = 12'h111;
rom[119402] = 12'h111;
rom[119403] = 12'h111;
rom[119404] = 12'h222;
rom[119405] = 12'h222;
rom[119406] = 12'h222;
rom[119407] = 12'h222;
rom[119408] = 12'h222;
rom[119409] = 12'h111;
rom[119410] = 12'h111;
rom[119411] = 12'h111;
rom[119412] = 12'h111;
rom[119413] = 12'h222;
rom[119414] = 12'h222;
rom[119415] = 12'h222;
rom[119416] = 12'h111;
rom[119417] = 12'h111;
rom[119418] = 12'h  0;
rom[119419] = 12'h111;
rom[119420] = 12'h222;
rom[119421] = 12'h111;
rom[119422] = 12'h  0;
rom[119423] = 12'h  0;
rom[119424] = 12'h  0;
rom[119425] = 12'h  0;
rom[119426] = 12'h  0;
rom[119427] = 12'h  0;
rom[119428] = 12'h  0;
rom[119429] = 12'h  0;
rom[119430] = 12'h222;
rom[119431] = 12'h444;
rom[119432] = 12'h444;
rom[119433] = 12'h333;
rom[119434] = 12'h222;
rom[119435] = 12'h222;
rom[119436] = 12'h444;
rom[119437] = 12'h666;
rom[119438] = 12'h666;
rom[119439] = 12'h666;
rom[119440] = 12'h222;
rom[119441] = 12'h  0;
rom[119442] = 12'h  0;
rom[119443] = 12'h  0;
rom[119444] = 12'h  0;
rom[119445] = 12'h  0;
rom[119446] = 12'h  0;
rom[119447] = 12'h  0;
rom[119448] = 12'h  0;
rom[119449] = 12'h  0;
rom[119450] = 12'h  0;
rom[119451] = 12'h  0;
rom[119452] = 12'h  0;
rom[119453] = 12'h  0;
rom[119454] = 12'h  0;
rom[119455] = 12'h  0;
rom[119456] = 12'h  0;
rom[119457] = 12'h  0;
rom[119458] = 12'h  0;
rom[119459] = 12'h  0;
rom[119460] = 12'h  0;
rom[119461] = 12'h  0;
rom[119462] = 12'h111;
rom[119463] = 12'h555;
rom[119464] = 12'hddd;
rom[119465] = 12'heee;
rom[119466] = 12'haaa;
rom[119467] = 12'h333;
rom[119468] = 12'h111;
rom[119469] = 12'h111;
rom[119470] = 12'h  0;
rom[119471] = 12'h  0;
rom[119472] = 12'h  0;
rom[119473] = 12'h  0;
rom[119474] = 12'h  0;
rom[119475] = 12'h  0;
rom[119476] = 12'h111;
rom[119477] = 12'h666;
rom[119478] = 12'haaa;
rom[119479] = 12'haaa;
rom[119480] = 12'h555;
rom[119481] = 12'h222;
rom[119482] = 12'h  0;
rom[119483] = 12'h  0;
rom[119484] = 12'h  0;
rom[119485] = 12'h  0;
rom[119486] = 12'h  0;
rom[119487] = 12'h  0;
rom[119488] = 12'h111;
rom[119489] = 12'h  0;
rom[119490] = 12'h111;
rom[119491] = 12'h222;
rom[119492] = 12'h444;
rom[119493] = 12'h444;
rom[119494] = 12'h222;
rom[119495] = 12'h111;
rom[119496] = 12'h111;
rom[119497] = 12'h222;
rom[119498] = 12'h444;
rom[119499] = 12'h555;
rom[119500] = 12'h555;
rom[119501] = 12'h222;
rom[119502] = 12'h  0;
rom[119503] = 12'h  0;
rom[119504] = 12'h  0;
rom[119505] = 12'h  0;
rom[119506] = 12'h  0;
rom[119507] = 12'h  0;
rom[119508] = 12'h  0;
rom[119509] = 12'h  0;
rom[119510] = 12'h  0;
rom[119511] = 12'h  0;
rom[119512] = 12'h  0;
rom[119513] = 12'h  0;
rom[119514] = 12'h111;
rom[119515] = 12'h111;
rom[119516] = 12'h222;
rom[119517] = 12'h333;
rom[119518] = 12'h666;
rom[119519] = 12'h888;
rom[119520] = 12'h888;
rom[119521] = 12'h666;
rom[119522] = 12'h333;
rom[119523] = 12'h111;
rom[119524] = 12'h111;
rom[119525] = 12'h  0;
rom[119526] = 12'h  0;
rom[119527] = 12'h  0;
rom[119528] = 12'h  0;
rom[119529] = 12'h  0;
rom[119530] = 12'h  0;
rom[119531] = 12'h  0;
rom[119532] = 12'h  0;
rom[119533] = 12'h  0;
rom[119534] = 12'h  0;
rom[119535] = 12'h  0;
rom[119536] = 12'h  0;
rom[119537] = 12'h  0;
rom[119538] = 12'h  0;
rom[119539] = 12'h  0;
rom[119540] = 12'h  0;
rom[119541] = 12'h  0;
rom[119542] = 12'h  0;
rom[119543] = 12'h  0;
rom[119544] = 12'h  0;
rom[119545] = 12'h  0;
rom[119546] = 12'h  0;
rom[119547] = 12'h  0;
rom[119548] = 12'h  0;
rom[119549] = 12'h  0;
rom[119550] = 12'h  0;
rom[119551] = 12'h  0;
rom[119552] = 12'h  0;
rom[119553] = 12'h  0;
rom[119554] = 12'h  0;
rom[119555] = 12'h  0;
rom[119556] = 12'h  0;
rom[119557] = 12'h  0;
rom[119558] = 12'h  0;
rom[119559] = 12'h  0;
rom[119560] = 12'h  0;
rom[119561] = 12'h  0;
rom[119562] = 12'h  0;
rom[119563] = 12'h  0;
rom[119564] = 12'h  0;
rom[119565] = 12'h  0;
rom[119566] = 12'h  0;
rom[119567] = 12'h  0;
rom[119568] = 12'h  0;
rom[119569] = 12'h  0;
rom[119570] = 12'h  0;
rom[119571] = 12'h111;
rom[119572] = 12'h111;
rom[119573] = 12'h222;
rom[119574] = 12'h444;
rom[119575] = 12'h666;
rom[119576] = 12'h888;
rom[119577] = 12'h666;
rom[119578] = 12'h333;
rom[119579] = 12'h111;
rom[119580] = 12'h  0;
rom[119581] = 12'h  0;
rom[119582] = 12'h  0;
rom[119583] = 12'h  0;
rom[119584] = 12'h  0;
rom[119585] = 12'h  0;
rom[119586] = 12'h  0;
rom[119587] = 12'h  0;
rom[119588] = 12'h  0;
rom[119589] = 12'h  0;
rom[119590] = 12'h  0;
rom[119591] = 12'h  0;
rom[119592] = 12'h  0;
rom[119593] = 12'h  0;
rom[119594] = 12'h  0;
rom[119595] = 12'h  0;
rom[119596] = 12'h  0;
rom[119597] = 12'h  0;
rom[119598] = 12'h  0;
rom[119599] = 12'h  0;
rom[119600] = 12'heee;
rom[119601] = 12'heee;
rom[119602] = 12'heee;
rom[119603] = 12'heee;
rom[119604] = 12'heee;
rom[119605] = 12'heee;
rom[119606] = 12'heee;
rom[119607] = 12'heee;
rom[119608] = 12'heee;
rom[119609] = 12'heee;
rom[119610] = 12'heee;
rom[119611] = 12'heee;
rom[119612] = 12'heee;
rom[119613] = 12'heee;
rom[119614] = 12'hddd;
rom[119615] = 12'hddd;
rom[119616] = 12'hddd;
rom[119617] = 12'hddd;
rom[119618] = 12'hddd;
rom[119619] = 12'hddd;
rom[119620] = 12'hddd;
rom[119621] = 12'hddd;
rom[119622] = 12'hddd;
rom[119623] = 12'hddd;
rom[119624] = 12'hddd;
rom[119625] = 12'hddd;
rom[119626] = 12'hddd;
rom[119627] = 12'hddd;
rom[119628] = 12'hddd;
rom[119629] = 12'hccc;
rom[119630] = 12'hccc;
rom[119631] = 12'hccc;
rom[119632] = 12'hccc;
rom[119633] = 12'hccc;
rom[119634] = 12'hccc;
rom[119635] = 12'hccc;
rom[119636] = 12'hccc;
rom[119637] = 12'hccc;
rom[119638] = 12'hccc;
rom[119639] = 12'hccc;
rom[119640] = 12'hccc;
rom[119641] = 12'hccc;
rom[119642] = 12'hccc;
rom[119643] = 12'hccc;
rom[119644] = 12'hccc;
rom[119645] = 12'hccc;
rom[119646] = 12'hbbb;
rom[119647] = 12'hbbb;
rom[119648] = 12'hbbb;
rom[119649] = 12'hbbb;
rom[119650] = 12'hbbb;
rom[119651] = 12'hbbb;
rom[119652] = 12'hbbb;
rom[119653] = 12'hbbb;
rom[119654] = 12'hbbb;
rom[119655] = 12'hbbb;
rom[119656] = 12'hbbb;
rom[119657] = 12'hbbb;
rom[119658] = 12'hbbb;
rom[119659] = 12'hbbb;
rom[119660] = 12'hbbb;
rom[119661] = 12'hbbb;
rom[119662] = 12'hbbb;
rom[119663] = 12'hbbb;
rom[119664] = 12'haaa;
rom[119665] = 12'hbbb;
rom[119666] = 12'hbbb;
rom[119667] = 12'hbbb;
rom[119668] = 12'haaa;
rom[119669] = 12'hbbb;
rom[119670] = 12'hccc;
rom[119671] = 12'hddd;
rom[119672] = 12'hfff;
rom[119673] = 12'hfff;
rom[119674] = 12'heee;
rom[119675] = 12'hddd;
rom[119676] = 12'hbbb;
rom[119677] = 12'haaa;
rom[119678] = 12'h999;
rom[119679] = 12'h999;
rom[119680] = 12'h999;
rom[119681] = 12'h888;
rom[119682] = 12'h888;
rom[119683] = 12'h777;
rom[119684] = 12'h777;
rom[119685] = 12'h777;
rom[119686] = 12'h777;
rom[119687] = 12'h777;
rom[119688] = 12'h777;
rom[119689] = 12'h666;
rom[119690] = 12'h777;
rom[119691] = 12'h999;
rom[119692] = 12'hbbb;
rom[119693] = 12'hbbb;
rom[119694] = 12'h999;
rom[119695] = 12'h777;
rom[119696] = 12'h666;
rom[119697] = 12'h666;
rom[119698] = 12'h777;
rom[119699] = 12'h888;
rom[119700] = 12'h777;
rom[119701] = 12'h777;
rom[119702] = 12'h777;
rom[119703] = 12'h666;
rom[119704] = 12'h666;
rom[119705] = 12'h666;
rom[119706] = 12'h666;
rom[119707] = 12'h666;
rom[119708] = 12'h666;
rom[119709] = 12'h666;
rom[119710] = 12'h555;
rom[119711] = 12'h555;
rom[119712] = 12'h444;
rom[119713] = 12'h555;
rom[119714] = 12'h555;
rom[119715] = 12'h555;
rom[119716] = 12'h444;
rom[119717] = 12'h444;
rom[119718] = 12'h555;
rom[119719] = 12'h666;
rom[119720] = 12'h666;
rom[119721] = 12'h666;
rom[119722] = 12'h555;
rom[119723] = 12'h555;
rom[119724] = 12'h555;
rom[119725] = 12'h555;
rom[119726] = 12'h555;
rom[119727] = 12'h555;
rom[119728] = 12'h444;
rom[119729] = 12'h444;
rom[119730] = 12'h444;
rom[119731] = 12'h444;
rom[119732] = 12'h555;
rom[119733] = 12'h555;
rom[119734] = 12'h555;
rom[119735] = 12'h444;
rom[119736] = 12'h333;
rom[119737] = 12'h333;
rom[119738] = 12'h333;
rom[119739] = 12'h333;
rom[119740] = 12'h333;
rom[119741] = 12'h333;
rom[119742] = 12'h333;
rom[119743] = 12'h333;
rom[119744] = 12'h333;
rom[119745] = 12'h333;
rom[119746] = 12'h333;
rom[119747] = 12'h333;
rom[119748] = 12'h333;
rom[119749] = 12'h333;
rom[119750] = 12'h333;
rom[119751] = 12'h333;
rom[119752] = 12'h333;
rom[119753] = 12'h333;
rom[119754] = 12'h444;
rom[119755] = 12'h444;
rom[119756] = 12'h444;
rom[119757] = 12'h333;
rom[119758] = 12'h333;
rom[119759] = 12'h333;
rom[119760] = 12'h333;
rom[119761] = 12'h333;
rom[119762] = 12'h333;
rom[119763] = 12'h333;
rom[119764] = 12'h333;
rom[119765] = 12'h333;
rom[119766] = 12'h444;
rom[119767] = 12'h444;
rom[119768] = 12'h444;
rom[119769] = 12'h444;
rom[119770] = 12'h333;
rom[119771] = 12'h333;
rom[119772] = 12'h333;
rom[119773] = 12'h333;
rom[119774] = 12'h222;
rom[119775] = 12'h222;
rom[119776] = 12'h222;
rom[119777] = 12'h222;
rom[119778] = 12'h222;
rom[119779] = 12'h333;
rom[119780] = 12'h333;
rom[119781] = 12'h333;
rom[119782] = 12'h333;
rom[119783] = 12'h222;
rom[119784] = 12'h222;
rom[119785] = 12'h222;
rom[119786] = 12'h222;
rom[119787] = 12'h222;
rom[119788] = 12'h222;
rom[119789] = 12'h222;
rom[119790] = 12'h222;
rom[119791] = 12'h222;
rom[119792] = 12'h444;
rom[119793] = 12'h444;
rom[119794] = 12'h444;
rom[119795] = 12'h444;
rom[119796] = 12'h333;
rom[119797] = 12'h222;
rom[119798] = 12'h222;
rom[119799] = 12'h222;
rom[119800] = 12'h111;
rom[119801] = 12'h111;
rom[119802] = 12'h111;
rom[119803] = 12'h111;
rom[119804] = 12'h111;
rom[119805] = 12'h111;
rom[119806] = 12'h111;
rom[119807] = 12'h111;
rom[119808] = 12'h111;
rom[119809] = 12'h111;
rom[119810] = 12'h111;
rom[119811] = 12'h111;
rom[119812] = 12'h111;
rom[119813] = 12'h111;
rom[119814] = 12'h222;
rom[119815] = 12'h222;
rom[119816] = 12'h222;
rom[119817] = 12'h111;
rom[119818] = 12'h  0;
rom[119819] = 12'h111;
rom[119820] = 12'h222;
rom[119821] = 12'h111;
rom[119822] = 12'h  0;
rom[119823] = 12'h  0;
rom[119824] = 12'h  0;
rom[119825] = 12'h  0;
rom[119826] = 12'h  0;
rom[119827] = 12'h  0;
rom[119828] = 12'h  0;
rom[119829] = 12'h  0;
rom[119830] = 12'h111;
rom[119831] = 12'h333;
rom[119832] = 12'h444;
rom[119833] = 12'h333;
rom[119834] = 12'h222;
rom[119835] = 12'h222;
rom[119836] = 12'h444;
rom[119837] = 12'h666;
rom[119838] = 12'h666;
rom[119839] = 12'h444;
rom[119840] = 12'h111;
rom[119841] = 12'h  0;
rom[119842] = 12'h  0;
rom[119843] = 12'h  0;
rom[119844] = 12'h  0;
rom[119845] = 12'h  0;
rom[119846] = 12'h  0;
rom[119847] = 12'h  0;
rom[119848] = 12'h  0;
rom[119849] = 12'h  0;
rom[119850] = 12'h  0;
rom[119851] = 12'h  0;
rom[119852] = 12'h  0;
rom[119853] = 12'h  0;
rom[119854] = 12'h  0;
rom[119855] = 12'h  0;
rom[119856] = 12'h  0;
rom[119857] = 12'h  0;
rom[119858] = 12'h  0;
rom[119859] = 12'h  0;
rom[119860] = 12'h  0;
rom[119861] = 12'h  0;
rom[119862] = 12'h111;
rom[119863] = 12'h555;
rom[119864] = 12'heee;
rom[119865] = 12'heee;
rom[119866] = 12'haaa;
rom[119867] = 12'h333;
rom[119868] = 12'h111;
rom[119869] = 12'h111;
rom[119870] = 12'h  0;
rom[119871] = 12'h  0;
rom[119872] = 12'h  0;
rom[119873] = 12'h  0;
rom[119874] = 12'h  0;
rom[119875] = 12'h  0;
rom[119876] = 12'h111;
rom[119877] = 12'h555;
rom[119878] = 12'h999;
rom[119879] = 12'hbbb;
rom[119880] = 12'h666;
rom[119881] = 12'h222;
rom[119882] = 12'h  0;
rom[119883] = 12'h  0;
rom[119884] = 12'h  0;
rom[119885] = 12'h  0;
rom[119886] = 12'h111;
rom[119887] = 12'h  0;
rom[119888] = 12'h  0;
rom[119889] = 12'h  0;
rom[119890] = 12'h  0;
rom[119891] = 12'h222;
rom[119892] = 12'h444;
rom[119893] = 12'h444;
rom[119894] = 12'h222;
rom[119895] = 12'h111;
rom[119896] = 12'h111;
rom[119897] = 12'h111;
rom[119898] = 12'h222;
rom[119899] = 12'h444;
rom[119900] = 12'h555;
rom[119901] = 12'h333;
rom[119902] = 12'h111;
rom[119903] = 12'h  0;
rom[119904] = 12'h  0;
rom[119905] = 12'h  0;
rom[119906] = 12'h  0;
rom[119907] = 12'h  0;
rom[119908] = 12'h  0;
rom[119909] = 12'h  0;
rom[119910] = 12'h  0;
rom[119911] = 12'h  0;
rom[119912] = 12'h  0;
rom[119913] = 12'h  0;
rom[119914] = 12'h111;
rom[119915] = 12'h111;
rom[119916] = 12'h111;
rom[119917] = 12'h222;
rom[119918] = 12'h555;
rom[119919] = 12'h777;
rom[119920] = 12'h888;
rom[119921] = 12'h666;
rom[119922] = 12'h333;
rom[119923] = 12'h222;
rom[119924] = 12'h111;
rom[119925] = 12'h  0;
rom[119926] = 12'h  0;
rom[119927] = 12'h  0;
rom[119928] = 12'h  0;
rom[119929] = 12'h  0;
rom[119930] = 12'h  0;
rom[119931] = 12'h  0;
rom[119932] = 12'h  0;
rom[119933] = 12'h  0;
rom[119934] = 12'h  0;
rom[119935] = 12'h  0;
rom[119936] = 12'h  0;
rom[119937] = 12'h  0;
rom[119938] = 12'h  0;
rom[119939] = 12'h  0;
rom[119940] = 12'h  0;
rom[119941] = 12'h  0;
rom[119942] = 12'h  0;
rom[119943] = 12'h  0;
rom[119944] = 12'h  0;
rom[119945] = 12'h  0;
rom[119946] = 12'h  0;
rom[119947] = 12'h  0;
rom[119948] = 12'h  0;
rom[119949] = 12'h  0;
rom[119950] = 12'h  0;
rom[119951] = 12'h  0;
rom[119952] = 12'h  0;
rom[119953] = 12'h  0;
rom[119954] = 12'h  0;
rom[119955] = 12'h  0;
rom[119956] = 12'h  0;
rom[119957] = 12'h  0;
rom[119958] = 12'h  0;
rom[119959] = 12'h  0;
rom[119960] = 12'h  0;
rom[119961] = 12'h  0;
rom[119962] = 12'h  0;
rom[119963] = 12'h  0;
rom[119964] = 12'h  0;
rom[119965] = 12'h  0;
rom[119966] = 12'h  0;
rom[119967] = 12'h  0;
rom[119968] = 12'h  0;
rom[119969] = 12'h  0;
rom[119970] = 12'h  0;
rom[119971] = 12'h  0;
rom[119972] = 12'h  0;
rom[119973] = 12'h111;
rom[119974] = 12'h333;
rom[119975] = 12'h555;
rom[119976] = 12'h777;
rom[119977] = 12'h666;
rom[119978] = 12'h444;
rom[119979] = 12'h222;
rom[119980] = 12'h111;
rom[119981] = 12'h111;
rom[119982] = 12'h  0;
rom[119983] = 12'h  0;
rom[119984] = 12'h  0;
rom[119985] = 12'h  0;
rom[119986] = 12'h  0;
rom[119987] = 12'h  0;
rom[119988] = 12'h  0;
rom[119989] = 12'h  0;
rom[119990] = 12'h  0;
rom[119991] = 12'h  0;
rom[119992] = 12'h  0;
rom[119993] = 12'h  0;
rom[119994] = 12'h  0;
rom[119995] = 12'h  0;
rom[119996] = 12'h  0;
rom[119997] = 12'h  0;
rom[119998] = 12'h  0;
rom[119999] = 12'h  0;
rom[120000] = 12'heee;
rom[120001] = 12'heee;
rom[120002] = 12'heee;
rom[120003] = 12'heee;
rom[120004] = 12'heee;
rom[120005] = 12'hddd;
rom[120006] = 12'hddd;
rom[120007] = 12'hddd;
rom[120008] = 12'hddd;
rom[120009] = 12'hddd;
rom[120010] = 12'hddd;
rom[120011] = 12'hddd;
rom[120012] = 12'hddd;
rom[120013] = 12'hddd;
rom[120014] = 12'hddd;
rom[120015] = 12'hddd;
rom[120016] = 12'hddd;
rom[120017] = 12'hddd;
rom[120018] = 12'hddd;
rom[120019] = 12'hddd;
rom[120020] = 12'hddd;
rom[120021] = 12'hddd;
rom[120022] = 12'hddd;
rom[120023] = 12'hddd;
rom[120024] = 12'hccc;
rom[120025] = 12'hccc;
rom[120026] = 12'hccc;
rom[120027] = 12'hccc;
rom[120028] = 12'hccc;
rom[120029] = 12'hccc;
rom[120030] = 12'hccc;
rom[120031] = 12'hccc;
rom[120032] = 12'hccc;
rom[120033] = 12'hccc;
rom[120034] = 12'hccc;
rom[120035] = 12'hccc;
rom[120036] = 12'hccc;
rom[120037] = 12'hccc;
rom[120038] = 12'hccc;
rom[120039] = 12'hccc;
rom[120040] = 12'hccc;
rom[120041] = 12'hccc;
rom[120042] = 12'hccc;
rom[120043] = 12'hccc;
rom[120044] = 12'hccc;
rom[120045] = 12'hccc;
rom[120046] = 12'hbbb;
rom[120047] = 12'hbbb;
rom[120048] = 12'hbbb;
rom[120049] = 12'hbbb;
rom[120050] = 12'hbbb;
rom[120051] = 12'hbbb;
rom[120052] = 12'hbbb;
rom[120053] = 12'hbbb;
rom[120054] = 12'hbbb;
rom[120055] = 12'hbbb;
rom[120056] = 12'hbbb;
rom[120057] = 12'hbbb;
rom[120058] = 12'hbbb;
rom[120059] = 12'hbbb;
rom[120060] = 12'hbbb;
rom[120061] = 12'hbbb;
rom[120062] = 12'haaa;
rom[120063] = 12'haaa;
rom[120064] = 12'haaa;
rom[120065] = 12'haaa;
rom[120066] = 12'hbbb;
rom[120067] = 12'haaa;
rom[120068] = 12'hbbb;
rom[120069] = 12'hccc;
rom[120070] = 12'hddd;
rom[120071] = 12'hfff;
rom[120072] = 12'hfff;
rom[120073] = 12'hfff;
rom[120074] = 12'hddd;
rom[120075] = 12'hccc;
rom[120076] = 12'haaa;
rom[120077] = 12'h999;
rom[120078] = 12'h999;
rom[120079] = 12'h999;
rom[120080] = 12'h999;
rom[120081] = 12'h888;
rom[120082] = 12'h888;
rom[120083] = 12'h777;
rom[120084] = 12'h777;
rom[120085] = 12'h777;
rom[120086] = 12'h777;
rom[120087] = 12'h666;
rom[120088] = 12'h666;
rom[120089] = 12'h777;
rom[120090] = 12'h999;
rom[120091] = 12'hbbb;
rom[120092] = 12'hbbb;
rom[120093] = 12'haaa;
rom[120094] = 12'h888;
rom[120095] = 12'h666;
rom[120096] = 12'h777;
rom[120097] = 12'h666;
rom[120098] = 12'h777;
rom[120099] = 12'h777;
rom[120100] = 12'h777;
rom[120101] = 12'h777;
rom[120102] = 12'h777;
rom[120103] = 12'h777;
rom[120104] = 12'h666;
rom[120105] = 12'h666;
rom[120106] = 12'h666;
rom[120107] = 12'h666;
rom[120108] = 12'h666;
rom[120109] = 12'h666;
rom[120110] = 12'h555;
rom[120111] = 12'h555;
rom[120112] = 12'h444;
rom[120113] = 12'h444;
rom[120114] = 12'h555;
rom[120115] = 12'h555;
rom[120116] = 12'h444;
rom[120117] = 12'h444;
rom[120118] = 12'h555;
rom[120119] = 12'h666;
rom[120120] = 12'h666;
rom[120121] = 12'h666;
rom[120122] = 12'h555;
rom[120123] = 12'h555;
rom[120124] = 12'h555;
rom[120125] = 12'h555;
rom[120126] = 12'h555;
rom[120127] = 12'h555;
rom[120128] = 12'h444;
rom[120129] = 12'h444;
rom[120130] = 12'h444;
rom[120131] = 12'h444;
rom[120132] = 12'h444;
rom[120133] = 12'h555;
rom[120134] = 12'h444;
rom[120135] = 12'h444;
rom[120136] = 12'h333;
rom[120137] = 12'h333;
rom[120138] = 12'h333;
rom[120139] = 12'h333;
rom[120140] = 12'h333;
rom[120141] = 12'h333;
rom[120142] = 12'h333;
rom[120143] = 12'h333;
rom[120144] = 12'h333;
rom[120145] = 12'h333;
rom[120146] = 12'h333;
rom[120147] = 12'h333;
rom[120148] = 12'h333;
rom[120149] = 12'h333;
rom[120150] = 12'h333;
rom[120151] = 12'h333;
rom[120152] = 12'h333;
rom[120153] = 12'h333;
rom[120154] = 12'h333;
rom[120155] = 12'h333;
rom[120156] = 12'h333;
rom[120157] = 12'h333;
rom[120158] = 12'h333;
rom[120159] = 12'h333;
rom[120160] = 12'h333;
rom[120161] = 12'h333;
rom[120162] = 12'h333;
rom[120163] = 12'h333;
rom[120164] = 12'h333;
rom[120165] = 12'h333;
rom[120166] = 12'h444;
rom[120167] = 12'h444;
rom[120168] = 12'h333;
rom[120169] = 12'h333;
rom[120170] = 12'h333;
rom[120171] = 12'h333;
rom[120172] = 12'h333;
rom[120173] = 12'h222;
rom[120174] = 12'h222;
rom[120175] = 12'h222;
rom[120176] = 12'h222;
rom[120177] = 12'h222;
rom[120178] = 12'h222;
rom[120179] = 12'h222;
rom[120180] = 12'h333;
rom[120181] = 12'h333;
rom[120182] = 12'h333;
rom[120183] = 12'h222;
rom[120184] = 12'h111;
rom[120185] = 12'h222;
rom[120186] = 12'h222;
rom[120187] = 12'h222;
rom[120188] = 12'h222;
rom[120189] = 12'h222;
rom[120190] = 12'h222;
rom[120191] = 12'h222;
rom[120192] = 12'h333;
rom[120193] = 12'h444;
rom[120194] = 12'h444;
rom[120195] = 12'h444;
rom[120196] = 12'h333;
rom[120197] = 12'h222;
rom[120198] = 12'h111;
rom[120199] = 12'h111;
rom[120200] = 12'h111;
rom[120201] = 12'h111;
rom[120202] = 12'h111;
rom[120203] = 12'h111;
rom[120204] = 12'h111;
rom[120205] = 12'h111;
rom[120206] = 12'h111;
rom[120207] = 12'h111;
rom[120208] = 12'h111;
rom[120209] = 12'h111;
rom[120210] = 12'h111;
rom[120211] = 12'h111;
rom[120212] = 12'h  0;
rom[120213] = 12'h111;
rom[120214] = 12'h111;
rom[120215] = 12'h222;
rom[120216] = 12'h222;
rom[120217] = 12'h111;
rom[120218] = 12'h  0;
rom[120219] = 12'h111;
rom[120220] = 12'h111;
rom[120221] = 12'h111;
rom[120222] = 12'h  0;
rom[120223] = 12'h  0;
rom[120224] = 12'h  0;
rom[120225] = 12'h  0;
rom[120226] = 12'h  0;
rom[120227] = 12'h  0;
rom[120228] = 12'h  0;
rom[120229] = 12'h  0;
rom[120230] = 12'h  0;
rom[120231] = 12'h111;
rom[120232] = 12'h333;
rom[120233] = 12'h333;
rom[120234] = 12'h333;
rom[120235] = 12'h222;
rom[120236] = 12'h444;
rom[120237] = 12'h666;
rom[120238] = 12'h555;
rom[120239] = 12'h333;
rom[120240] = 12'h111;
rom[120241] = 12'h  0;
rom[120242] = 12'h  0;
rom[120243] = 12'h  0;
rom[120244] = 12'h  0;
rom[120245] = 12'h  0;
rom[120246] = 12'h  0;
rom[120247] = 12'h  0;
rom[120248] = 12'h  0;
rom[120249] = 12'h  0;
rom[120250] = 12'h  0;
rom[120251] = 12'h  0;
rom[120252] = 12'h  0;
rom[120253] = 12'h  0;
rom[120254] = 12'h  0;
rom[120255] = 12'h  0;
rom[120256] = 12'h  0;
rom[120257] = 12'h  0;
rom[120258] = 12'h  0;
rom[120259] = 12'h  0;
rom[120260] = 12'h  0;
rom[120261] = 12'h  0;
rom[120262] = 12'h111;
rom[120263] = 12'h666;
rom[120264] = 12'heee;
rom[120265] = 12'heee;
rom[120266] = 12'h999;
rom[120267] = 12'h333;
rom[120268] = 12'h111;
rom[120269] = 12'h111;
rom[120270] = 12'h  0;
rom[120271] = 12'h  0;
rom[120272] = 12'h  0;
rom[120273] = 12'h  0;
rom[120274] = 12'h  0;
rom[120275] = 12'h  0;
rom[120276] = 12'h  0;
rom[120277] = 12'h444;
rom[120278] = 12'h888;
rom[120279] = 12'hbbb;
rom[120280] = 12'h666;
rom[120281] = 12'h333;
rom[120282] = 12'h  0;
rom[120283] = 12'h  0;
rom[120284] = 12'h  0;
rom[120285] = 12'h  0;
rom[120286] = 12'h111;
rom[120287] = 12'h  0;
rom[120288] = 12'h  0;
rom[120289] = 12'h  0;
rom[120290] = 12'h  0;
rom[120291] = 12'h111;
rom[120292] = 12'h333;
rom[120293] = 12'h444;
rom[120294] = 12'h222;
rom[120295] = 12'h111;
rom[120296] = 12'h111;
rom[120297] = 12'h111;
rom[120298] = 12'h111;
rom[120299] = 12'h333;
rom[120300] = 12'h444;
rom[120301] = 12'h333;
rom[120302] = 12'h222;
rom[120303] = 12'h  0;
rom[120304] = 12'h  0;
rom[120305] = 12'h  0;
rom[120306] = 12'h  0;
rom[120307] = 12'h  0;
rom[120308] = 12'h  0;
rom[120309] = 12'h  0;
rom[120310] = 12'h  0;
rom[120311] = 12'h  0;
rom[120312] = 12'h  0;
rom[120313] = 12'h  0;
rom[120314] = 12'h111;
rom[120315] = 12'h111;
rom[120316] = 12'h111;
rom[120317] = 12'h222;
rom[120318] = 12'h444;
rom[120319] = 12'h666;
rom[120320] = 12'h888;
rom[120321] = 12'h666;
rom[120322] = 12'h444;
rom[120323] = 12'h333;
rom[120324] = 12'h111;
rom[120325] = 12'h  0;
rom[120326] = 12'h  0;
rom[120327] = 12'h  0;
rom[120328] = 12'h  0;
rom[120329] = 12'h  0;
rom[120330] = 12'h  0;
rom[120331] = 12'h  0;
rom[120332] = 12'h  0;
rom[120333] = 12'h  0;
rom[120334] = 12'h  0;
rom[120335] = 12'h  0;
rom[120336] = 12'h  0;
rom[120337] = 12'h  0;
rom[120338] = 12'h  0;
rom[120339] = 12'h  0;
rom[120340] = 12'h  0;
rom[120341] = 12'h  0;
rom[120342] = 12'h  0;
rom[120343] = 12'h  0;
rom[120344] = 12'h  0;
rom[120345] = 12'h  0;
rom[120346] = 12'h  0;
rom[120347] = 12'h  0;
rom[120348] = 12'h  0;
rom[120349] = 12'h  0;
rom[120350] = 12'h  0;
rom[120351] = 12'h  0;
rom[120352] = 12'h  0;
rom[120353] = 12'h  0;
rom[120354] = 12'h  0;
rom[120355] = 12'h  0;
rom[120356] = 12'h  0;
rom[120357] = 12'h  0;
rom[120358] = 12'h  0;
rom[120359] = 12'h  0;
rom[120360] = 12'h  0;
rom[120361] = 12'h  0;
rom[120362] = 12'h  0;
rom[120363] = 12'h  0;
rom[120364] = 12'h  0;
rom[120365] = 12'h  0;
rom[120366] = 12'h  0;
rom[120367] = 12'h  0;
rom[120368] = 12'h  0;
rom[120369] = 12'h  0;
rom[120370] = 12'h  0;
rom[120371] = 12'h  0;
rom[120372] = 12'h  0;
rom[120373] = 12'h111;
rom[120374] = 12'h222;
rom[120375] = 12'h444;
rom[120376] = 12'h777;
rom[120377] = 12'h777;
rom[120378] = 12'h666;
rom[120379] = 12'h333;
rom[120380] = 12'h111;
rom[120381] = 12'h111;
rom[120382] = 12'h  0;
rom[120383] = 12'h  0;
rom[120384] = 12'h  0;
rom[120385] = 12'h  0;
rom[120386] = 12'h  0;
rom[120387] = 12'h  0;
rom[120388] = 12'h  0;
rom[120389] = 12'h  0;
rom[120390] = 12'h  0;
rom[120391] = 12'h  0;
rom[120392] = 12'h  0;
rom[120393] = 12'h  0;
rom[120394] = 12'h  0;
rom[120395] = 12'h  0;
rom[120396] = 12'h  0;
rom[120397] = 12'h  0;
rom[120398] = 12'h  0;
rom[120399] = 12'h  0;
rom[120400] = 12'heee;
rom[120401] = 12'heee;
rom[120402] = 12'heee;
rom[120403] = 12'heee;
rom[120404] = 12'hddd;
rom[120405] = 12'hddd;
rom[120406] = 12'hddd;
rom[120407] = 12'hddd;
rom[120408] = 12'hddd;
rom[120409] = 12'hddd;
rom[120410] = 12'hddd;
rom[120411] = 12'hddd;
rom[120412] = 12'hddd;
rom[120413] = 12'hddd;
rom[120414] = 12'hddd;
rom[120415] = 12'hddd;
rom[120416] = 12'hddd;
rom[120417] = 12'hddd;
rom[120418] = 12'hddd;
rom[120419] = 12'hddd;
rom[120420] = 12'hddd;
rom[120421] = 12'hddd;
rom[120422] = 12'hddd;
rom[120423] = 12'hddd;
rom[120424] = 12'hccc;
rom[120425] = 12'hccc;
rom[120426] = 12'hccc;
rom[120427] = 12'hccc;
rom[120428] = 12'hccc;
rom[120429] = 12'hccc;
rom[120430] = 12'hccc;
rom[120431] = 12'hccc;
rom[120432] = 12'hccc;
rom[120433] = 12'hccc;
rom[120434] = 12'hccc;
rom[120435] = 12'hccc;
rom[120436] = 12'hccc;
rom[120437] = 12'hccc;
rom[120438] = 12'hccc;
rom[120439] = 12'hccc;
rom[120440] = 12'hccc;
rom[120441] = 12'hccc;
rom[120442] = 12'hccc;
rom[120443] = 12'hccc;
rom[120444] = 12'hccc;
rom[120445] = 12'hbbb;
rom[120446] = 12'hbbb;
rom[120447] = 12'hbbb;
rom[120448] = 12'hbbb;
rom[120449] = 12'hbbb;
rom[120450] = 12'hbbb;
rom[120451] = 12'hbbb;
rom[120452] = 12'hbbb;
rom[120453] = 12'hbbb;
rom[120454] = 12'hbbb;
rom[120455] = 12'hbbb;
rom[120456] = 12'haaa;
rom[120457] = 12'haaa;
rom[120458] = 12'hbbb;
rom[120459] = 12'hbbb;
rom[120460] = 12'haaa;
rom[120461] = 12'haaa;
rom[120462] = 12'haaa;
rom[120463] = 12'haaa;
rom[120464] = 12'haaa;
rom[120465] = 12'haaa;
rom[120466] = 12'haaa;
rom[120467] = 12'haaa;
rom[120468] = 12'hbbb;
rom[120469] = 12'hddd;
rom[120470] = 12'heee;
rom[120471] = 12'hfff;
rom[120472] = 12'hfff;
rom[120473] = 12'heee;
rom[120474] = 12'hccc;
rom[120475] = 12'haaa;
rom[120476] = 12'h999;
rom[120477] = 12'h888;
rom[120478] = 12'h888;
rom[120479] = 12'h888;
rom[120480] = 12'h888;
rom[120481] = 12'h888;
rom[120482] = 12'h888;
rom[120483] = 12'h777;
rom[120484] = 12'h777;
rom[120485] = 12'h777;
rom[120486] = 12'h666;
rom[120487] = 12'h666;
rom[120488] = 12'h666;
rom[120489] = 12'h888;
rom[120490] = 12'haaa;
rom[120491] = 12'hbbb;
rom[120492] = 12'haaa;
rom[120493] = 12'h888;
rom[120494] = 12'h777;
rom[120495] = 12'h666;
rom[120496] = 12'h777;
rom[120497] = 12'h666;
rom[120498] = 12'h666;
rom[120499] = 12'h666;
rom[120500] = 12'h777;
rom[120501] = 12'h777;
rom[120502] = 12'h777;
rom[120503] = 12'h777;
rom[120504] = 12'h666;
rom[120505] = 12'h666;
rom[120506] = 12'h666;
rom[120507] = 12'h666;
rom[120508] = 12'h666;
rom[120509] = 12'h666;
rom[120510] = 12'h555;
rom[120511] = 12'h555;
rom[120512] = 12'h444;
rom[120513] = 12'h444;
rom[120514] = 12'h444;
rom[120515] = 12'h444;
rom[120516] = 12'h444;
rom[120517] = 12'h444;
rom[120518] = 12'h555;
rom[120519] = 12'h666;
rom[120520] = 12'h666;
rom[120521] = 12'h666;
rom[120522] = 12'h555;
rom[120523] = 12'h555;
rom[120524] = 12'h555;
rom[120525] = 12'h555;
rom[120526] = 12'h555;
rom[120527] = 12'h555;
rom[120528] = 12'h555;
rom[120529] = 12'h555;
rom[120530] = 12'h444;
rom[120531] = 12'h444;
rom[120532] = 12'h444;
rom[120533] = 12'h555;
rom[120534] = 12'h444;
rom[120535] = 12'h444;
rom[120536] = 12'h333;
rom[120537] = 12'h333;
rom[120538] = 12'h333;
rom[120539] = 12'h333;
rom[120540] = 12'h333;
rom[120541] = 12'h333;
rom[120542] = 12'h333;
rom[120543] = 12'h333;
rom[120544] = 12'h333;
rom[120545] = 12'h333;
rom[120546] = 12'h333;
rom[120547] = 12'h333;
rom[120548] = 12'h333;
rom[120549] = 12'h333;
rom[120550] = 12'h333;
rom[120551] = 12'h333;
rom[120552] = 12'h333;
rom[120553] = 12'h333;
rom[120554] = 12'h333;
rom[120555] = 12'h333;
rom[120556] = 12'h333;
rom[120557] = 12'h333;
rom[120558] = 12'h333;
rom[120559] = 12'h333;
rom[120560] = 12'h333;
rom[120561] = 12'h333;
rom[120562] = 12'h333;
rom[120563] = 12'h333;
rom[120564] = 12'h333;
rom[120565] = 12'h333;
rom[120566] = 12'h333;
rom[120567] = 12'h333;
rom[120568] = 12'h333;
rom[120569] = 12'h333;
rom[120570] = 12'h333;
rom[120571] = 12'h222;
rom[120572] = 12'h222;
rom[120573] = 12'h222;
rom[120574] = 12'h222;
rom[120575] = 12'h111;
rom[120576] = 12'h111;
rom[120577] = 12'h111;
rom[120578] = 12'h222;
rom[120579] = 12'h222;
rom[120580] = 12'h222;
rom[120581] = 12'h333;
rom[120582] = 12'h222;
rom[120583] = 12'h222;
rom[120584] = 12'h111;
rom[120585] = 12'h111;
rom[120586] = 12'h111;
rom[120587] = 12'h111;
rom[120588] = 12'h111;
rom[120589] = 12'h222;
rom[120590] = 12'h222;
rom[120591] = 12'h222;
rom[120592] = 12'h333;
rom[120593] = 12'h333;
rom[120594] = 12'h333;
rom[120595] = 12'h333;
rom[120596] = 12'h222;
rom[120597] = 12'h222;
rom[120598] = 12'h111;
rom[120599] = 12'h111;
rom[120600] = 12'h111;
rom[120601] = 12'h111;
rom[120602] = 12'h111;
rom[120603] = 12'h111;
rom[120604] = 12'h111;
rom[120605] = 12'h111;
rom[120606] = 12'h111;
rom[120607] = 12'h111;
rom[120608] = 12'h111;
rom[120609] = 12'h111;
rom[120610] = 12'h111;
rom[120611] = 12'h  0;
rom[120612] = 12'h  0;
rom[120613] = 12'h  0;
rom[120614] = 12'h111;
rom[120615] = 12'h111;
rom[120616] = 12'h111;
rom[120617] = 12'h111;
rom[120618] = 12'h  0;
rom[120619] = 12'h111;
rom[120620] = 12'h111;
rom[120621] = 12'h111;
rom[120622] = 12'h  0;
rom[120623] = 12'h  0;
rom[120624] = 12'h  0;
rom[120625] = 12'h  0;
rom[120626] = 12'h  0;
rom[120627] = 12'h  0;
rom[120628] = 12'h  0;
rom[120629] = 12'h  0;
rom[120630] = 12'h  0;
rom[120631] = 12'h  0;
rom[120632] = 12'h333;
rom[120633] = 12'h333;
rom[120634] = 12'h333;
rom[120635] = 12'h333;
rom[120636] = 12'h444;
rom[120637] = 12'h555;
rom[120638] = 12'h444;
rom[120639] = 12'h222;
rom[120640] = 12'h  0;
rom[120641] = 12'h  0;
rom[120642] = 12'h  0;
rom[120643] = 12'h  0;
rom[120644] = 12'h  0;
rom[120645] = 12'h  0;
rom[120646] = 12'h  0;
rom[120647] = 12'h  0;
rom[120648] = 12'h  0;
rom[120649] = 12'h  0;
rom[120650] = 12'h  0;
rom[120651] = 12'h  0;
rom[120652] = 12'h  0;
rom[120653] = 12'h  0;
rom[120654] = 12'h  0;
rom[120655] = 12'h  0;
rom[120656] = 12'h  0;
rom[120657] = 12'h  0;
rom[120658] = 12'h  0;
rom[120659] = 12'h  0;
rom[120660] = 12'h  0;
rom[120661] = 12'h  0;
rom[120662] = 12'h222;
rom[120663] = 12'h666;
rom[120664] = 12'heee;
rom[120665] = 12'heee;
rom[120666] = 12'h888;
rom[120667] = 12'h222;
rom[120668] = 12'h111;
rom[120669] = 12'h111;
rom[120670] = 12'h  0;
rom[120671] = 12'h  0;
rom[120672] = 12'h  0;
rom[120673] = 12'h  0;
rom[120674] = 12'h  0;
rom[120675] = 12'h  0;
rom[120676] = 12'h  0;
rom[120677] = 12'h333;
rom[120678] = 12'h888;
rom[120679] = 12'hbbb;
rom[120680] = 12'h777;
rom[120681] = 12'h333;
rom[120682] = 12'h  0;
rom[120683] = 12'h  0;
rom[120684] = 12'h  0;
rom[120685] = 12'h  0;
rom[120686] = 12'h111;
rom[120687] = 12'h  0;
rom[120688] = 12'h  0;
rom[120689] = 12'h  0;
rom[120690] = 12'h  0;
rom[120691] = 12'h111;
rom[120692] = 12'h333;
rom[120693] = 12'h333;
rom[120694] = 12'h222;
rom[120695] = 12'h111;
rom[120696] = 12'h111;
rom[120697] = 12'h  0;
rom[120698] = 12'h111;
rom[120699] = 12'h222;
rom[120700] = 12'h444;
rom[120701] = 12'h444;
rom[120702] = 12'h222;
rom[120703] = 12'h111;
rom[120704] = 12'h  0;
rom[120705] = 12'h  0;
rom[120706] = 12'h  0;
rom[120707] = 12'h  0;
rom[120708] = 12'h  0;
rom[120709] = 12'h  0;
rom[120710] = 12'h  0;
rom[120711] = 12'h  0;
rom[120712] = 12'h  0;
rom[120713] = 12'h  0;
rom[120714] = 12'h111;
rom[120715] = 12'h111;
rom[120716] = 12'h111;
rom[120717] = 12'h111;
rom[120718] = 12'h333;
rom[120719] = 12'h444;
rom[120720] = 12'h777;
rom[120721] = 12'h666;
rom[120722] = 12'h555;
rom[120723] = 12'h333;
rom[120724] = 12'h111;
rom[120725] = 12'h  0;
rom[120726] = 12'h  0;
rom[120727] = 12'h  0;
rom[120728] = 12'h  0;
rom[120729] = 12'h  0;
rom[120730] = 12'h  0;
rom[120731] = 12'h  0;
rom[120732] = 12'h  0;
rom[120733] = 12'h  0;
rom[120734] = 12'h  0;
rom[120735] = 12'h  0;
rom[120736] = 12'h  0;
rom[120737] = 12'h  0;
rom[120738] = 12'h  0;
rom[120739] = 12'h  0;
rom[120740] = 12'h  0;
rom[120741] = 12'h  0;
rom[120742] = 12'h  0;
rom[120743] = 12'h  0;
rom[120744] = 12'h  0;
rom[120745] = 12'h  0;
rom[120746] = 12'h  0;
rom[120747] = 12'h  0;
rom[120748] = 12'h  0;
rom[120749] = 12'h  0;
rom[120750] = 12'h  0;
rom[120751] = 12'h  0;
rom[120752] = 12'h  0;
rom[120753] = 12'h  0;
rom[120754] = 12'h  0;
rom[120755] = 12'h  0;
rom[120756] = 12'h  0;
rom[120757] = 12'h  0;
rom[120758] = 12'h  0;
rom[120759] = 12'h  0;
rom[120760] = 12'h  0;
rom[120761] = 12'h  0;
rom[120762] = 12'h  0;
rom[120763] = 12'h  0;
rom[120764] = 12'h  0;
rom[120765] = 12'h  0;
rom[120766] = 12'h  0;
rom[120767] = 12'h  0;
rom[120768] = 12'h  0;
rom[120769] = 12'h  0;
rom[120770] = 12'h  0;
rom[120771] = 12'h  0;
rom[120772] = 12'h  0;
rom[120773] = 12'h111;
rom[120774] = 12'h222;
rom[120775] = 12'h333;
rom[120776] = 12'h666;
rom[120777] = 12'h777;
rom[120778] = 12'h666;
rom[120779] = 12'h444;
rom[120780] = 12'h222;
rom[120781] = 12'h  0;
rom[120782] = 12'h  0;
rom[120783] = 12'h  0;
rom[120784] = 12'h  0;
rom[120785] = 12'h  0;
rom[120786] = 12'h  0;
rom[120787] = 12'h  0;
rom[120788] = 12'h  0;
rom[120789] = 12'h  0;
rom[120790] = 12'h  0;
rom[120791] = 12'h  0;
rom[120792] = 12'h  0;
rom[120793] = 12'h  0;
rom[120794] = 12'h  0;
rom[120795] = 12'h  0;
rom[120796] = 12'h  0;
rom[120797] = 12'h  0;
rom[120798] = 12'h  0;
rom[120799] = 12'h  0;
rom[120800] = 12'heee;
rom[120801] = 12'heee;
rom[120802] = 12'heee;
rom[120803] = 12'heee;
rom[120804] = 12'hddd;
rom[120805] = 12'hddd;
rom[120806] = 12'hddd;
rom[120807] = 12'hddd;
rom[120808] = 12'hddd;
rom[120809] = 12'hddd;
rom[120810] = 12'hddd;
rom[120811] = 12'hddd;
rom[120812] = 12'hddd;
rom[120813] = 12'hddd;
rom[120814] = 12'hddd;
rom[120815] = 12'hddd;
rom[120816] = 12'hddd;
rom[120817] = 12'hddd;
rom[120818] = 12'hddd;
rom[120819] = 12'hddd;
rom[120820] = 12'hddd;
rom[120821] = 12'hddd;
rom[120822] = 12'hddd;
rom[120823] = 12'hccc;
rom[120824] = 12'hccc;
rom[120825] = 12'hccc;
rom[120826] = 12'hccc;
rom[120827] = 12'hccc;
rom[120828] = 12'hccc;
rom[120829] = 12'hccc;
rom[120830] = 12'hccc;
rom[120831] = 12'hccc;
rom[120832] = 12'hccc;
rom[120833] = 12'hccc;
rom[120834] = 12'hccc;
rom[120835] = 12'hccc;
rom[120836] = 12'hccc;
rom[120837] = 12'hccc;
rom[120838] = 12'hccc;
rom[120839] = 12'hccc;
rom[120840] = 12'hbbb;
rom[120841] = 12'hbbb;
rom[120842] = 12'hbbb;
rom[120843] = 12'hbbb;
rom[120844] = 12'hbbb;
rom[120845] = 12'hbbb;
rom[120846] = 12'hbbb;
rom[120847] = 12'hbbb;
rom[120848] = 12'hbbb;
rom[120849] = 12'hbbb;
rom[120850] = 12'hbbb;
rom[120851] = 12'hbbb;
rom[120852] = 12'haaa;
rom[120853] = 12'haaa;
rom[120854] = 12'haaa;
rom[120855] = 12'haaa;
rom[120856] = 12'haaa;
rom[120857] = 12'haaa;
rom[120858] = 12'haaa;
rom[120859] = 12'haaa;
rom[120860] = 12'haaa;
rom[120861] = 12'haaa;
rom[120862] = 12'haaa;
rom[120863] = 12'haaa;
rom[120864] = 12'haaa;
rom[120865] = 12'haaa;
rom[120866] = 12'haaa;
rom[120867] = 12'haaa;
rom[120868] = 12'hccc;
rom[120869] = 12'heee;
rom[120870] = 12'hfff;
rom[120871] = 12'hfff;
rom[120872] = 12'heee;
rom[120873] = 12'hccc;
rom[120874] = 12'haaa;
rom[120875] = 12'h999;
rom[120876] = 12'h888;
rom[120877] = 12'h888;
rom[120878] = 12'h888;
rom[120879] = 12'h888;
rom[120880] = 12'h888;
rom[120881] = 12'h888;
rom[120882] = 12'h888;
rom[120883] = 12'h888;
rom[120884] = 12'h777;
rom[120885] = 12'h666;
rom[120886] = 12'h666;
rom[120887] = 12'h666;
rom[120888] = 12'h666;
rom[120889] = 12'h999;
rom[120890] = 12'hbbb;
rom[120891] = 12'haaa;
rom[120892] = 12'h888;
rom[120893] = 12'h777;
rom[120894] = 12'h666;
rom[120895] = 12'h666;
rom[120896] = 12'h666;
rom[120897] = 12'h555;
rom[120898] = 12'h666;
rom[120899] = 12'h666;
rom[120900] = 12'h666;
rom[120901] = 12'h777;
rom[120902] = 12'h777;
rom[120903] = 12'h777;
rom[120904] = 12'h777;
rom[120905] = 12'h666;
rom[120906] = 12'h666;
rom[120907] = 12'h666;
rom[120908] = 12'h666;
rom[120909] = 12'h666;
rom[120910] = 12'h666;
rom[120911] = 12'h555;
rom[120912] = 12'h444;
rom[120913] = 12'h444;
rom[120914] = 12'h444;
rom[120915] = 12'h444;
rom[120916] = 12'h444;
rom[120917] = 12'h444;
rom[120918] = 12'h555;
rom[120919] = 12'h555;
rom[120920] = 12'h666;
rom[120921] = 12'h555;
rom[120922] = 12'h555;
rom[120923] = 12'h555;
rom[120924] = 12'h555;
rom[120925] = 12'h555;
rom[120926] = 12'h555;
rom[120927] = 12'h555;
rom[120928] = 12'h555;
rom[120929] = 12'h555;
rom[120930] = 12'h444;
rom[120931] = 12'h444;
rom[120932] = 12'h444;
rom[120933] = 12'h444;
rom[120934] = 12'h444;
rom[120935] = 12'h333;
rom[120936] = 12'h333;
rom[120937] = 12'h333;
rom[120938] = 12'h333;
rom[120939] = 12'h333;
rom[120940] = 12'h333;
rom[120941] = 12'h333;
rom[120942] = 12'h333;
rom[120943] = 12'h333;
rom[120944] = 12'h333;
rom[120945] = 12'h333;
rom[120946] = 12'h333;
rom[120947] = 12'h333;
rom[120948] = 12'h333;
rom[120949] = 12'h333;
rom[120950] = 12'h333;
rom[120951] = 12'h333;
rom[120952] = 12'h333;
rom[120953] = 12'h333;
rom[120954] = 12'h333;
rom[120955] = 12'h333;
rom[120956] = 12'h333;
rom[120957] = 12'h333;
rom[120958] = 12'h333;
rom[120959] = 12'h222;
rom[120960] = 12'h333;
rom[120961] = 12'h333;
rom[120962] = 12'h333;
rom[120963] = 12'h333;
rom[120964] = 12'h333;
rom[120965] = 12'h333;
rom[120966] = 12'h333;
rom[120967] = 12'h333;
rom[120968] = 12'h333;
rom[120969] = 12'h222;
rom[120970] = 12'h222;
rom[120971] = 12'h222;
rom[120972] = 12'h222;
rom[120973] = 12'h222;
rom[120974] = 12'h111;
rom[120975] = 12'h111;
rom[120976] = 12'h111;
rom[120977] = 12'h111;
rom[120978] = 12'h111;
rom[120979] = 12'h111;
rom[120980] = 12'h222;
rom[120981] = 12'h222;
rom[120982] = 12'h222;
rom[120983] = 12'h222;
rom[120984] = 12'h111;
rom[120985] = 12'h111;
rom[120986] = 12'h111;
rom[120987] = 12'h111;
rom[120988] = 12'h111;
rom[120989] = 12'h111;
rom[120990] = 12'h222;
rom[120991] = 12'h222;
rom[120992] = 12'h222;
rom[120993] = 12'h333;
rom[120994] = 12'h333;
rom[120995] = 12'h333;
rom[120996] = 12'h222;
rom[120997] = 12'h111;
rom[120998] = 12'h111;
rom[120999] = 12'h  0;
rom[121000] = 12'h  0;
rom[121001] = 12'h  0;
rom[121002] = 12'h  0;
rom[121003] = 12'h111;
rom[121004] = 12'h111;
rom[121005] = 12'h  0;
rom[121006] = 12'h  0;
rom[121007] = 12'h  0;
rom[121008] = 12'h  0;
rom[121009] = 12'h  0;
rom[121010] = 12'h  0;
rom[121011] = 12'h  0;
rom[121012] = 12'h  0;
rom[121013] = 12'h  0;
rom[121014] = 12'h  0;
rom[121015] = 12'h111;
rom[121016] = 12'h111;
rom[121017] = 12'h111;
rom[121018] = 12'h111;
rom[121019] = 12'h  0;
rom[121020] = 12'h  0;
rom[121021] = 12'h  0;
rom[121022] = 12'h  0;
rom[121023] = 12'h  0;
rom[121024] = 12'h  0;
rom[121025] = 12'h  0;
rom[121026] = 12'h  0;
rom[121027] = 12'h  0;
rom[121028] = 12'h  0;
rom[121029] = 12'h  0;
rom[121030] = 12'h  0;
rom[121031] = 12'h  0;
rom[121032] = 12'h222;
rom[121033] = 12'h222;
rom[121034] = 12'h222;
rom[121035] = 12'h333;
rom[121036] = 12'h444;
rom[121037] = 12'h444;
rom[121038] = 12'h333;
rom[121039] = 12'h111;
rom[121040] = 12'h  0;
rom[121041] = 12'h  0;
rom[121042] = 12'h  0;
rom[121043] = 12'h  0;
rom[121044] = 12'h  0;
rom[121045] = 12'h  0;
rom[121046] = 12'h  0;
rom[121047] = 12'h  0;
rom[121048] = 12'h  0;
rom[121049] = 12'h  0;
rom[121050] = 12'h  0;
rom[121051] = 12'h  0;
rom[121052] = 12'h  0;
rom[121053] = 12'h  0;
rom[121054] = 12'h  0;
rom[121055] = 12'h  0;
rom[121056] = 12'h  0;
rom[121057] = 12'h  0;
rom[121058] = 12'h  0;
rom[121059] = 12'h  0;
rom[121060] = 12'h  0;
rom[121061] = 12'h  0;
rom[121062] = 12'h222;
rom[121063] = 12'h777;
rom[121064] = 12'heee;
rom[121065] = 12'hddd;
rom[121066] = 12'h888;
rom[121067] = 12'h222;
rom[121068] = 12'h111;
rom[121069] = 12'h111;
rom[121070] = 12'h  0;
rom[121071] = 12'h  0;
rom[121072] = 12'h  0;
rom[121073] = 12'h  0;
rom[121074] = 12'h  0;
rom[121075] = 12'h  0;
rom[121076] = 12'h  0;
rom[121077] = 12'h222;
rom[121078] = 12'h777;
rom[121079] = 12'hbbb;
rom[121080] = 12'h888;
rom[121081] = 12'h333;
rom[121082] = 12'h  0;
rom[121083] = 12'h  0;
rom[121084] = 12'h  0;
rom[121085] = 12'h  0;
rom[121086] = 12'h  0;
rom[121087] = 12'h  0;
rom[121088] = 12'h  0;
rom[121089] = 12'h  0;
rom[121090] = 12'h  0;
rom[121091] = 12'h111;
rom[121092] = 12'h222;
rom[121093] = 12'h333;
rom[121094] = 12'h222;
rom[121095] = 12'h111;
rom[121096] = 12'h  0;
rom[121097] = 12'h  0;
rom[121098] = 12'h  0;
rom[121099] = 12'h111;
rom[121100] = 12'h333;
rom[121101] = 12'h444;
rom[121102] = 12'h333;
rom[121103] = 12'h111;
rom[121104] = 12'h  0;
rom[121105] = 12'h  0;
rom[121106] = 12'h  0;
rom[121107] = 12'h  0;
rom[121108] = 12'h  0;
rom[121109] = 12'h  0;
rom[121110] = 12'h  0;
rom[121111] = 12'h  0;
rom[121112] = 12'h  0;
rom[121113] = 12'h  0;
rom[121114] = 12'h111;
rom[121115] = 12'h111;
rom[121116] = 12'h111;
rom[121117] = 12'h111;
rom[121118] = 12'h222;
rom[121119] = 12'h333;
rom[121120] = 12'h666;
rom[121121] = 12'h777;
rom[121122] = 12'h666;
rom[121123] = 12'h333;
rom[121124] = 12'h111;
rom[121125] = 12'h  0;
rom[121126] = 12'h  0;
rom[121127] = 12'h  0;
rom[121128] = 12'h  0;
rom[121129] = 12'h  0;
rom[121130] = 12'h  0;
rom[121131] = 12'h  0;
rom[121132] = 12'h  0;
rom[121133] = 12'h  0;
rom[121134] = 12'h  0;
rom[121135] = 12'h  0;
rom[121136] = 12'h  0;
rom[121137] = 12'h  0;
rom[121138] = 12'h  0;
rom[121139] = 12'h  0;
rom[121140] = 12'h  0;
rom[121141] = 12'h  0;
rom[121142] = 12'h  0;
rom[121143] = 12'h  0;
rom[121144] = 12'h  0;
rom[121145] = 12'h  0;
rom[121146] = 12'h  0;
rom[121147] = 12'h  0;
rom[121148] = 12'h  0;
rom[121149] = 12'h  0;
rom[121150] = 12'h  0;
rom[121151] = 12'h  0;
rom[121152] = 12'h  0;
rom[121153] = 12'h  0;
rom[121154] = 12'h  0;
rom[121155] = 12'h  0;
rom[121156] = 12'h  0;
rom[121157] = 12'h  0;
rom[121158] = 12'h  0;
rom[121159] = 12'h  0;
rom[121160] = 12'h  0;
rom[121161] = 12'h  0;
rom[121162] = 12'h  0;
rom[121163] = 12'h  0;
rom[121164] = 12'h  0;
rom[121165] = 12'h  0;
rom[121166] = 12'h  0;
rom[121167] = 12'h  0;
rom[121168] = 12'h  0;
rom[121169] = 12'h  0;
rom[121170] = 12'h  0;
rom[121171] = 12'h  0;
rom[121172] = 12'h  0;
rom[121173] = 12'h  0;
rom[121174] = 12'h111;
rom[121175] = 12'h222;
rom[121176] = 12'h555;
rom[121177] = 12'h666;
rom[121178] = 12'h777;
rom[121179] = 12'h555;
rom[121180] = 12'h222;
rom[121181] = 12'h111;
rom[121182] = 12'h  0;
rom[121183] = 12'h  0;
rom[121184] = 12'h  0;
rom[121185] = 12'h  0;
rom[121186] = 12'h  0;
rom[121187] = 12'h  0;
rom[121188] = 12'h  0;
rom[121189] = 12'h  0;
rom[121190] = 12'h  0;
rom[121191] = 12'h  0;
rom[121192] = 12'h  0;
rom[121193] = 12'h  0;
rom[121194] = 12'h  0;
rom[121195] = 12'h  0;
rom[121196] = 12'h  0;
rom[121197] = 12'h  0;
rom[121198] = 12'h  0;
rom[121199] = 12'h  0;
rom[121200] = 12'heee;
rom[121201] = 12'heee;
rom[121202] = 12'heee;
rom[121203] = 12'heee;
rom[121204] = 12'hddd;
rom[121205] = 12'hddd;
rom[121206] = 12'hddd;
rom[121207] = 12'hddd;
rom[121208] = 12'hddd;
rom[121209] = 12'hddd;
rom[121210] = 12'hddd;
rom[121211] = 12'hddd;
rom[121212] = 12'hddd;
rom[121213] = 12'hddd;
rom[121214] = 12'hddd;
rom[121215] = 12'hddd;
rom[121216] = 12'hddd;
rom[121217] = 12'hddd;
rom[121218] = 12'hddd;
rom[121219] = 12'hddd;
rom[121220] = 12'hddd;
rom[121221] = 12'hddd;
rom[121222] = 12'hccc;
rom[121223] = 12'hccc;
rom[121224] = 12'hccc;
rom[121225] = 12'hccc;
rom[121226] = 12'hccc;
rom[121227] = 12'hccc;
rom[121228] = 12'hccc;
rom[121229] = 12'hccc;
rom[121230] = 12'hccc;
rom[121231] = 12'hccc;
rom[121232] = 12'hccc;
rom[121233] = 12'hccc;
rom[121234] = 12'hccc;
rom[121235] = 12'hccc;
rom[121236] = 12'hccc;
rom[121237] = 12'hccc;
rom[121238] = 12'hccc;
rom[121239] = 12'hccc;
rom[121240] = 12'hbbb;
rom[121241] = 12'hbbb;
rom[121242] = 12'hbbb;
rom[121243] = 12'hbbb;
rom[121244] = 12'hbbb;
rom[121245] = 12'hbbb;
rom[121246] = 12'hbbb;
rom[121247] = 12'hbbb;
rom[121248] = 12'hbbb;
rom[121249] = 12'hbbb;
rom[121250] = 12'haaa;
rom[121251] = 12'haaa;
rom[121252] = 12'haaa;
rom[121253] = 12'haaa;
rom[121254] = 12'haaa;
rom[121255] = 12'haaa;
rom[121256] = 12'haaa;
rom[121257] = 12'haaa;
rom[121258] = 12'haaa;
rom[121259] = 12'haaa;
rom[121260] = 12'haaa;
rom[121261] = 12'haaa;
rom[121262] = 12'h999;
rom[121263] = 12'h999;
rom[121264] = 12'haaa;
rom[121265] = 12'haaa;
rom[121266] = 12'haaa;
rom[121267] = 12'hbbb;
rom[121268] = 12'hddd;
rom[121269] = 12'hfff;
rom[121270] = 12'hfff;
rom[121271] = 12'hfff;
rom[121272] = 12'hddd;
rom[121273] = 12'hbbb;
rom[121274] = 12'h888;
rom[121275] = 12'h888;
rom[121276] = 12'h888;
rom[121277] = 12'h888;
rom[121278] = 12'h888;
rom[121279] = 12'h888;
rom[121280] = 12'h888;
rom[121281] = 12'h888;
rom[121282] = 12'h888;
rom[121283] = 12'h888;
rom[121284] = 12'h777;
rom[121285] = 12'h666;
rom[121286] = 12'h666;
rom[121287] = 12'h666;
rom[121288] = 12'h888;
rom[121289] = 12'haaa;
rom[121290] = 12'hbbb;
rom[121291] = 12'haaa;
rom[121292] = 12'h777;
rom[121293] = 12'h666;
rom[121294] = 12'h555;
rom[121295] = 12'h555;
rom[121296] = 12'h555;
rom[121297] = 12'h555;
rom[121298] = 12'h666;
rom[121299] = 12'h666;
rom[121300] = 12'h666;
rom[121301] = 12'h666;
rom[121302] = 12'h777;
rom[121303] = 12'h777;
rom[121304] = 12'h777;
rom[121305] = 12'h666;
rom[121306] = 12'h666;
rom[121307] = 12'h666;
rom[121308] = 12'h666;
rom[121309] = 12'h666;
rom[121310] = 12'h666;
rom[121311] = 12'h555;
rom[121312] = 12'h444;
rom[121313] = 12'h444;
rom[121314] = 12'h444;
rom[121315] = 12'h444;
rom[121316] = 12'h444;
rom[121317] = 12'h444;
rom[121318] = 12'h555;
rom[121319] = 12'h555;
rom[121320] = 12'h555;
rom[121321] = 12'h555;
rom[121322] = 12'h555;
rom[121323] = 12'h555;
rom[121324] = 12'h555;
rom[121325] = 12'h555;
rom[121326] = 12'h555;
rom[121327] = 12'h555;
rom[121328] = 12'h555;
rom[121329] = 12'h555;
rom[121330] = 12'h444;
rom[121331] = 12'h444;
rom[121332] = 12'h444;
rom[121333] = 12'h444;
rom[121334] = 12'h444;
rom[121335] = 12'h333;
rom[121336] = 12'h333;
rom[121337] = 12'h333;
rom[121338] = 12'h333;
rom[121339] = 12'h333;
rom[121340] = 12'h333;
rom[121341] = 12'h333;
rom[121342] = 12'h333;
rom[121343] = 12'h333;
rom[121344] = 12'h333;
rom[121345] = 12'h333;
rom[121346] = 12'h333;
rom[121347] = 12'h333;
rom[121348] = 12'h333;
rom[121349] = 12'h333;
rom[121350] = 12'h333;
rom[121351] = 12'h333;
rom[121352] = 12'h333;
rom[121353] = 12'h333;
rom[121354] = 12'h333;
rom[121355] = 12'h333;
rom[121356] = 12'h333;
rom[121357] = 12'h333;
rom[121358] = 12'h222;
rom[121359] = 12'h222;
rom[121360] = 12'h222;
rom[121361] = 12'h333;
rom[121362] = 12'h333;
rom[121363] = 12'h333;
rom[121364] = 12'h333;
rom[121365] = 12'h333;
rom[121366] = 12'h333;
rom[121367] = 12'h222;
rom[121368] = 12'h222;
rom[121369] = 12'h222;
rom[121370] = 12'h222;
rom[121371] = 12'h222;
rom[121372] = 12'h222;
rom[121373] = 12'h222;
rom[121374] = 12'h111;
rom[121375] = 12'h111;
rom[121376] = 12'h111;
rom[121377] = 12'h111;
rom[121378] = 12'h111;
rom[121379] = 12'h111;
rom[121380] = 12'h222;
rom[121381] = 12'h222;
rom[121382] = 12'h222;
rom[121383] = 12'h222;
rom[121384] = 12'h111;
rom[121385] = 12'h111;
rom[121386] = 12'h111;
rom[121387] = 12'h111;
rom[121388] = 12'h111;
rom[121389] = 12'h111;
rom[121390] = 12'h111;
rom[121391] = 12'h222;
rom[121392] = 12'h222;
rom[121393] = 12'h222;
rom[121394] = 12'h222;
rom[121395] = 12'h222;
rom[121396] = 12'h222;
rom[121397] = 12'h111;
rom[121398] = 12'h  0;
rom[121399] = 12'h  0;
rom[121400] = 12'h  0;
rom[121401] = 12'h  0;
rom[121402] = 12'h  0;
rom[121403] = 12'h  0;
rom[121404] = 12'h  0;
rom[121405] = 12'h  0;
rom[121406] = 12'h  0;
rom[121407] = 12'h  0;
rom[121408] = 12'h  0;
rom[121409] = 12'h  0;
rom[121410] = 12'h  0;
rom[121411] = 12'h  0;
rom[121412] = 12'h  0;
rom[121413] = 12'h  0;
rom[121414] = 12'h  0;
rom[121415] = 12'h  0;
rom[121416] = 12'h  0;
rom[121417] = 12'h  0;
rom[121418] = 12'h111;
rom[121419] = 12'h  0;
rom[121420] = 12'h  0;
rom[121421] = 12'h  0;
rom[121422] = 12'h  0;
rom[121423] = 12'h111;
rom[121424] = 12'h  0;
rom[121425] = 12'h  0;
rom[121426] = 12'h  0;
rom[121427] = 12'h  0;
rom[121428] = 12'h  0;
rom[121429] = 12'h  0;
rom[121430] = 12'h  0;
rom[121431] = 12'h  0;
rom[121432] = 12'h111;
rom[121433] = 12'h111;
rom[121434] = 12'h222;
rom[121435] = 12'h333;
rom[121436] = 12'h444;
rom[121437] = 12'h333;
rom[121438] = 12'h222;
rom[121439] = 12'h  0;
rom[121440] = 12'h  0;
rom[121441] = 12'h  0;
rom[121442] = 12'h  0;
rom[121443] = 12'h  0;
rom[121444] = 12'h  0;
rom[121445] = 12'h  0;
rom[121446] = 12'h  0;
rom[121447] = 12'h  0;
rom[121448] = 12'h  0;
rom[121449] = 12'h  0;
rom[121450] = 12'h  0;
rom[121451] = 12'h  0;
rom[121452] = 12'h  0;
rom[121453] = 12'h  0;
rom[121454] = 12'h  0;
rom[121455] = 12'h  0;
rom[121456] = 12'h  0;
rom[121457] = 12'h  0;
rom[121458] = 12'h  0;
rom[121459] = 12'h  0;
rom[121460] = 12'h  0;
rom[121461] = 12'h  0;
rom[121462] = 12'h222;
rom[121463] = 12'h777;
rom[121464] = 12'heee;
rom[121465] = 12'hddd;
rom[121466] = 12'h777;
rom[121467] = 12'h222;
rom[121468] = 12'h111;
rom[121469] = 12'h111;
rom[121470] = 12'h  0;
rom[121471] = 12'h  0;
rom[121472] = 12'h  0;
rom[121473] = 12'h  0;
rom[121474] = 12'h  0;
rom[121475] = 12'h  0;
rom[121476] = 12'h  0;
rom[121477] = 12'h222;
rom[121478] = 12'h777;
rom[121479] = 12'haaa;
rom[121480] = 12'h999;
rom[121481] = 12'h444;
rom[121482] = 12'h111;
rom[121483] = 12'h  0;
rom[121484] = 12'h111;
rom[121485] = 12'h111;
rom[121486] = 12'h111;
rom[121487] = 12'h  0;
rom[121488] = 12'h  0;
rom[121489] = 12'h  0;
rom[121490] = 12'h  0;
rom[121491] = 12'h  0;
rom[121492] = 12'h222;
rom[121493] = 12'h333;
rom[121494] = 12'h222;
rom[121495] = 12'h111;
rom[121496] = 12'h  0;
rom[121497] = 12'h  0;
rom[121498] = 12'h  0;
rom[121499] = 12'h  0;
rom[121500] = 12'h222;
rom[121501] = 12'h444;
rom[121502] = 12'h333;
rom[121503] = 12'h222;
rom[121504] = 12'h  0;
rom[121505] = 12'h  0;
rom[121506] = 12'h  0;
rom[121507] = 12'h  0;
rom[121508] = 12'h  0;
rom[121509] = 12'h  0;
rom[121510] = 12'h  0;
rom[121511] = 12'h  0;
rom[121512] = 12'h  0;
rom[121513] = 12'h  0;
rom[121514] = 12'h  0;
rom[121515] = 12'h  0;
rom[121516] = 12'h  0;
rom[121517] = 12'h  0;
rom[121518] = 12'h111;
rom[121519] = 12'h333;
rom[121520] = 12'h666;
rom[121521] = 12'h777;
rom[121522] = 12'h666;
rom[121523] = 12'h333;
rom[121524] = 12'h111;
rom[121525] = 12'h111;
rom[121526] = 12'h111;
rom[121527] = 12'h  0;
rom[121528] = 12'h  0;
rom[121529] = 12'h  0;
rom[121530] = 12'h  0;
rom[121531] = 12'h  0;
rom[121532] = 12'h  0;
rom[121533] = 12'h  0;
rom[121534] = 12'h  0;
rom[121535] = 12'h  0;
rom[121536] = 12'h  0;
rom[121537] = 12'h  0;
rom[121538] = 12'h  0;
rom[121539] = 12'h  0;
rom[121540] = 12'h  0;
rom[121541] = 12'h  0;
rom[121542] = 12'h  0;
rom[121543] = 12'h  0;
rom[121544] = 12'h  0;
rom[121545] = 12'h  0;
rom[121546] = 12'h  0;
rom[121547] = 12'h  0;
rom[121548] = 12'h  0;
rom[121549] = 12'h  0;
rom[121550] = 12'h  0;
rom[121551] = 12'h  0;
rom[121552] = 12'h  0;
rom[121553] = 12'h  0;
rom[121554] = 12'h  0;
rom[121555] = 12'h  0;
rom[121556] = 12'h  0;
rom[121557] = 12'h  0;
rom[121558] = 12'h  0;
rom[121559] = 12'h  0;
rom[121560] = 12'h  0;
rom[121561] = 12'h  0;
rom[121562] = 12'h  0;
rom[121563] = 12'h  0;
rom[121564] = 12'h  0;
rom[121565] = 12'h  0;
rom[121566] = 12'h  0;
rom[121567] = 12'h  0;
rom[121568] = 12'h  0;
rom[121569] = 12'h  0;
rom[121570] = 12'h  0;
rom[121571] = 12'h  0;
rom[121572] = 12'h  0;
rom[121573] = 12'h  0;
rom[121574] = 12'h111;
rom[121575] = 12'h111;
rom[121576] = 12'h444;
rom[121577] = 12'h555;
rom[121578] = 12'h666;
rom[121579] = 12'h555;
rom[121580] = 12'h333;
rom[121581] = 12'h111;
rom[121582] = 12'h  0;
rom[121583] = 12'h111;
rom[121584] = 12'h  0;
rom[121585] = 12'h  0;
rom[121586] = 12'h  0;
rom[121587] = 12'h  0;
rom[121588] = 12'h  0;
rom[121589] = 12'h  0;
rom[121590] = 12'h  0;
rom[121591] = 12'h  0;
rom[121592] = 12'h  0;
rom[121593] = 12'h  0;
rom[121594] = 12'h  0;
rom[121595] = 12'h  0;
rom[121596] = 12'h  0;
rom[121597] = 12'h  0;
rom[121598] = 12'h  0;
rom[121599] = 12'h  0;
rom[121600] = 12'heee;
rom[121601] = 12'heee;
rom[121602] = 12'heee;
rom[121603] = 12'heee;
rom[121604] = 12'hddd;
rom[121605] = 12'hddd;
rom[121606] = 12'hddd;
rom[121607] = 12'hddd;
rom[121608] = 12'hddd;
rom[121609] = 12'hddd;
rom[121610] = 12'hddd;
rom[121611] = 12'hddd;
rom[121612] = 12'hddd;
rom[121613] = 12'hddd;
rom[121614] = 12'hddd;
rom[121615] = 12'hddd;
rom[121616] = 12'hddd;
rom[121617] = 12'hddd;
rom[121618] = 12'hddd;
rom[121619] = 12'hddd;
rom[121620] = 12'hddd;
rom[121621] = 12'hddd;
rom[121622] = 12'hccc;
rom[121623] = 12'hccc;
rom[121624] = 12'hccc;
rom[121625] = 12'hccc;
rom[121626] = 12'hccc;
rom[121627] = 12'hccc;
rom[121628] = 12'hccc;
rom[121629] = 12'hccc;
rom[121630] = 12'hccc;
rom[121631] = 12'hccc;
rom[121632] = 12'hccc;
rom[121633] = 12'hccc;
rom[121634] = 12'hccc;
rom[121635] = 12'hccc;
rom[121636] = 12'hbbb;
rom[121637] = 12'hbbb;
rom[121638] = 12'hbbb;
rom[121639] = 12'hbbb;
rom[121640] = 12'hbbb;
rom[121641] = 12'hbbb;
rom[121642] = 12'hbbb;
rom[121643] = 12'hbbb;
rom[121644] = 12'hbbb;
rom[121645] = 12'hbbb;
rom[121646] = 12'haaa;
rom[121647] = 12'haaa;
rom[121648] = 12'haaa;
rom[121649] = 12'haaa;
rom[121650] = 12'haaa;
rom[121651] = 12'haaa;
rom[121652] = 12'haaa;
rom[121653] = 12'haaa;
rom[121654] = 12'haaa;
rom[121655] = 12'h999;
rom[121656] = 12'h999;
rom[121657] = 12'haaa;
rom[121658] = 12'haaa;
rom[121659] = 12'haaa;
rom[121660] = 12'h999;
rom[121661] = 12'h999;
rom[121662] = 12'h999;
rom[121663] = 12'h999;
rom[121664] = 12'haaa;
rom[121665] = 12'haaa;
rom[121666] = 12'haaa;
rom[121667] = 12'hccc;
rom[121668] = 12'hfff;
rom[121669] = 12'hfff;
rom[121670] = 12'hfff;
rom[121671] = 12'hddd;
rom[121672] = 12'hbbb;
rom[121673] = 12'h999;
rom[121674] = 12'h888;
rom[121675] = 12'h777;
rom[121676] = 12'h777;
rom[121677] = 12'h777;
rom[121678] = 12'h777;
rom[121679] = 12'h777;
rom[121680] = 12'h888;
rom[121681] = 12'h777;
rom[121682] = 12'h777;
rom[121683] = 12'h888;
rom[121684] = 12'h777;
rom[121685] = 12'h666;
rom[121686] = 12'h666;
rom[121687] = 12'h666;
rom[121688] = 12'haaa;
rom[121689] = 12'hbbb;
rom[121690] = 12'haaa;
rom[121691] = 12'h888;
rom[121692] = 12'h666;
rom[121693] = 12'h666;
rom[121694] = 12'h555;
rom[121695] = 12'h444;
rom[121696] = 12'h555;
rom[121697] = 12'h555;
rom[121698] = 12'h666;
rom[121699] = 12'h666;
rom[121700] = 12'h666;
rom[121701] = 12'h666;
rom[121702] = 12'h666;
rom[121703] = 12'h666;
rom[121704] = 12'h666;
rom[121705] = 12'h777;
rom[121706] = 12'h666;
rom[121707] = 12'h666;
rom[121708] = 12'h555;
rom[121709] = 12'h666;
rom[121710] = 12'h666;
rom[121711] = 12'h555;
rom[121712] = 12'h555;
rom[121713] = 12'h444;
rom[121714] = 12'h444;
rom[121715] = 12'h444;
rom[121716] = 12'h444;
rom[121717] = 12'h444;
rom[121718] = 12'h555;
rom[121719] = 12'h555;
rom[121720] = 12'h555;
rom[121721] = 12'h555;
rom[121722] = 12'h555;
rom[121723] = 12'h555;
rom[121724] = 12'h555;
rom[121725] = 12'h555;
rom[121726] = 12'h555;
rom[121727] = 12'h555;
rom[121728] = 12'h666;
rom[121729] = 12'h555;
rom[121730] = 12'h444;
rom[121731] = 12'h444;
rom[121732] = 12'h444;
rom[121733] = 12'h444;
rom[121734] = 12'h333;
rom[121735] = 12'h333;
rom[121736] = 12'h333;
rom[121737] = 12'h333;
rom[121738] = 12'h333;
rom[121739] = 12'h333;
rom[121740] = 12'h333;
rom[121741] = 12'h333;
rom[121742] = 12'h222;
rom[121743] = 12'h222;
rom[121744] = 12'h333;
rom[121745] = 12'h333;
rom[121746] = 12'h333;
rom[121747] = 12'h333;
rom[121748] = 12'h333;
rom[121749] = 12'h333;
rom[121750] = 12'h333;
rom[121751] = 12'h333;
rom[121752] = 12'h333;
rom[121753] = 12'h333;
rom[121754] = 12'h333;
rom[121755] = 12'h222;
rom[121756] = 12'h222;
rom[121757] = 12'h222;
rom[121758] = 12'h222;
rom[121759] = 12'h222;
rom[121760] = 12'h333;
rom[121761] = 12'h333;
rom[121762] = 12'h333;
rom[121763] = 12'h333;
rom[121764] = 12'h333;
rom[121765] = 12'h333;
rom[121766] = 12'h222;
rom[121767] = 12'h222;
rom[121768] = 12'h222;
rom[121769] = 12'h222;
rom[121770] = 12'h111;
rom[121771] = 12'h111;
rom[121772] = 12'h111;
rom[121773] = 12'h111;
rom[121774] = 12'h111;
rom[121775] = 12'h111;
rom[121776] = 12'h111;
rom[121777] = 12'h111;
rom[121778] = 12'h111;
rom[121779] = 12'h111;
rom[121780] = 12'h111;
rom[121781] = 12'h222;
rom[121782] = 12'h222;
rom[121783] = 12'h222;
rom[121784] = 12'h111;
rom[121785] = 12'h111;
rom[121786] = 12'h  0;
rom[121787] = 12'h  0;
rom[121788] = 12'h111;
rom[121789] = 12'h111;
rom[121790] = 12'h111;
rom[121791] = 12'h111;
rom[121792] = 12'h222;
rom[121793] = 12'h222;
rom[121794] = 12'h333;
rom[121795] = 12'h222;
rom[121796] = 12'h222;
rom[121797] = 12'h111;
rom[121798] = 12'h  0;
rom[121799] = 12'h  0;
rom[121800] = 12'h  0;
rom[121801] = 12'h  0;
rom[121802] = 12'h  0;
rom[121803] = 12'h  0;
rom[121804] = 12'h  0;
rom[121805] = 12'h  0;
rom[121806] = 12'h  0;
rom[121807] = 12'h  0;
rom[121808] = 12'h  0;
rom[121809] = 12'h  0;
rom[121810] = 12'h  0;
rom[121811] = 12'h  0;
rom[121812] = 12'h  0;
rom[121813] = 12'h  0;
rom[121814] = 12'h  0;
rom[121815] = 12'h  0;
rom[121816] = 12'h  0;
rom[121817] = 12'h  0;
rom[121818] = 12'h  0;
rom[121819] = 12'h  0;
rom[121820] = 12'h  0;
rom[121821] = 12'h  0;
rom[121822] = 12'h  0;
rom[121823] = 12'h111;
rom[121824] = 12'h  0;
rom[121825] = 12'h  0;
rom[121826] = 12'h  0;
rom[121827] = 12'h  0;
rom[121828] = 12'h  0;
rom[121829] = 12'h  0;
rom[121830] = 12'h  0;
rom[121831] = 12'h  0;
rom[121832] = 12'h111;
rom[121833] = 12'h111;
rom[121834] = 12'h222;
rom[121835] = 12'h333;
rom[121836] = 12'h444;
rom[121837] = 12'h222;
rom[121838] = 12'h111;
rom[121839] = 12'h  0;
rom[121840] = 12'h  0;
rom[121841] = 12'h  0;
rom[121842] = 12'h  0;
rom[121843] = 12'h  0;
rom[121844] = 12'h  0;
rom[121845] = 12'h  0;
rom[121846] = 12'h  0;
rom[121847] = 12'h  0;
rom[121848] = 12'h  0;
rom[121849] = 12'h  0;
rom[121850] = 12'h  0;
rom[121851] = 12'h  0;
rom[121852] = 12'h  0;
rom[121853] = 12'h  0;
rom[121854] = 12'h  0;
rom[121855] = 12'h  0;
rom[121856] = 12'h  0;
rom[121857] = 12'h  0;
rom[121858] = 12'h  0;
rom[121859] = 12'h  0;
rom[121860] = 12'h  0;
rom[121861] = 12'h  0;
rom[121862] = 12'h333;
rom[121863] = 12'h888;
rom[121864] = 12'heee;
rom[121865] = 12'hccc;
rom[121866] = 12'h666;
rom[121867] = 12'h111;
rom[121868] = 12'h111;
rom[121869] = 12'h  0;
rom[121870] = 12'h  0;
rom[121871] = 12'h  0;
rom[121872] = 12'h  0;
rom[121873] = 12'h  0;
rom[121874] = 12'h  0;
rom[121875] = 12'h  0;
rom[121876] = 12'h  0;
rom[121877] = 12'h111;
rom[121878] = 12'h555;
rom[121879] = 12'haaa;
rom[121880] = 12'h999;
rom[121881] = 12'h444;
rom[121882] = 12'h111;
rom[121883] = 12'h111;
rom[121884] = 12'h  0;
rom[121885] = 12'h  0;
rom[121886] = 12'h111;
rom[121887] = 12'h  0;
rom[121888] = 12'h  0;
rom[121889] = 12'h  0;
rom[121890] = 12'h  0;
rom[121891] = 12'h  0;
rom[121892] = 12'h111;
rom[121893] = 12'h333;
rom[121894] = 12'h333;
rom[121895] = 12'h111;
rom[121896] = 12'h  0;
rom[121897] = 12'h  0;
rom[121898] = 12'h  0;
rom[121899] = 12'h  0;
rom[121900] = 12'h111;
rom[121901] = 12'h222;
rom[121902] = 12'h333;
rom[121903] = 12'h222;
rom[121904] = 12'h  0;
rom[121905] = 12'h  0;
rom[121906] = 12'h  0;
rom[121907] = 12'h  0;
rom[121908] = 12'h  0;
rom[121909] = 12'h  0;
rom[121910] = 12'h  0;
rom[121911] = 12'h  0;
rom[121912] = 12'h  0;
rom[121913] = 12'h  0;
rom[121914] = 12'h  0;
rom[121915] = 12'h  0;
rom[121916] = 12'h  0;
rom[121917] = 12'h  0;
rom[121918] = 12'h111;
rom[121919] = 12'h222;
rom[121920] = 12'h444;
rom[121921] = 12'h666;
rom[121922] = 12'h666;
rom[121923] = 12'h333;
rom[121924] = 12'h111;
rom[121925] = 12'h  0;
rom[121926] = 12'h  0;
rom[121927] = 12'h  0;
rom[121928] = 12'h  0;
rom[121929] = 12'h  0;
rom[121930] = 12'h  0;
rom[121931] = 12'h  0;
rom[121932] = 12'h  0;
rom[121933] = 12'h  0;
rom[121934] = 12'h  0;
rom[121935] = 12'h  0;
rom[121936] = 12'h  0;
rom[121937] = 12'h  0;
rom[121938] = 12'h  0;
rom[121939] = 12'h  0;
rom[121940] = 12'h  0;
rom[121941] = 12'h  0;
rom[121942] = 12'h  0;
rom[121943] = 12'h  0;
rom[121944] = 12'h  0;
rom[121945] = 12'h  0;
rom[121946] = 12'h  0;
rom[121947] = 12'h  0;
rom[121948] = 12'h  0;
rom[121949] = 12'h  0;
rom[121950] = 12'h  0;
rom[121951] = 12'h  0;
rom[121952] = 12'h  0;
rom[121953] = 12'h  0;
rom[121954] = 12'h  0;
rom[121955] = 12'h  0;
rom[121956] = 12'h  0;
rom[121957] = 12'h  0;
rom[121958] = 12'h  0;
rom[121959] = 12'h  0;
rom[121960] = 12'h  0;
rom[121961] = 12'h  0;
rom[121962] = 12'h  0;
rom[121963] = 12'h  0;
rom[121964] = 12'h  0;
rom[121965] = 12'h  0;
rom[121966] = 12'h  0;
rom[121967] = 12'h  0;
rom[121968] = 12'h  0;
rom[121969] = 12'h  0;
rom[121970] = 12'h  0;
rom[121971] = 12'h  0;
rom[121972] = 12'h  0;
rom[121973] = 12'h  0;
rom[121974] = 12'h111;
rom[121975] = 12'h111;
rom[121976] = 12'h333;
rom[121977] = 12'h555;
rom[121978] = 12'h666;
rom[121979] = 12'h666;
rom[121980] = 12'h444;
rom[121981] = 12'h111;
rom[121982] = 12'h  0;
rom[121983] = 12'h  0;
rom[121984] = 12'h  0;
rom[121985] = 12'h  0;
rom[121986] = 12'h  0;
rom[121987] = 12'h  0;
rom[121988] = 12'h  0;
rom[121989] = 12'h  0;
rom[121990] = 12'h  0;
rom[121991] = 12'h  0;
rom[121992] = 12'h  0;
rom[121993] = 12'h  0;
rom[121994] = 12'h  0;
rom[121995] = 12'h  0;
rom[121996] = 12'h  0;
rom[121997] = 12'h  0;
rom[121998] = 12'h  0;
rom[121999] = 12'h  0;
rom[122000] = 12'heee;
rom[122001] = 12'heee;
rom[122002] = 12'heee;
rom[122003] = 12'heee;
rom[122004] = 12'hddd;
rom[122005] = 12'hddd;
rom[122006] = 12'hddd;
rom[122007] = 12'hddd;
rom[122008] = 12'hddd;
rom[122009] = 12'hddd;
rom[122010] = 12'hddd;
rom[122011] = 12'hddd;
rom[122012] = 12'hddd;
rom[122013] = 12'hddd;
rom[122014] = 12'hddd;
rom[122015] = 12'hddd;
rom[122016] = 12'hddd;
rom[122017] = 12'hddd;
rom[122018] = 12'hddd;
rom[122019] = 12'hddd;
rom[122020] = 12'hccc;
rom[122021] = 12'hccc;
rom[122022] = 12'hccc;
rom[122023] = 12'hccc;
rom[122024] = 12'hccc;
rom[122025] = 12'hccc;
rom[122026] = 12'hccc;
rom[122027] = 12'hccc;
rom[122028] = 12'hccc;
rom[122029] = 12'hccc;
rom[122030] = 12'hccc;
rom[122031] = 12'hccc;
rom[122032] = 12'hccc;
rom[122033] = 12'hbbb;
rom[122034] = 12'hbbb;
rom[122035] = 12'hbbb;
rom[122036] = 12'hbbb;
rom[122037] = 12'hbbb;
rom[122038] = 12'hbbb;
rom[122039] = 12'hbbb;
rom[122040] = 12'hbbb;
rom[122041] = 12'hbbb;
rom[122042] = 12'haaa;
rom[122043] = 12'haaa;
rom[122044] = 12'haaa;
rom[122045] = 12'haaa;
rom[122046] = 12'haaa;
rom[122047] = 12'haaa;
rom[122048] = 12'haaa;
rom[122049] = 12'haaa;
rom[122050] = 12'h999;
rom[122051] = 12'h999;
rom[122052] = 12'h999;
rom[122053] = 12'h999;
rom[122054] = 12'h999;
rom[122055] = 12'h999;
rom[122056] = 12'h999;
rom[122057] = 12'h999;
rom[122058] = 12'h999;
rom[122059] = 12'h999;
rom[122060] = 12'h999;
rom[122061] = 12'h999;
rom[122062] = 12'h999;
rom[122063] = 12'h999;
rom[122064] = 12'h999;
rom[122065] = 12'haaa;
rom[122066] = 12'hbbb;
rom[122067] = 12'hddd;
rom[122068] = 12'hfff;
rom[122069] = 12'hfff;
rom[122070] = 12'heee;
rom[122071] = 12'hccc;
rom[122072] = 12'h999;
rom[122073] = 12'h888;
rom[122074] = 12'h777;
rom[122075] = 12'h777;
rom[122076] = 12'h777;
rom[122077] = 12'h777;
rom[122078] = 12'h666;
rom[122079] = 12'h777;
rom[122080] = 12'h777;
rom[122081] = 12'h777;
rom[122082] = 12'h777;
rom[122083] = 12'h888;
rom[122084] = 12'h777;
rom[122085] = 12'h777;
rom[122086] = 12'h777;
rom[122087] = 12'h777;
rom[122088] = 12'hbbb;
rom[122089] = 12'haaa;
rom[122090] = 12'h999;
rom[122091] = 12'h666;
rom[122092] = 12'h555;
rom[122093] = 12'h555;
rom[122094] = 12'h555;
rom[122095] = 12'h555;
rom[122096] = 12'h444;
rom[122097] = 12'h555;
rom[122098] = 12'h666;
rom[122099] = 12'h666;
rom[122100] = 12'h666;
rom[122101] = 12'h666;
rom[122102] = 12'h666;
rom[122103] = 12'h666;
rom[122104] = 12'h666;
rom[122105] = 12'h666;
rom[122106] = 12'h666;
rom[122107] = 12'h666;
rom[122108] = 12'h666;
rom[122109] = 12'h666;
rom[122110] = 12'h666;
rom[122111] = 12'h555;
rom[122112] = 12'h555;
rom[122113] = 12'h444;
rom[122114] = 12'h444;
rom[122115] = 12'h444;
rom[122116] = 12'h444;
rom[122117] = 12'h444;
rom[122118] = 12'h555;
rom[122119] = 12'h555;
rom[122120] = 12'h555;
rom[122121] = 12'h555;
rom[122122] = 12'h555;
rom[122123] = 12'h555;
rom[122124] = 12'h555;
rom[122125] = 12'h444;
rom[122126] = 12'h444;
rom[122127] = 12'h555;
rom[122128] = 12'h555;
rom[122129] = 12'h555;
rom[122130] = 12'h444;
rom[122131] = 12'h444;
rom[122132] = 12'h444;
rom[122133] = 12'h444;
rom[122134] = 12'h333;
rom[122135] = 12'h333;
rom[122136] = 12'h333;
rom[122137] = 12'h333;
rom[122138] = 12'h333;
rom[122139] = 12'h333;
rom[122140] = 12'h333;
rom[122141] = 12'h333;
rom[122142] = 12'h222;
rom[122143] = 12'h222;
rom[122144] = 12'h333;
rom[122145] = 12'h333;
rom[122146] = 12'h333;
rom[122147] = 12'h333;
rom[122148] = 12'h333;
rom[122149] = 12'h333;
rom[122150] = 12'h333;
rom[122151] = 12'h333;
rom[122152] = 12'h333;
rom[122153] = 12'h333;
rom[122154] = 12'h222;
rom[122155] = 12'h222;
rom[122156] = 12'h222;
rom[122157] = 12'h222;
rom[122158] = 12'h222;
rom[122159] = 12'h222;
rom[122160] = 12'h333;
rom[122161] = 12'h333;
rom[122162] = 12'h333;
rom[122163] = 12'h333;
rom[122164] = 12'h333;
rom[122165] = 12'h222;
rom[122166] = 12'h222;
rom[122167] = 12'h222;
rom[122168] = 12'h222;
rom[122169] = 12'h111;
rom[122170] = 12'h111;
rom[122171] = 12'h111;
rom[122172] = 12'h111;
rom[122173] = 12'h111;
rom[122174] = 12'h111;
rom[122175] = 12'h111;
rom[122176] = 12'h111;
rom[122177] = 12'h111;
rom[122178] = 12'h111;
rom[122179] = 12'h111;
rom[122180] = 12'h111;
rom[122181] = 12'h222;
rom[122182] = 12'h222;
rom[122183] = 12'h222;
rom[122184] = 12'h111;
rom[122185] = 12'h111;
rom[122186] = 12'h  0;
rom[122187] = 12'h  0;
rom[122188] = 12'h111;
rom[122189] = 12'h111;
rom[122190] = 12'h111;
rom[122191] = 12'h111;
rom[122192] = 12'h222;
rom[122193] = 12'h222;
rom[122194] = 12'h222;
rom[122195] = 12'h222;
rom[122196] = 12'h222;
rom[122197] = 12'h111;
rom[122198] = 12'h  0;
rom[122199] = 12'h  0;
rom[122200] = 12'h  0;
rom[122201] = 12'h  0;
rom[122202] = 12'h  0;
rom[122203] = 12'h  0;
rom[122204] = 12'h  0;
rom[122205] = 12'h  0;
rom[122206] = 12'h  0;
rom[122207] = 12'h  0;
rom[122208] = 12'h  0;
rom[122209] = 12'h  0;
rom[122210] = 12'h  0;
rom[122211] = 12'h  0;
rom[122212] = 12'h  0;
rom[122213] = 12'h  0;
rom[122214] = 12'h  0;
rom[122215] = 12'h  0;
rom[122216] = 12'h  0;
rom[122217] = 12'h  0;
rom[122218] = 12'h  0;
rom[122219] = 12'h  0;
rom[122220] = 12'h  0;
rom[122221] = 12'h  0;
rom[122222] = 12'h  0;
rom[122223] = 12'h  0;
rom[122224] = 12'h  0;
rom[122225] = 12'h  0;
rom[122226] = 12'h  0;
rom[122227] = 12'h  0;
rom[122228] = 12'h  0;
rom[122229] = 12'h  0;
rom[122230] = 12'h  0;
rom[122231] = 12'h  0;
rom[122232] = 12'h  0;
rom[122233] = 12'h111;
rom[122234] = 12'h222;
rom[122235] = 12'h333;
rom[122236] = 12'h333;
rom[122237] = 12'h222;
rom[122238] = 12'h111;
rom[122239] = 12'h  0;
rom[122240] = 12'h  0;
rom[122241] = 12'h  0;
rom[122242] = 12'h  0;
rom[122243] = 12'h  0;
rom[122244] = 12'h  0;
rom[122245] = 12'h  0;
rom[122246] = 12'h  0;
rom[122247] = 12'h  0;
rom[122248] = 12'h  0;
rom[122249] = 12'h  0;
rom[122250] = 12'h  0;
rom[122251] = 12'h  0;
rom[122252] = 12'h  0;
rom[122253] = 12'h  0;
rom[122254] = 12'h  0;
rom[122255] = 12'h  0;
rom[122256] = 12'h  0;
rom[122257] = 12'h  0;
rom[122258] = 12'h  0;
rom[122259] = 12'h  0;
rom[122260] = 12'h  0;
rom[122261] = 12'h  0;
rom[122262] = 12'h333;
rom[122263] = 12'h999;
rom[122264] = 12'heee;
rom[122265] = 12'hccc;
rom[122266] = 12'h666;
rom[122267] = 12'h111;
rom[122268] = 12'h111;
rom[122269] = 12'h  0;
rom[122270] = 12'h  0;
rom[122271] = 12'h  0;
rom[122272] = 12'h  0;
rom[122273] = 12'h  0;
rom[122274] = 12'h  0;
rom[122275] = 12'h  0;
rom[122276] = 12'h  0;
rom[122277] = 12'h111;
rom[122278] = 12'h555;
rom[122279] = 12'haaa;
rom[122280] = 12'haaa;
rom[122281] = 12'h555;
rom[122282] = 12'h222;
rom[122283] = 12'h111;
rom[122284] = 12'h  0;
rom[122285] = 12'h  0;
rom[122286] = 12'h111;
rom[122287] = 12'h  0;
rom[122288] = 12'h  0;
rom[122289] = 12'h  0;
rom[122290] = 12'h  0;
rom[122291] = 12'h  0;
rom[122292] = 12'h111;
rom[122293] = 12'h333;
rom[122294] = 12'h333;
rom[122295] = 12'h111;
rom[122296] = 12'h  0;
rom[122297] = 12'h  0;
rom[122298] = 12'h  0;
rom[122299] = 12'h  0;
rom[122300] = 12'h  0;
rom[122301] = 12'h222;
rom[122302] = 12'h222;
rom[122303] = 12'h222;
rom[122304] = 12'h111;
rom[122305] = 12'h  0;
rom[122306] = 12'h  0;
rom[122307] = 12'h  0;
rom[122308] = 12'h  0;
rom[122309] = 12'h  0;
rom[122310] = 12'h  0;
rom[122311] = 12'h  0;
rom[122312] = 12'h  0;
rom[122313] = 12'h  0;
rom[122314] = 12'h  0;
rom[122315] = 12'h  0;
rom[122316] = 12'h  0;
rom[122317] = 12'h  0;
rom[122318] = 12'h111;
rom[122319] = 12'h222;
rom[122320] = 12'h444;
rom[122321] = 12'h555;
rom[122322] = 12'h555;
rom[122323] = 12'h333;
rom[122324] = 12'h111;
rom[122325] = 12'h  0;
rom[122326] = 12'h  0;
rom[122327] = 12'h  0;
rom[122328] = 12'h  0;
rom[122329] = 12'h  0;
rom[122330] = 12'h  0;
rom[122331] = 12'h  0;
rom[122332] = 12'h  0;
rom[122333] = 12'h  0;
rom[122334] = 12'h  0;
rom[122335] = 12'h  0;
rom[122336] = 12'h  0;
rom[122337] = 12'h  0;
rom[122338] = 12'h  0;
rom[122339] = 12'h  0;
rom[122340] = 12'h  0;
rom[122341] = 12'h  0;
rom[122342] = 12'h  0;
rom[122343] = 12'h  0;
rom[122344] = 12'h  0;
rom[122345] = 12'h  0;
rom[122346] = 12'h  0;
rom[122347] = 12'h  0;
rom[122348] = 12'h  0;
rom[122349] = 12'h  0;
rom[122350] = 12'h  0;
rom[122351] = 12'h  0;
rom[122352] = 12'h  0;
rom[122353] = 12'h  0;
rom[122354] = 12'h  0;
rom[122355] = 12'h  0;
rom[122356] = 12'h  0;
rom[122357] = 12'h  0;
rom[122358] = 12'h  0;
rom[122359] = 12'h  0;
rom[122360] = 12'h  0;
rom[122361] = 12'h  0;
rom[122362] = 12'h  0;
rom[122363] = 12'h  0;
rom[122364] = 12'h  0;
rom[122365] = 12'h  0;
rom[122366] = 12'h  0;
rom[122367] = 12'h  0;
rom[122368] = 12'h  0;
rom[122369] = 12'h  0;
rom[122370] = 12'h  0;
rom[122371] = 12'h  0;
rom[122372] = 12'h  0;
rom[122373] = 12'h  0;
rom[122374] = 12'h  0;
rom[122375] = 12'h111;
rom[122376] = 12'h222;
rom[122377] = 12'h444;
rom[122378] = 12'h666;
rom[122379] = 12'h666;
rom[122380] = 12'h444;
rom[122381] = 12'h222;
rom[122382] = 12'h111;
rom[122383] = 12'h  0;
rom[122384] = 12'h  0;
rom[122385] = 12'h  0;
rom[122386] = 12'h  0;
rom[122387] = 12'h  0;
rom[122388] = 12'h  0;
rom[122389] = 12'h  0;
rom[122390] = 12'h  0;
rom[122391] = 12'h  0;
rom[122392] = 12'h  0;
rom[122393] = 12'h  0;
rom[122394] = 12'h  0;
rom[122395] = 12'h  0;
rom[122396] = 12'h  0;
rom[122397] = 12'h  0;
rom[122398] = 12'h  0;
rom[122399] = 12'h  0;
rom[122400] = 12'heee;
rom[122401] = 12'heee;
rom[122402] = 12'heee;
rom[122403] = 12'heee;
rom[122404] = 12'hddd;
rom[122405] = 12'hddd;
rom[122406] = 12'hddd;
rom[122407] = 12'hddd;
rom[122408] = 12'hddd;
rom[122409] = 12'hddd;
rom[122410] = 12'hddd;
rom[122411] = 12'hddd;
rom[122412] = 12'hddd;
rom[122413] = 12'hddd;
rom[122414] = 12'hddd;
rom[122415] = 12'hddd;
rom[122416] = 12'hddd;
rom[122417] = 12'hddd;
rom[122418] = 12'hddd;
rom[122419] = 12'hccc;
rom[122420] = 12'hccc;
rom[122421] = 12'hccc;
rom[122422] = 12'hccc;
rom[122423] = 12'hccc;
rom[122424] = 12'hccc;
rom[122425] = 12'hccc;
rom[122426] = 12'hccc;
rom[122427] = 12'hccc;
rom[122428] = 12'hccc;
rom[122429] = 12'hccc;
rom[122430] = 12'hccc;
rom[122431] = 12'hbbb;
rom[122432] = 12'hbbb;
rom[122433] = 12'hbbb;
rom[122434] = 12'hbbb;
rom[122435] = 12'hbbb;
rom[122436] = 12'hbbb;
rom[122437] = 12'hbbb;
rom[122438] = 12'hbbb;
rom[122439] = 12'hbbb;
rom[122440] = 12'haaa;
rom[122441] = 12'haaa;
rom[122442] = 12'haaa;
rom[122443] = 12'haaa;
rom[122444] = 12'h999;
rom[122445] = 12'h999;
rom[122446] = 12'h999;
rom[122447] = 12'h999;
rom[122448] = 12'h999;
rom[122449] = 12'h999;
rom[122450] = 12'h999;
rom[122451] = 12'h999;
rom[122452] = 12'h999;
rom[122453] = 12'h999;
rom[122454] = 12'h999;
rom[122455] = 12'h999;
rom[122456] = 12'h999;
rom[122457] = 12'h999;
rom[122458] = 12'h999;
rom[122459] = 12'h999;
rom[122460] = 12'h999;
rom[122461] = 12'h999;
rom[122462] = 12'h999;
rom[122463] = 12'h999;
rom[122464] = 12'h999;
rom[122465] = 12'haaa;
rom[122466] = 12'hccc;
rom[122467] = 12'heee;
rom[122468] = 12'hfff;
rom[122469] = 12'hfff;
rom[122470] = 12'hddd;
rom[122471] = 12'haaa;
rom[122472] = 12'h888;
rom[122473] = 12'h777;
rom[122474] = 12'h666;
rom[122475] = 12'h666;
rom[122476] = 12'h666;
rom[122477] = 12'h666;
rom[122478] = 12'h666;
rom[122479] = 12'h666;
rom[122480] = 12'h666;
rom[122481] = 12'h666;
rom[122482] = 12'h777;
rom[122483] = 12'h777;
rom[122484] = 12'h777;
rom[122485] = 12'h777;
rom[122486] = 12'h777;
rom[122487] = 12'h888;
rom[122488] = 12'hbbb;
rom[122489] = 12'h999;
rom[122490] = 12'h777;
rom[122491] = 12'h555;
rom[122492] = 12'h555;
rom[122493] = 12'h555;
rom[122494] = 12'h555;
rom[122495] = 12'h555;
rom[122496] = 12'h444;
rom[122497] = 12'h555;
rom[122498] = 12'h666;
rom[122499] = 12'h666;
rom[122500] = 12'h555;
rom[122501] = 12'h555;
rom[122502] = 12'h555;
rom[122503] = 12'h666;
rom[122504] = 12'h666;
rom[122505] = 12'h666;
rom[122506] = 12'h666;
rom[122507] = 12'h666;
rom[122508] = 12'h666;
rom[122509] = 12'h666;
rom[122510] = 12'h666;
rom[122511] = 12'h555;
rom[122512] = 12'h555;
rom[122513] = 12'h444;
rom[122514] = 12'h444;
rom[122515] = 12'h444;
rom[122516] = 12'h444;
rom[122517] = 12'h444;
rom[122518] = 12'h555;
rom[122519] = 12'h555;
rom[122520] = 12'h555;
rom[122521] = 12'h444;
rom[122522] = 12'h444;
rom[122523] = 12'h555;
rom[122524] = 12'h555;
rom[122525] = 12'h444;
rom[122526] = 12'h444;
rom[122527] = 12'h444;
rom[122528] = 12'h555;
rom[122529] = 12'h555;
rom[122530] = 12'h555;
rom[122531] = 12'h444;
rom[122532] = 12'h444;
rom[122533] = 12'h444;
rom[122534] = 12'h333;
rom[122535] = 12'h333;
rom[122536] = 12'h333;
rom[122537] = 12'h333;
rom[122538] = 12'h333;
rom[122539] = 12'h333;
rom[122540] = 12'h333;
rom[122541] = 12'h333;
rom[122542] = 12'h222;
rom[122543] = 12'h222;
rom[122544] = 12'h333;
rom[122545] = 12'h333;
rom[122546] = 12'h333;
rom[122547] = 12'h333;
rom[122548] = 12'h333;
rom[122549] = 12'h333;
rom[122550] = 12'h333;
rom[122551] = 12'h333;
rom[122552] = 12'h222;
rom[122553] = 12'h222;
rom[122554] = 12'h222;
rom[122555] = 12'h222;
rom[122556] = 12'h222;
rom[122557] = 12'h222;
rom[122558] = 12'h222;
rom[122559] = 12'h222;
rom[122560] = 12'h222;
rom[122561] = 12'h333;
rom[122562] = 12'h333;
rom[122563] = 12'h333;
rom[122564] = 12'h333;
rom[122565] = 12'h222;
rom[122566] = 12'h222;
rom[122567] = 12'h222;
rom[122568] = 12'h111;
rom[122569] = 12'h111;
rom[122570] = 12'h111;
rom[122571] = 12'h111;
rom[122572] = 12'h111;
rom[122573] = 12'h111;
rom[122574] = 12'h111;
rom[122575] = 12'h111;
rom[122576] = 12'h  0;
rom[122577] = 12'h111;
rom[122578] = 12'h111;
rom[122579] = 12'h111;
rom[122580] = 12'h111;
rom[122581] = 12'h111;
rom[122582] = 12'h111;
rom[122583] = 12'h222;
rom[122584] = 12'h111;
rom[122585] = 12'h111;
rom[122586] = 12'h  0;
rom[122587] = 12'h  0;
rom[122588] = 12'h111;
rom[122589] = 12'h111;
rom[122590] = 12'h111;
rom[122591] = 12'h111;
rom[122592] = 12'h222;
rom[122593] = 12'h222;
rom[122594] = 12'h222;
rom[122595] = 12'h222;
rom[122596] = 12'h222;
rom[122597] = 12'h111;
rom[122598] = 12'h  0;
rom[122599] = 12'h  0;
rom[122600] = 12'h  0;
rom[122601] = 12'h  0;
rom[122602] = 12'h  0;
rom[122603] = 12'h  0;
rom[122604] = 12'h  0;
rom[122605] = 12'h  0;
rom[122606] = 12'h  0;
rom[122607] = 12'h  0;
rom[122608] = 12'h  0;
rom[122609] = 12'h  0;
rom[122610] = 12'h  0;
rom[122611] = 12'h  0;
rom[122612] = 12'h  0;
rom[122613] = 12'h  0;
rom[122614] = 12'h  0;
rom[122615] = 12'h  0;
rom[122616] = 12'h  0;
rom[122617] = 12'h  0;
rom[122618] = 12'h  0;
rom[122619] = 12'h  0;
rom[122620] = 12'h  0;
rom[122621] = 12'h  0;
rom[122622] = 12'h  0;
rom[122623] = 12'h  0;
rom[122624] = 12'h  0;
rom[122625] = 12'h  0;
rom[122626] = 12'h  0;
rom[122627] = 12'h  0;
rom[122628] = 12'h  0;
rom[122629] = 12'h  0;
rom[122630] = 12'h  0;
rom[122631] = 12'h  0;
rom[122632] = 12'h  0;
rom[122633] = 12'h111;
rom[122634] = 12'h222;
rom[122635] = 12'h222;
rom[122636] = 12'h222;
rom[122637] = 12'h111;
rom[122638] = 12'h111;
rom[122639] = 12'h  0;
rom[122640] = 12'h  0;
rom[122641] = 12'h  0;
rom[122642] = 12'h  0;
rom[122643] = 12'h  0;
rom[122644] = 12'h  0;
rom[122645] = 12'h  0;
rom[122646] = 12'h  0;
rom[122647] = 12'h  0;
rom[122648] = 12'h  0;
rom[122649] = 12'h  0;
rom[122650] = 12'h  0;
rom[122651] = 12'h  0;
rom[122652] = 12'h  0;
rom[122653] = 12'h  0;
rom[122654] = 12'h  0;
rom[122655] = 12'h  0;
rom[122656] = 12'h  0;
rom[122657] = 12'h  0;
rom[122658] = 12'h  0;
rom[122659] = 12'h  0;
rom[122660] = 12'h  0;
rom[122661] = 12'h  0;
rom[122662] = 12'h444;
rom[122663] = 12'haaa;
rom[122664] = 12'heee;
rom[122665] = 12'hbbb;
rom[122666] = 12'h555;
rom[122667] = 12'h111;
rom[122668] = 12'h111;
rom[122669] = 12'h  0;
rom[122670] = 12'h  0;
rom[122671] = 12'h  0;
rom[122672] = 12'h  0;
rom[122673] = 12'h  0;
rom[122674] = 12'h  0;
rom[122675] = 12'h  0;
rom[122676] = 12'h  0;
rom[122677] = 12'h111;
rom[122678] = 12'h444;
rom[122679] = 12'h999;
rom[122680] = 12'haaa;
rom[122681] = 12'h666;
rom[122682] = 12'h222;
rom[122683] = 12'h111;
rom[122684] = 12'h  0;
rom[122685] = 12'h  0;
rom[122686] = 12'h  0;
rom[122687] = 12'h  0;
rom[122688] = 12'h  0;
rom[122689] = 12'h  0;
rom[122690] = 12'h  0;
rom[122691] = 12'h  0;
rom[122692] = 12'h111;
rom[122693] = 12'h222;
rom[122694] = 12'h333;
rom[122695] = 12'h111;
rom[122696] = 12'h  0;
rom[122697] = 12'h  0;
rom[122698] = 12'h  0;
rom[122699] = 12'h  0;
rom[122700] = 12'h  0;
rom[122701] = 12'h111;
rom[122702] = 12'h111;
rom[122703] = 12'h222;
rom[122704] = 12'h222;
rom[122705] = 12'h111;
rom[122706] = 12'h  0;
rom[122707] = 12'h  0;
rom[122708] = 12'h  0;
rom[122709] = 12'h  0;
rom[122710] = 12'h  0;
rom[122711] = 12'h  0;
rom[122712] = 12'h  0;
rom[122713] = 12'h  0;
rom[122714] = 12'h  0;
rom[122715] = 12'h  0;
rom[122716] = 12'h  0;
rom[122717] = 12'h  0;
rom[122718] = 12'h111;
rom[122719] = 12'h222;
rom[122720] = 12'h333;
rom[122721] = 12'h555;
rom[122722] = 12'h555;
rom[122723] = 12'h333;
rom[122724] = 12'h111;
rom[122725] = 12'h  0;
rom[122726] = 12'h  0;
rom[122727] = 12'h  0;
rom[122728] = 12'h  0;
rom[122729] = 12'h  0;
rom[122730] = 12'h  0;
rom[122731] = 12'h  0;
rom[122732] = 12'h  0;
rom[122733] = 12'h  0;
rom[122734] = 12'h  0;
rom[122735] = 12'h  0;
rom[122736] = 12'h  0;
rom[122737] = 12'h  0;
rom[122738] = 12'h  0;
rom[122739] = 12'h  0;
rom[122740] = 12'h  0;
rom[122741] = 12'h  0;
rom[122742] = 12'h  0;
rom[122743] = 12'h  0;
rom[122744] = 12'h  0;
rom[122745] = 12'h  0;
rom[122746] = 12'h  0;
rom[122747] = 12'h  0;
rom[122748] = 12'h  0;
rom[122749] = 12'h  0;
rom[122750] = 12'h  0;
rom[122751] = 12'h  0;
rom[122752] = 12'h  0;
rom[122753] = 12'h  0;
rom[122754] = 12'h  0;
rom[122755] = 12'h  0;
rom[122756] = 12'h  0;
rom[122757] = 12'h  0;
rom[122758] = 12'h  0;
rom[122759] = 12'h  0;
rom[122760] = 12'h  0;
rom[122761] = 12'h  0;
rom[122762] = 12'h  0;
rom[122763] = 12'h  0;
rom[122764] = 12'h  0;
rom[122765] = 12'h  0;
rom[122766] = 12'h  0;
rom[122767] = 12'h  0;
rom[122768] = 12'h  0;
rom[122769] = 12'h  0;
rom[122770] = 12'h  0;
rom[122771] = 12'h  0;
rom[122772] = 12'h  0;
rom[122773] = 12'h  0;
rom[122774] = 12'h  0;
rom[122775] = 12'h  0;
rom[122776] = 12'h111;
rom[122777] = 12'h333;
rom[122778] = 12'h666;
rom[122779] = 12'h666;
rom[122780] = 12'h555;
rom[122781] = 12'h333;
rom[122782] = 12'h111;
rom[122783] = 12'h  0;
rom[122784] = 12'h  0;
rom[122785] = 12'h  0;
rom[122786] = 12'h  0;
rom[122787] = 12'h  0;
rom[122788] = 12'h  0;
rom[122789] = 12'h  0;
rom[122790] = 12'h  0;
rom[122791] = 12'h  0;
rom[122792] = 12'h  0;
rom[122793] = 12'h  0;
rom[122794] = 12'h  0;
rom[122795] = 12'h  0;
rom[122796] = 12'h  0;
rom[122797] = 12'h  0;
rom[122798] = 12'h  0;
rom[122799] = 12'h  0;
rom[122800] = 12'heee;
rom[122801] = 12'heee;
rom[122802] = 12'heee;
rom[122803] = 12'hddd;
rom[122804] = 12'hddd;
rom[122805] = 12'hddd;
rom[122806] = 12'hddd;
rom[122807] = 12'hddd;
rom[122808] = 12'hddd;
rom[122809] = 12'hddd;
rom[122810] = 12'hddd;
rom[122811] = 12'hddd;
rom[122812] = 12'hddd;
rom[122813] = 12'hddd;
rom[122814] = 12'hddd;
rom[122815] = 12'hddd;
rom[122816] = 12'hddd;
rom[122817] = 12'hddd;
rom[122818] = 12'hccc;
rom[122819] = 12'hccc;
rom[122820] = 12'hccc;
rom[122821] = 12'hccc;
rom[122822] = 12'hccc;
rom[122823] = 12'hccc;
rom[122824] = 12'hccc;
rom[122825] = 12'hccc;
rom[122826] = 12'hccc;
rom[122827] = 12'hbbb;
rom[122828] = 12'hbbb;
rom[122829] = 12'hbbb;
rom[122830] = 12'hbbb;
rom[122831] = 12'hbbb;
rom[122832] = 12'hbbb;
rom[122833] = 12'hbbb;
rom[122834] = 12'hbbb;
rom[122835] = 12'hbbb;
rom[122836] = 12'hbbb;
rom[122837] = 12'haaa;
rom[122838] = 12'haaa;
rom[122839] = 12'haaa;
rom[122840] = 12'haaa;
rom[122841] = 12'haaa;
rom[122842] = 12'h999;
rom[122843] = 12'h999;
rom[122844] = 12'h999;
rom[122845] = 12'h999;
rom[122846] = 12'h999;
rom[122847] = 12'h999;
rom[122848] = 12'h999;
rom[122849] = 12'h888;
rom[122850] = 12'h888;
rom[122851] = 12'h888;
rom[122852] = 12'h888;
rom[122853] = 12'h888;
rom[122854] = 12'h888;
rom[122855] = 12'h888;
rom[122856] = 12'h888;
rom[122857] = 12'h888;
rom[122858] = 12'h999;
rom[122859] = 12'h999;
rom[122860] = 12'h999;
rom[122861] = 12'h999;
rom[122862] = 12'h999;
rom[122863] = 12'h999;
rom[122864] = 12'h999;
rom[122865] = 12'hbbb;
rom[122866] = 12'heee;
rom[122867] = 12'hfff;
rom[122868] = 12'hfff;
rom[122869] = 12'heee;
rom[122870] = 12'hbbb;
rom[122871] = 12'h999;
rom[122872] = 12'h777;
rom[122873] = 12'h777;
rom[122874] = 12'h666;
rom[122875] = 12'h666;
rom[122876] = 12'h666;
rom[122877] = 12'h666;
rom[122878] = 12'h666;
rom[122879] = 12'h666;
rom[122880] = 12'h666;
rom[122881] = 12'h666;
rom[122882] = 12'h777;
rom[122883] = 12'h777;
rom[122884] = 12'h777;
rom[122885] = 12'h777;
rom[122886] = 12'h999;
rom[122887] = 12'h999;
rom[122888] = 12'haaa;
rom[122889] = 12'h777;
rom[122890] = 12'h555;
rom[122891] = 12'h555;
rom[122892] = 12'h555;
rom[122893] = 12'h555;
rom[122894] = 12'h444;
rom[122895] = 12'h444;
rom[122896] = 12'h444;
rom[122897] = 12'h555;
rom[122898] = 12'h666;
rom[122899] = 12'h666;
rom[122900] = 12'h555;
rom[122901] = 12'h555;
rom[122902] = 12'h555;
rom[122903] = 12'h555;
rom[122904] = 12'h666;
rom[122905] = 12'h666;
rom[122906] = 12'h666;
rom[122907] = 12'h666;
rom[122908] = 12'h666;
rom[122909] = 12'h666;
rom[122910] = 12'h555;
rom[122911] = 12'h555;
rom[122912] = 12'h555;
rom[122913] = 12'h444;
rom[122914] = 12'h444;
rom[122915] = 12'h444;
rom[122916] = 12'h444;
rom[122917] = 12'h444;
rom[122918] = 12'h555;
rom[122919] = 12'h555;
rom[122920] = 12'h444;
rom[122921] = 12'h444;
rom[122922] = 12'h444;
rom[122923] = 12'h555;
rom[122924] = 12'h444;
rom[122925] = 12'h444;
rom[122926] = 12'h444;
rom[122927] = 12'h444;
rom[122928] = 12'h444;
rom[122929] = 12'h555;
rom[122930] = 12'h555;
rom[122931] = 12'h555;
rom[122932] = 12'h444;
rom[122933] = 12'h444;
rom[122934] = 12'h333;
rom[122935] = 12'h333;
rom[122936] = 12'h333;
rom[122937] = 12'h333;
rom[122938] = 12'h333;
rom[122939] = 12'h333;
rom[122940] = 12'h333;
rom[122941] = 12'h333;
rom[122942] = 12'h222;
rom[122943] = 12'h222;
rom[122944] = 12'h333;
rom[122945] = 12'h333;
rom[122946] = 12'h333;
rom[122947] = 12'h333;
rom[122948] = 12'h333;
rom[122949] = 12'h333;
rom[122950] = 12'h333;
rom[122951] = 12'h333;
rom[122952] = 12'h222;
rom[122953] = 12'h222;
rom[122954] = 12'h222;
rom[122955] = 12'h222;
rom[122956] = 12'h222;
rom[122957] = 12'h222;
rom[122958] = 12'h222;
rom[122959] = 12'h333;
rom[122960] = 12'h222;
rom[122961] = 12'h222;
rom[122962] = 12'h333;
rom[122963] = 12'h333;
rom[122964] = 12'h222;
rom[122965] = 12'h222;
rom[122966] = 12'h111;
rom[122967] = 12'h111;
rom[122968] = 12'h111;
rom[122969] = 12'h111;
rom[122970] = 12'h111;
rom[122971] = 12'h111;
rom[122972] = 12'h111;
rom[122973] = 12'h111;
rom[122974] = 12'h111;
rom[122975] = 12'h111;
rom[122976] = 12'h  0;
rom[122977] = 12'h  0;
rom[122978] = 12'h  0;
rom[122979] = 12'h111;
rom[122980] = 12'h111;
rom[122981] = 12'h111;
rom[122982] = 12'h111;
rom[122983] = 12'h111;
rom[122984] = 12'h111;
rom[122985] = 12'h111;
rom[122986] = 12'h  0;
rom[122987] = 12'h  0;
rom[122988] = 12'h111;
rom[122989] = 12'h111;
rom[122990] = 12'h111;
rom[122991] = 12'h111;
rom[122992] = 12'h111;
rom[122993] = 12'h111;
rom[122994] = 12'h111;
rom[122995] = 12'h111;
rom[122996] = 12'h111;
rom[122997] = 12'h111;
rom[122998] = 12'h  0;
rom[122999] = 12'h  0;
rom[123000] = 12'h  0;
rom[123001] = 12'h  0;
rom[123002] = 12'h  0;
rom[123003] = 12'h  0;
rom[123004] = 12'h  0;
rom[123005] = 12'h  0;
rom[123006] = 12'h  0;
rom[123007] = 12'h  0;
rom[123008] = 12'h  0;
rom[123009] = 12'h  0;
rom[123010] = 12'h  0;
rom[123011] = 12'h  0;
rom[123012] = 12'h  0;
rom[123013] = 12'h  0;
rom[123014] = 12'h  0;
rom[123015] = 12'h  0;
rom[123016] = 12'h  0;
rom[123017] = 12'h  0;
rom[123018] = 12'h  0;
rom[123019] = 12'h  0;
rom[123020] = 12'h  0;
rom[123021] = 12'h  0;
rom[123022] = 12'h  0;
rom[123023] = 12'h  0;
rom[123024] = 12'h  0;
rom[123025] = 12'h  0;
rom[123026] = 12'h  0;
rom[123027] = 12'h  0;
rom[123028] = 12'h  0;
rom[123029] = 12'h  0;
rom[123030] = 12'h  0;
rom[123031] = 12'h  0;
rom[123032] = 12'h  0;
rom[123033] = 12'h111;
rom[123034] = 12'h222;
rom[123035] = 12'h222;
rom[123036] = 12'h111;
rom[123037] = 12'h111;
rom[123038] = 12'h111;
rom[123039] = 12'h  0;
rom[123040] = 12'h  0;
rom[123041] = 12'h  0;
rom[123042] = 12'h  0;
rom[123043] = 12'h  0;
rom[123044] = 12'h  0;
rom[123045] = 12'h  0;
rom[123046] = 12'h  0;
rom[123047] = 12'h  0;
rom[123048] = 12'h  0;
rom[123049] = 12'h  0;
rom[123050] = 12'h  0;
rom[123051] = 12'h  0;
rom[123052] = 12'h  0;
rom[123053] = 12'h  0;
rom[123054] = 12'h  0;
rom[123055] = 12'h  0;
rom[123056] = 12'h  0;
rom[123057] = 12'h  0;
rom[123058] = 12'h  0;
rom[123059] = 12'h  0;
rom[123060] = 12'h  0;
rom[123061] = 12'h  0;
rom[123062] = 12'h555;
rom[123063] = 12'hbbb;
rom[123064] = 12'heee;
rom[123065] = 12'haaa;
rom[123066] = 12'h444;
rom[123067] = 12'h111;
rom[123068] = 12'h111;
rom[123069] = 12'h111;
rom[123070] = 12'h  0;
rom[123071] = 12'h  0;
rom[123072] = 12'h  0;
rom[123073] = 12'h  0;
rom[123074] = 12'h  0;
rom[123075] = 12'h  0;
rom[123076] = 12'h  0;
rom[123077] = 12'h111;
rom[123078] = 12'h444;
rom[123079] = 12'h888;
rom[123080] = 12'haaa;
rom[123081] = 12'h666;
rom[123082] = 12'h222;
rom[123083] = 12'h  0;
rom[123084] = 12'h  0;
rom[123085] = 12'h  0;
rom[123086] = 12'h  0;
rom[123087] = 12'h  0;
rom[123088] = 12'h  0;
rom[123089] = 12'h  0;
rom[123090] = 12'h  0;
rom[123091] = 12'h  0;
rom[123092] = 12'h111;
rom[123093] = 12'h222;
rom[123094] = 12'h222;
rom[123095] = 12'h111;
rom[123096] = 12'h  0;
rom[123097] = 12'h  0;
rom[123098] = 12'h  0;
rom[123099] = 12'h  0;
rom[123100] = 12'h  0;
rom[123101] = 12'h  0;
rom[123102] = 12'h111;
rom[123103] = 12'h111;
rom[123104] = 12'h222;
rom[123105] = 12'h111;
rom[123106] = 12'h  0;
rom[123107] = 12'h  0;
rom[123108] = 12'h  0;
rom[123109] = 12'h  0;
rom[123110] = 12'h  0;
rom[123111] = 12'h  0;
rom[123112] = 12'h  0;
rom[123113] = 12'h  0;
rom[123114] = 12'h  0;
rom[123115] = 12'h  0;
rom[123116] = 12'h  0;
rom[123117] = 12'h  0;
rom[123118] = 12'h  0;
rom[123119] = 12'h111;
rom[123120] = 12'h333;
rom[123121] = 12'h444;
rom[123122] = 12'h555;
rom[123123] = 12'h333;
rom[123124] = 12'h111;
rom[123125] = 12'h  0;
rom[123126] = 12'h  0;
rom[123127] = 12'h  0;
rom[123128] = 12'h  0;
rom[123129] = 12'h  0;
rom[123130] = 12'h  0;
rom[123131] = 12'h  0;
rom[123132] = 12'h  0;
rom[123133] = 12'h  0;
rom[123134] = 12'h  0;
rom[123135] = 12'h  0;
rom[123136] = 12'h  0;
rom[123137] = 12'h  0;
rom[123138] = 12'h  0;
rom[123139] = 12'h  0;
rom[123140] = 12'h  0;
rom[123141] = 12'h  0;
rom[123142] = 12'h  0;
rom[123143] = 12'h  0;
rom[123144] = 12'h  0;
rom[123145] = 12'h  0;
rom[123146] = 12'h  0;
rom[123147] = 12'h  0;
rom[123148] = 12'h  0;
rom[123149] = 12'h  0;
rom[123150] = 12'h  0;
rom[123151] = 12'h  0;
rom[123152] = 12'h  0;
rom[123153] = 12'h  0;
rom[123154] = 12'h  0;
rom[123155] = 12'h  0;
rom[123156] = 12'h  0;
rom[123157] = 12'h  0;
rom[123158] = 12'h  0;
rom[123159] = 12'h  0;
rom[123160] = 12'h  0;
rom[123161] = 12'h  0;
rom[123162] = 12'h  0;
rom[123163] = 12'h  0;
rom[123164] = 12'h  0;
rom[123165] = 12'h  0;
rom[123166] = 12'h  0;
rom[123167] = 12'h  0;
rom[123168] = 12'h  0;
rom[123169] = 12'h  0;
rom[123170] = 12'h  0;
rom[123171] = 12'h  0;
rom[123172] = 12'h  0;
rom[123173] = 12'h  0;
rom[123174] = 12'h  0;
rom[123175] = 12'h  0;
rom[123176] = 12'h111;
rom[123177] = 12'h333;
rom[123178] = 12'h555;
rom[123179] = 12'h666;
rom[123180] = 12'h555;
rom[123181] = 12'h444;
rom[123182] = 12'h111;
rom[123183] = 12'h  0;
rom[123184] = 12'h  0;
rom[123185] = 12'h  0;
rom[123186] = 12'h  0;
rom[123187] = 12'h  0;
rom[123188] = 12'h  0;
rom[123189] = 12'h  0;
rom[123190] = 12'h  0;
rom[123191] = 12'h  0;
rom[123192] = 12'h  0;
rom[123193] = 12'h  0;
rom[123194] = 12'h  0;
rom[123195] = 12'h  0;
rom[123196] = 12'h  0;
rom[123197] = 12'h  0;
rom[123198] = 12'h  0;
rom[123199] = 12'h  0;
rom[123200] = 12'heee;
rom[123201] = 12'heee;
rom[123202] = 12'hddd;
rom[123203] = 12'hddd;
rom[123204] = 12'hddd;
rom[123205] = 12'hddd;
rom[123206] = 12'hddd;
rom[123207] = 12'hddd;
rom[123208] = 12'hddd;
rom[123209] = 12'hddd;
rom[123210] = 12'hddd;
rom[123211] = 12'hddd;
rom[123212] = 12'hccc;
rom[123213] = 12'hccc;
rom[123214] = 12'hccc;
rom[123215] = 12'hccc;
rom[123216] = 12'hccc;
rom[123217] = 12'hccc;
rom[123218] = 12'hccc;
rom[123219] = 12'hccc;
rom[123220] = 12'hccc;
rom[123221] = 12'hccc;
rom[123222] = 12'hccc;
rom[123223] = 12'hccc;
rom[123224] = 12'hccc;
rom[123225] = 12'hbbb;
rom[123226] = 12'hbbb;
rom[123227] = 12'hbbb;
rom[123228] = 12'hbbb;
rom[123229] = 12'hbbb;
rom[123230] = 12'hbbb;
rom[123231] = 12'hbbb;
rom[123232] = 12'haaa;
rom[123233] = 12'haaa;
rom[123234] = 12'haaa;
rom[123235] = 12'haaa;
rom[123236] = 12'haaa;
rom[123237] = 12'haaa;
rom[123238] = 12'haaa;
rom[123239] = 12'h999;
rom[123240] = 12'h999;
rom[123241] = 12'h999;
rom[123242] = 12'h999;
rom[123243] = 12'h999;
rom[123244] = 12'h999;
rom[123245] = 12'h888;
rom[123246] = 12'h888;
rom[123247] = 12'h888;
rom[123248] = 12'h888;
rom[123249] = 12'h888;
rom[123250] = 12'h888;
rom[123251] = 12'h888;
rom[123252] = 12'h777;
rom[123253] = 12'h888;
rom[123254] = 12'h888;
rom[123255] = 12'h888;
rom[123256] = 12'h888;
rom[123257] = 12'h888;
rom[123258] = 12'h888;
rom[123259] = 12'h999;
rom[123260] = 12'h999;
rom[123261] = 12'h999;
rom[123262] = 12'h999;
rom[123263] = 12'h999;
rom[123264] = 12'haaa;
rom[123265] = 12'hddd;
rom[123266] = 12'hfff;
rom[123267] = 12'hfff;
rom[123268] = 12'heee;
rom[123269] = 12'hbbb;
rom[123270] = 12'h999;
rom[123271] = 12'h777;
rom[123272] = 12'h666;
rom[123273] = 12'h666;
rom[123274] = 12'h666;
rom[123275] = 12'h666;
rom[123276] = 12'h666;
rom[123277] = 12'h666;
rom[123278] = 12'h666;
rom[123279] = 12'h555;
rom[123280] = 12'h666;
rom[123281] = 12'h666;
rom[123282] = 12'h666;
rom[123283] = 12'h666;
rom[123284] = 12'h777;
rom[123285] = 12'h888;
rom[123286] = 12'h999;
rom[123287] = 12'haaa;
rom[123288] = 12'h888;
rom[123289] = 12'h666;
rom[123290] = 12'h555;
rom[123291] = 12'h555;
rom[123292] = 12'h555;
rom[123293] = 12'h555;
rom[123294] = 12'h444;
rom[123295] = 12'h444;
rom[123296] = 12'h444;
rom[123297] = 12'h555;
rom[123298] = 12'h666;
rom[123299] = 12'h555;
rom[123300] = 12'h555;
rom[123301] = 12'h444;
rom[123302] = 12'h555;
rom[123303] = 12'h555;
rom[123304] = 12'h555;
rom[123305] = 12'h555;
rom[123306] = 12'h666;
rom[123307] = 12'h666;
rom[123308] = 12'h666;
rom[123309] = 12'h666;
rom[123310] = 12'h555;
rom[123311] = 12'h555;
rom[123312] = 12'h555;
rom[123313] = 12'h444;
rom[123314] = 12'h444;
rom[123315] = 12'h444;
rom[123316] = 12'h444;
rom[123317] = 12'h555;
rom[123318] = 12'h555;
rom[123319] = 12'h555;
rom[123320] = 12'h444;
rom[123321] = 12'h444;
rom[123322] = 12'h444;
rom[123323] = 12'h555;
rom[123324] = 12'h444;
rom[123325] = 12'h444;
rom[123326] = 12'h444;
rom[123327] = 12'h444;
rom[123328] = 12'h444;
rom[123329] = 12'h444;
rom[123330] = 12'h555;
rom[123331] = 12'h555;
rom[123332] = 12'h555;
rom[123333] = 12'h444;
rom[123334] = 12'h333;
rom[123335] = 12'h333;
rom[123336] = 12'h333;
rom[123337] = 12'h333;
rom[123338] = 12'h333;
rom[123339] = 12'h333;
rom[123340] = 12'h333;
rom[123341] = 12'h333;
rom[123342] = 12'h222;
rom[123343] = 12'h222;
rom[123344] = 12'h222;
rom[123345] = 12'h333;
rom[123346] = 12'h333;
rom[123347] = 12'h333;
rom[123348] = 12'h333;
rom[123349] = 12'h333;
rom[123350] = 12'h333;
rom[123351] = 12'h333;
rom[123352] = 12'h222;
rom[123353] = 12'h222;
rom[123354] = 12'h222;
rom[123355] = 12'h222;
rom[123356] = 12'h222;
rom[123357] = 12'h222;
rom[123358] = 12'h222;
rom[123359] = 12'h333;
rom[123360] = 12'h222;
rom[123361] = 12'h222;
rom[123362] = 12'h222;
rom[123363] = 12'h222;
rom[123364] = 12'h222;
rom[123365] = 12'h222;
rom[123366] = 12'h111;
rom[123367] = 12'h111;
rom[123368] = 12'h111;
rom[123369] = 12'h111;
rom[123370] = 12'h111;
rom[123371] = 12'h111;
rom[123372] = 12'h111;
rom[123373] = 12'h111;
rom[123374] = 12'h111;
rom[123375] = 12'h  0;
rom[123376] = 12'h  0;
rom[123377] = 12'h  0;
rom[123378] = 12'h  0;
rom[123379] = 12'h  0;
rom[123380] = 12'h111;
rom[123381] = 12'h111;
rom[123382] = 12'h111;
rom[123383] = 12'h111;
rom[123384] = 12'h111;
rom[123385] = 12'h111;
rom[123386] = 12'h111;
rom[123387] = 12'h  0;
rom[123388] = 12'h111;
rom[123389] = 12'h111;
rom[123390] = 12'h111;
rom[123391] = 12'h111;
rom[123392] = 12'h111;
rom[123393] = 12'h111;
rom[123394] = 12'h111;
rom[123395] = 12'h111;
rom[123396] = 12'h111;
rom[123397] = 12'h111;
rom[123398] = 12'h  0;
rom[123399] = 12'h  0;
rom[123400] = 12'h  0;
rom[123401] = 12'h  0;
rom[123402] = 12'h  0;
rom[123403] = 12'h  0;
rom[123404] = 12'h  0;
rom[123405] = 12'h  0;
rom[123406] = 12'h  0;
rom[123407] = 12'h  0;
rom[123408] = 12'h  0;
rom[123409] = 12'h  0;
rom[123410] = 12'h  0;
rom[123411] = 12'h  0;
rom[123412] = 12'h  0;
rom[123413] = 12'h  0;
rom[123414] = 12'h  0;
rom[123415] = 12'h  0;
rom[123416] = 12'h  0;
rom[123417] = 12'h  0;
rom[123418] = 12'h  0;
rom[123419] = 12'h  0;
rom[123420] = 12'h  0;
rom[123421] = 12'h  0;
rom[123422] = 12'h  0;
rom[123423] = 12'h  0;
rom[123424] = 12'h  0;
rom[123425] = 12'h  0;
rom[123426] = 12'h  0;
rom[123427] = 12'h  0;
rom[123428] = 12'h  0;
rom[123429] = 12'h  0;
rom[123430] = 12'h  0;
rom[123431] = 12'h  0;
rom[123432] = 12'h  0;
rom[123433] = 12'h111;
rom[123434] = 12'h222;
rom[123435] = 12'h111;
rom[123436] = 12'h  0;
rom[123437] = 12'h  0;
rom[123438] = 12'h111;
rom[123439] = 12'h  0;
rom[123440] = 12'h  0;
rom[123441] = 12'h  0;
rom[123442] = 12'h  0;
rom[123443] = 12'h  0;
rom[123444] = 12'h  0;
rom[123445] = 12'h  0;
rom[123446] = 12'h  0;
rom[123447] = 12'h  0;
rom[123448] = 12'h  0;
rom[123449] = 12'h  0;
rom[123450] = 12'h  0;
rom[123451] = 12'h  0;
rom[123452] = 12'h  0;
rom[123453] = 12'h  0;
rom[123454] = 12'h  0;
rom[123455] = 12'h  0;
rom[123456] = 12'h  0;
rom[123457] = 12'h  0;
rom[123458] = 12'h  0;
rom[123459] = 12'h  0;
rom[123460] = 12'h  0;
rom[123461] = 12'h111;
rom[123462] = 12'h555;
rom[123463] = 12'hbbb;
rom[123464] = 12'heee;
rom[123465] = 12'h999;
rom[123466] = 12'h444;
rom[123467] = 12'h111;
rom[123468] = 12'h111;
rom[123469] = 12'h111;
rom[123470] = 12'h  0;
rom[123471] = 12'h  0;
rom[123472] = 12'h  0;
rom[123473] = 12'h  0;
rom[123474] = 12'h  0;
rom[123475] = 12'h  0;
rom[123476] = 12'h  0;
rom[123477] = 12'h111;
rom[123478] = 12'h333;
rom[123479] = 12'h777;
rom[123480] = 12'haaa;
rom[123481] = 12'h777;
rom[123482] = 12'h222;
rom[123483] = 12'h  0;
rom[123484] = 12'h  0;
rom[123485] = 12'h  0;
rom[123486] = 12'h  0;
rom[123487] = 12'h  0;
rom[123488] = 12'h  0;
rom[123489] = 12'h  0;
rom[123490] = 12'h  0;
rom[123491] = 12'h  0;
rom[123492] = 12'h  0;
rom[123493] = 12'h222;
rom[123494] = 12'h222;
rom[123495] = 12'h111;
rom[123496] = 12'h  0;
rom[123497] = 12'h  0;
rom[123498] = 12'h  0;
rom[123499] = 12'h  0;
rom[123500] = 12'h  0;
rom[123501] = 12'h  0;
rom[123502] = 12'h  0;
rom[123503] = 12'h111;
rom[123504] = 12'h222;
rom[123505] = 12'h222;
rom[123506] = 12'h111;
rom[123507] = 12'h  0;
rom[123508] = 12'h  0;
rom[123509] = 12'h  0;
rom[123510] = 12'h  0;
rom[123511] = 12'h  0;
rom[123512] = 12'h  0;
rom[123513] = 12'h  0;
rom[123514] = 12'h  0;
rom[123515] = 12'h  0;
rom[123516] = 12'h  0;
rom[123517] = 12'h  0;
rom[123518] = 12'h  0;
rom[123519] = 12'h111;
rom[123520] = 12'h333;
rom[123521] = 12'h444;
rom[123522] = 12'h555;
rom[123523] = 12'h444;
rom[123524] = 12'h222;
rom[123525] = 12'h  0;
rom[123526] = 12'h  0;
rom[123527] = 12'h  0;
rom[123528] = 12'h  0;
rom[123529] = 12'h  0;
rom[123530] = 12'h  0;
rom[123531] = 12'h  0;
rom[123532] = 12'h  0;
rom[123533] = 12'h  0;
rom[123534] = 12'h  0;
rom[123535] = 12'h  0;
rom[123536] = 12'h  0;
rom[123537] = 12'h  0;
rom[123538] = 12'h  0;
rom[123539] = 12'h  0;
rom[123540] = 12'h  0;
rom[123541] = 12'h  0;
rom[123542] = 12'h  0;
rom[123543] = 12'h  0;
rom[123544] = 12'h  0;
rom[123545] = 12'h  0;
rom[123546] = 12'h  0;
rom[123547] = 12'h  0;
rom[123548] = 12'h  0;
rom[123549] = 12'h  0;
rom[123550] = 12'h  0;
rom[123551] = 12'h  0;
rom[123552] = 12'h  0;
rom[123553] = 12'h  0;
rom[123554] = 12'h  0;
rom[123555] = 12'h  0;
rom[123556] = 12'h  0;
rom[123557] = 12'h  0;
rom[123558] = 12'h  0;
rom[123559] = 12'h  0;
rom[123560] = 12'h  0;
rom[123561] = 12'h  0;
rom[123562] = 12'h  0;
rom[123563] = 12'h  0;
rom[123564] = 12'h  0;
rom[123565] = 12'h  0;
rom[123566] = 12'h  0;
rom[123567] = 12'h  0;
rom[123568] = 12'h  0;
rom[123569] = 12'h  0;
rom[123570] = 12'h  0;
rom[123571] = 12'h  0;
rom[123572] = 12'h  0;
rom[123573] = 12'h  0;
rom[123574] = 12'h  0;
rom[123575] = 12'h  0;
rom[123576] = 12'h111;
rom[123577] = 12'h222;
rom[123578] = 12'h444;
rom[123579] = 12'h555;
rom[123580] = 12'h666;
rom[123581] = 12'h444;
rom[123582] = 12'h222;
rom[123583] = 12'h111;
rom[123584] = 12'h  0;
rom[123585] = 12'h  0;
rom[123586] = 12'h  0;
rom[123587] = 12'h  0;
rom[123588] = 12'h  0;
rom[123589] = 12'h  0;
rom[123590] = 12'h  0;
rom[123591] = 12'h  0;
rom[123592] = 12'h  0;
rom[123593] = 12'h  0;
rom[123594] = 12'h  0;
rom[123595] = 12'h  0;
rom[123596] = 12'h  0;
rom[123597] = 12'h  0;
rom[123598] = 12'h  0;
rom[123599] = 12'h  0;
rom[123600] = 12'hddd;
rom[123601] = 12'hddd;
rom[123602] = 12'hddd;
rom[123603] = 12'hddd;
rom[123604] = 12'hddd;
rom[123605] = 12'hddd;
rom[123606] = 12'hddd;
rom[123607] = 12'hddd;
rom[123608] = 12'hddd;
rom[123609] = 12'hddd;
rom[123610] = 12'hddd;
rom[123611] = 12'hccc;
rom[123612] = 12'hccc;
rom[123613] = 12'hccc;
rom[123614] = 12'hccc;
rom[123615] = 12'hccc;
rom[123616] = 12'hccc;
rom[123617] = 12'hccc;
rom[123618] = 12'hccc;
rom[123619] = 12'hccc;
rom[123620] = 12'hccc;
rom[123621] = 12'hccc;
rom[123622] = 12'hbbb;
rom[123623] = 12'hbbb;
rom[123624] = 12'hbbb;
rom[123625] = 12'hbbb;
rom[123626] = 12'hbbb;
rom[123627] = 12'hbbb;
rom[123628] = 12'hbbb;
rom[123629] = 12'hbbb;
rom[123630] = 12'haaa;
rom[123631] = 12'haaa;
rom[123632] = 12'haaa;
rom[123633] = 12'haaa;
rom[123634] = 12'haaa;
rom[123635] = 12'haaa;
rom[123636] = 12'haaa;
rom[123637] = 12'h999;
rom[123638] = 12'h999;
rom[123639] = 12'h999;
rom[123640] = 12'h999;
rom[123641] = 12'h999;
rom[123642] = 12'h888;
rom[123643] = 12'h888;
rom[123644] = 12'h888;
rom[123645] = 12'h888;
rom[123646] = 12'h888;
rom[123647] = 12'h888;
rom[123648] = 12'h888;
rom[123649] = 12'h888;
rom[123650] = 12'h888;
rom[123651] = 12'h777;
rom[123652] = 12'h777;
rom[123653] = 12'h777;
rom[123654] = 12'h777;
rom[123655] = 12'h777;
rom[123656] = 12'h888;
rom[123657] = 12'h777;
rom[123658] = 12'h888;
rom[123659] = 12'h888;
rom[123660] = 12'h999;
rom[123661] = 12'h888;
rom[123662] = 12'h999;
rom[123663] = 12'h999;
rom[123664] = 12'hbbb;
rom[123665] = 12'heee;
rom[123666] = 12'hfff;
rom[123667] = 12'hfff;
rom[123668] = 12'hccc;
rom[123669] = 12'h999;
rom[123670] = 12'h888;
rom[123671] = 12'h666;
rom[123672] = 12'h666;
rom[123673] = 12'h666;
rom[123674] = 12'h666;
rom[123675] = 12'h666;
rom[123676] = 12'h666;
rom[123677] = 12'h666;
rom[123678] = 12'h555;
rom[123679] = 12'h555;
rom[123680] = 12'h666;
rom[123681] = 12'h666;
rom[123682] = 12'h666;
rom[123683] = 12'h666;
rom[123684] = 12'h777;
rom[123685] = 12'h999;
rom[123686] = 12'h999;
rom[123687] = 12'h999;
rom[123688] = 12'h666;
rom[123689] = 12'h555;
rom[123690] = 12'h555;
rom[123691] = 12'h555;
rom[123692] = 12'h555;
rom[123693] = 12'h444;
rom[123694] = 12'h444;
rom[123695] = 12'h555;
rom[123696] = 12'h444;
rom[123697] = 12'h555;
rom[123698] = 12'h555;
rom[123699] = 12'h555;
rom[123700] = 12'h555;
rom[123701] = 12'h444;
rom[123702] = 12'h444;
rom[123703] = 12'h555;
rom[123704] = 12'h555;
rom[123705] = 12'h555;
rom[123706] = 12'h555;
rom[123707] = 12'h666;
rom[123708] = 12'h666;
rom[123709] = 12'h666;
rom[123710] = 12'h555;
rom[123711] = 12'h555;
rom[123712] = 12'h555;
rom[123713] = 12'h555;
rom[123714] = 12'h444;
rom[123715] = 12'h444;
rom[123716] = 12'h444;
rom[123717] = 12'h555;
rom[123718] = 12'h555;
rom[123719] = 12'h555;
rom[123720] = 12'h444;
rom[123721] = 12'h444;
rom[123722] = 12'h444;
rom[123723] = 12'h555;
rom[123724] = 12'h444;
rom[123725] = 12'h444;
rom[123726] = 12'h444;
rom[123727] = 12'h444;
rom[123728] = 12'h444;
rom[123729] = 12'h444;
rom[123730] = 12'h444;
rom[123731] = 12'h555;
rom[123732] = 12'h555;
rom[123733] = 12'h444;
rom[123734] = 12'h444;
rom[123735] = 12'h333;
rom[123736] = 12'h333;
rom[123737] = 12'h333;
rom[123738] = 12'h333;
rom[123739] = 12'h333;
rom[123740] = 12'h333;
rom[123741] = 12'h333;
rom[123742] = 12'h222;
rom[123743] = 12'h222;
rom[123744] = 12'h222;
rom[123745] = 12'h222;
rom[123746] = 12'h333;
rom[123747] = 12'h333;
rom[123748] = 12'h333;
rom[123749] = 12'h333;
rom[123750] = 12'h333;
rom[123751] = 12'h333;
rom[123752] = 12'h222;
rom[123753] = 12'h222;
rom[123754] = 12'h222;
rom[123755] = 12'h222;
rom[123756] = 12'h222;
rom[123757] = 12'h222;
rom[123758] = 12'h222;
rom[123759] = 12'h222;
rom[123760] = 12'h222;
rom[123761] = 12'h222;
rom[123762] = 12'h222;
rom[123763] = 12'h222;
rom[123764] = 12'h222;
rom[123765] = 12'h111;
rom[123766] = 12'h111;
rom[123767] = 12'h111;
rom[123768] = 12'h111;
rom[123769] = 12'h111;
rom[123770] = 12'h111;
rom[123771] = 12'h111;
rom[123772] = 12'h111;
rom[123773] = 12'h111;
rom[123774] = 12'h111;
rom[123775] = 12'h  0;
rom[123776] = 12'h  0;
rom[123777] = 12'h  0;
rom[123778] = 12'h  0;
rom[123779] = 12'h  0;
rom[123780] = 12'h  0;
rom[123781] = 12'h111;
rom[123782] = 12'h111;
rom[123783] = 12'h111;
rom[123784] = 12'h111;
rom[123785] = 12'h111;
rom[123786] = 12'h111;
rom[123787] = 12'h111;
rom[123788] = 12'h111;
rom[123789] = 12'h111;
rom[123790] = 12'h111;
rom[123791] = 12'h111;
rom[123792] = 12'h111;
rom[123793] = 12'h111;
rom[123794] = 12'h111;
rom[123795] = 12'h111;
rom[123796] = 12'h111;
rom[123797] = 12'h111;
rom[123798] = 12'h  0;
rom[123799] = 12'h  0;
rom[123800] = 12'h  0;
rom[123801] = 12'h  0;
rom[123802] = 12'h  0;
rom[123803] = 12'h  0;
rom[123804] = 12'h  0;
rom[123805] = 12'h  0;
rom[123806] = 12'h  0;
rom[123807] = 12'h  0;
rom[123808] = 12'h  0;
rom[123809] = 12'h  0;
rom[123810] = 12'h  0;
rom[123811] = 12'h  0;
rom[123812] = 12'h  0;
rom[123813] = 12'h  0;
rom[123814] = 12'h  0;
rom[123815] = 12'h  0;
rom[123816] = 12'h  0;
rom[123817] = 12'h  0;
rom[123818] = 12'h  0;
rom[123819] = 12'h  0;
rom[123820] = 12'h  0;
rom[123821] = 12'h  0;
rom[123822] = 12'h  0;
rom[123823] = 12'h  0;
rom[123824] = 12'h  0;
rom[123825] = 12'h  0;
rom[123826] = 12'h  0;
rom[123827] = 12'h  0;
rom[123828] = 12'h  0;
rom[123829] = 12'h  0;
rom[123830] = 12'h  0;
rom[123831] = 12'h  0;
rom[123832] = 12'h  0;
rom[123833] = 12'h111;
rom[123834] = 12'h111;
rom[123835] = 12'h  0;
rom[123836] = 12'h  0;
rom[123837] = 12'h  0;
rom[123838] = 12'h  0;
rom[123839] = 12'h  0;
rom[123840] = 12'h  0;
rom[123841] = 12'h  0;
rom[123842] = 12'h  0;
rom[123843] = 12'h  0;
rom[123844] = 12'h  0;
rom[123845] = 12'h  0;
rom[123846] = 12'h  0;
rom[123847] = 12'h  0;
rom[123848] = 12'h  0;
rom[123849] = 12'h  0;
rom[123850] = 12'h  0;
rom[123851] = 12'h  0;
rom[123852] = 12'h  0;
rom[123853] = 12'h  0;
rom[123854] = 12'h  0;
rom[123855] = 12'h  0;
rom[123856] = 12'h  0;
rom[123857] = 12'h  0;
rom[123858] = 12'h  0;
rom[123859] = 12'h  0;
rom[123860] = 12'h  0;
rom[123861] = 12'h111;
rom[123862] = 12'h666;
rom[123863] = 12'hccc;
rom[123864] = 12'hddd;
rom[123865] = 12'h888;
rom[123866] = 12'h333;
rom[123867] = 12'h111;
rom[123868] = 12'h111;
rom[123869] = 12'h111;
rom[123870] = 12'h  0;
rom[123871] = 12'h  0;
rom[123872] = 12'h  0;
rom[123873] = 12'h  0;
rom[123874] = 12'h  0;
rom[123875] = 12'h  0;
rom[123876] = 12'h  0;
rom[123877] = 12'h111;
rom[123878] = 12'h333;
rom[123879] = 12'h777;
rom[123880] = 12'haaa;
rom[123881] = 12'h777;
rom[123882] = 12'h333;
rom[123883] = 12'h  0;
rom[123884] = 12'h  0;
rom[123885] = 12'h  0;
rom[123886] = 12'h  0;
rom[123887] = 12'h  0;
rom[123888] = 12'h  0;
rom[123889] = 12'h  0;
rom[123890] = 12'h  0;
rom[123891] = 12'h  0;
rom[123892] = 12'h  0;
rom[123893] = 12'h222;
rom[123894] = 12'h222;
rom[123895] = 12'h111;
rom[123896] = 12'h  0;
rom[123897] = 12'h  0;
rom[123898] = 12'h  0;
rom[123899] = 12'h  0;
rom[123900] = 12'h  0;
rom[123901] = 12'h  0;
rom[123902] = 12'h  0;
rom[123903] = 12'h  0;
rom[123904] = 12'h222;
rom[123905] = 12'h111;
rom[123906] = 12'h111;
rom[123907] = 12'h  0;
rom[123908] = 12'h  0;
rom[123909] = 12'h  0;
rom[123910] = 12'h  0;
rom[123911] = 12'h  0;
rom[123912] = 12'h  0;
rom[123913] = 12'h  0;
rom[123914] = 12'h  0;
rom[123915] = 12'h  0;
rom[123916] = 12'h  0;
rom[123917] = 12'h  0;
rom[123918] = 12'h  0;
rom[123919] = 12'h  0;
rom[123920] = 12'h333;
rom[123921] = 12'h444;
rom[123922] = 12'h555;
rom[123923] = 12'h444;
rom[123924] = 12'h222;
rom[123925] = 12'h111;
rom[123926] = 12'h  0;
rom[123927] = 12'h  0;
rom[123928] = 12'h  0;
rom[123929] = 12'h  0;
rom[123930] = 12'h  0;
rom[123931] = 12'h  0;
rom[123932] = 12'h  0;
rom[123933] = 12'h  0;
rom[123934] = 12'h  0;
rom[123935] = 12'h  0;
rom[123936] = 12'h  0;
rom[123937] = 12'h  0;
rom[123938] = 12'h  0;
rom[123939] = 12'h  0;
rom[123940] = 12'h  0;
rom[123941] = 12'h  0;
rom[123942] = 12'h  0;
rom[123943] = 12'h  0;
rom[123944] = 12'h  0;
rom[123945] = 12'h  0;
rom[123946] = 12'h  0;
rom[123947] = 12'h  0;
rom[123948] = 12'h  0;
rom[123949] = 12'h  0;
rom[123950] = 12'h  0;
rom[123951] = 12'h  0;
rom[123952] = 12'h  0;
rom[123953] = 12'h  0;
rom[123954] = 12'h  0;
rom[123955] = 12'h  0;
rom[123956] = 12'h  0;
rom[123957] = 12'h  0;
rom[123958] = 12'h  0;
rom[123959] = 12'h  0;
rom[123960] = 12'h  0;
rom[123961] = 12'h  0;
rom[123962] = 12'h  0;
rom[123963] = 12'h  0;
rom[123964] = 12'h  0;
rom[123965] = 12'h  0;
rom[123966] = 12'h  0;
rom[123967] = 12'h  0;
rom[123968] = 12'h  0;
rom[123969] = 12'h  0;
rom[123970] = 12'h  0;
rom[123971] = 12'h  0;
rom[123972] = 12'h  0;
rom[123973] = 12'h  0;
rom[123974] = 12'h  0;
rom[123975] = 12'h  0;
rom[123976] = 12'h  0;
rom[123977] = 12'h111;
rom[123978] = 12'h333;
rom[123979] = 12'h555;
rom[123980] = 12'h666;
rom[123981] = 12'h555;
rom[123982] = 12'h333;
rom[123983] = 12'h111;
rom[123984] = 12'h  0;
rom[123985] = 12'h  0;
rom[123986] = 12'h  0;
rom[123987] = 12'h  0;
rom[123988] = 12'h  0;
rom[123989] = 12'h  0;
rom[123990] = 12'h  0;
rom[123991] = 12'h  0;
rom[123992] = 12'h  0;
rom[123993] = 12'h  0;
rom[123994] = 12'h  0;
rom[123995] = 12'h  0;
rom[123996] = 12'h  0;
rom[123997] = 12'h  0;
rom[123998] = 12'h  0;
rom[123999] = 12'h  0;
rom[124000] = 12'hddd;
rom[124001] = 12'hddd;
rom[124002] = 12'hddd;
rom[124003] = 12'hddd;
rom[124004] = 12'hddd;
rom[124005] = 12'hddd;
rom[124006] = 12'hddd;
rom[124007] = 12'hddd;
rom[124008] = 12'hddd;
rom[124009] = 12'hccc;
rom[124010] = 12'hccc;
rom[124011] = 12'hccc;
rom[124012] = 12'hccc;
rom[124013] = 12'hccc;
rom[124014] = 12'hccc;
rom[124015] = 12'hccc;
rom[124016] = 12'hccc;
rom[124017] = 12'hccc;
rom[124018] = 12'hccc;
rom[124019] = 12'hbbb;
rom[124020] = 12'hbbb;
rom[124021] = 12'hbbb;
rom[124022] = 12'hbbb;
rom[124023] = 12'hbbb;
rom[124024] = 12'hbbb;
rom[124025] = 12'haaa;
rom[124026] = 12'haaa;
rom[124027] = 12'haaa;
rom[124028] = 12'haaa;
rom[124029] = 12'haaa;
rom[124030] = 12'haaa;
rom[124031] = 12'haaa;
rom[124032] = 12'h999;
rom[124033] = 12'h999;
rom[124034] = 12'haaa;
rom[124035] = 12'haaa;
rom[124036] = 12'h999;
rom[124037] = 12'h999;
rom[124038] = 12'h999;
rom[124039] = 12'h999;
rom[124040] = 12'h888;
rom[124041] = 12'h888;
rom[124042] = 12'h888;
rom[124043] = 12'h888;
rom[124044] = 12'h888;
rom[124045] = 12'h777;
rom[124046] = 12'h777;
rom[124047] = 12'h777;
rom[124048] = 12'h777;
rom[124049] = 12'h777;
rom[124050] = 12'h777;
rom[124051] = 12'h777;
rom[124052] = 12'h777;
rom[124053] = 12'h777;
rom[124054] = 12'h777;
rom[124055] = 12'h777;
rom[124056] = 12'h777;
rom[124057] = 12'h777;
rom[124058] = 12'h888;
rom[124059] = 12'h888;
rom[124060] = 12'h888;
rom[124061] = 12'h888;
rom[124062] = 12'h999;
rom[124063] = 12'haaa;
rom[124064] = 12'hddd;
rom[124065] = 12'hfff;
rom[124066] = 12'hfff;
rom[124067] = 12'hddd;
rom[124068] = 12'haaa;
rom[124069] = 12'h888;
rom[124070] = 12'h777;
rom[124071] = 12'h666;
rom[124072] = 12'h555;
rom[124073] = 12'h666;
rom[124074] = 12'h666;
rom[124075] = 12'h555;
rom[124076] = 12'h555;
rom[124077] = 12'h666;
rom[124078] = 12'h555;
rom[124079] = 12'h555;
rom[124080] = 12'h555;
rom[124081] = 12'h666;
rom[124082] = 12'h666;
rom[124083] = 12'h666;
rom[124084] = 12'h777;
rom[124085] = 12'h999;
rom[124086] = 12'h999;
rom[124087] = 12'h888;
rom[124088] = 12'h666;
rom[124089] = 12'h555;
rom[124090] = 12'h555;
rom[124091] = 12'h555;
rom[124092] = 12'h444;
rom[124093] = 12'h444;
rom[124094] = 12'h444;
rom[124095] = 12'h555;
rom[124096] = 12'h444;
rom[124097] = 12'h555;
rom[124098] = 12'h555;
rom[124099] = 12'h555;
rom[124100] = 12'h555;
rom[124101] = 12'h444;
rom[124102] = 12'h444;
rom[124103] = 12'h444;
rom[124104] = 12'h555;
rom[124105] = 12'h555;
rom[124106] = 12'h555;
rom[124107] = 12'h666;
rom[124108] = 12'h666;
rom[124109] = 12'h666;
rom[124110] = 12'h555;
rom[124111] = 12'h555;
rom[124112] = 12'h555;
rom[124113] = 12'h555;
rom[124114] = 12'h444;
rom[124115] = 12'h444;
rom[124116] = 12'h444;
rom[124117] = 12'h555;
rom[124118] = 12'h555;
rom[124119] = 12'h444;
rom[124120] = 12'h444;
rom[124121] = 12'h444;
rom[124122] = 12'h444;
rom[124123] = 12'h444;
rom[124124] = 12'h444;
rom[124125] = 12'h444;
rom[124126] = 12'h444;
rom[124127] = 12'h444;
rom[124128] = 12'h444;
rom[124129] = 12'h444;
rom[124130] = 12'h444;
rom[124131] = 12'h444;
rom[124132] = 12'h555;
rom[124133] = 12'h444;
rom[124134] = 12'h444;
rom[124135] = 12'h333;
rom[124136] = 12'h333;
rom[124137] = 12'h333;
rom[124138] = 12'h333;
rom[124139] = 12'h333;
rom[124140] = 12'h333;
rom[124141] = 12'h333;
rom[124142] = 12'h222;
rom[124143] = 12'h222;
rom[124144] = 12'h222;
rom[124145] = 12'h222;
rom[124146] = 12'h333;
rom[124147] = 12'h333;
rom[124148] = 12'h333;
rom[124149] = 12'h333;
rom[124150] = 12'h333;
rom[124151] = 12'h333;
rom[124152] = 12'h222;
rom[124153] = 12'h222;
rom[124154] = 12'h222;
rom[124155] = 12'h222;
rom[124156] = 12'h222;
rom[124157] = 12'h222;
rom[124158] = 12'h222;
rom[124159] = 12'h222;
rom[124160] = 12'h222;
rom[124161] = 12'h222;
rom[124162] = 12'h222;
rom[124163] = 12'h111;
rom[124164] = 12'h111;
rom[124165] = 12'h111;
rom[124166] = 12'h111;
rom[124167] = 12'h111;
rom[124168] = 12'h111;
rom[124169] = 12'h111;
rom[124170] = 12'h111;
rom[124171] = 12'h111;
rom[124172] = 12'h111;
rom[124173] = 12'h111;
rom[124174] = 12'h111;
rom[124175] = 12'h  0;
rom[124176] = 12'h  0;
rom[124177] = 12'h  0;
rom[124178] = 12'h  0;
rom[124179] = 12'h  0;
rom[124180] = 12'h  0;
rom[124181] = 12'h111;
rom[124182] = 12'h111;
rom[124183] = 12'h111;
rom[124184] = 12'h111;
rom[124185] = 12'h111;
rom[124186] = 12'h111;
rom[124187] = 12'h111;
rom[124188] = 12'h111;
rom[124189] = 12'h111;
rom[124190] = 12'h111;
rom[124191] = 12'h111;
rom[124192] = 12'h111;
rom[124193] = 12'h  0;
rom[124194] = 12'h  0;
rom[124195] = 12'h111;
rom[124196] = 12'h111;
rom[124197] = 12'h111;
rom[124198] = 12'h111;
rom[124199] = 12'h  0;
rom[124200] = 12'h  0;
rom[124201] = 12'h  0;
rom[124202] = 12'h  0;
rom[124203] = 12'h  0;
rom[124204] = 12'h  0;
rom[124205] = 12'h  0;
rom[124206] = 12'h  0;
rom[124207] = 12'h  0;
rom[124208] = 12'h  0;
rom[124209] = 12'h  0;
rom[124210] = 12'h  0;
rom[124211] = 12'h  0;
rom[124212] = 12'h  0;
rom[124213] = 12'h  0;
rom[124214] = 12'h  0;
rom[124215] = 12'h  0;
rom[124216] = 12'h  0;
rom[124217] = 12'h  0;
rom[124218] = 12'h  0;
rom[124219] = 12'h  0;
rom[124220] = 12'h  0;
rom[124221] = 12'h  0;
rom[124222] = 12'h  0;
rom[124223] = 12'h  0;
rom[124224] = 12'h  0;
rom[124225] = 12'h  0;
rom[124226] = 12'h  0;
rom[124227] = 12'h  0;
rom[124228] = 12'h  0;
rom[124229] = 12'h  0;
rom[124230] = 12'h  0;
rom[124231] = 12'h  0;
rom[124232] = 12'h  0;
rom[124233] = 12'h111;
rom[124234] = 12'h111;
rom[124235] = 12'h  0;
rom[124236] = 12'h  0;
rom[124237] = 12'h  0;
rom[124238] = 12'h  0;
rom[124239] = 12'h  0;
rom[124240] = 12'h  0;
rom[124241] = 12'h  0;
rom[124242] = 12'h  0;
rom[124243] = 12'h  0;
rom[124244] = 12'h  0;
rom[124245] = 12'h  0;
rom[124246] = 12'h  0;
rom[124247] = 12'h  0;
rom[124248] = 12'h  0;
rom[124249] = 12'h  0;
rom[124250] = 12'h  0;
rom[124251] = 12'h  0;
rom[124252] = 12'h  0;
rom[124253] = 12'h  0;
rom[124254] = 12'h  0;
rom[124255] = 12'h  0;
rom[124256] = 12'h  0;
rom[124257] = 12'h  0;
rom[124258] = 12'h  0;
rom[124259] = 12'h  0;
rom[124260] = 12'h  0;
rom[124261] = 12'h222;
rom[124262] = 12'h777;
rom[124263] = 12'hccc;
rom[124264] = 12'hccc;
rom[124265] = 12'h777;
rom[124266] = 12'h333;
rom[124267] = 12'h111;
rom[124268] = 12'h  0;
rom[124269] = 12'h  0;
rom[124270] = 12'h  0;
rom[124271] = 12'h  0;
rom[124272] = 12'h  0;
rom[124273] = 12'h  0;
rom[124274] = 12'h  0;
rom[124275] = 12'h  0;
rom[124276] = 12'h  0;
rom[124277] = 12'h  0;
rom[124278] = 12'h222;
rom[124279] = 12'h666;
rom[124280] = 12'haaa;
rom[124281] = 12'h777;
rom[124282] = 12'h333;
rom[124283] = 12'h  0;
rom[124284] = 12'h  0;
rom[124285] = 12'h  0;
rom[124286] = 12'h  0;
rom[124287] = 12'h  0;
rom[124288] = 12'h  0;
rom[124289] = 12'h  0;
rom[124290] = 12'h  0;
rom[124291] = 12'h  0;
rom[124292] = 12'h  0;
rom[124293] = 12'h111;
rom[124294] = 12'h222;
rom[124295] = 12'h111;
rom[124296] = 12'h  0;
rom[124297] = 12'h  0;
rom[124298] = 12'h  0;
rom[124299] = 12'h  0;
rom[124300] = 12'h  0;
rom[124301] = 12'h  0;
rom[124302] = 12'h  0;
rom[124303] = 12'h  0;
rom[124304] = 12'h111;
rom[124305] = 12'h111;
rom[124306] = 12'h111;
rom[124307] = 12'h  0;
rom[124308] = 12'h  0;
rom[124309] = 12'h  0;
rom[124310] = 12'h  0;
rom[124311] = 12'h  0;
rom[124312] = 12'h  0;
rom[124313] = 12'h  0;
rom[124314] = 12'h  0;
rom[124315] = 12'h  0;
rom[124316] = 12'h  0;
rom[124317] = 12'h  0;
rom[124318] = 12'h  0;
rom[124319] = 12'h  0;
rom[124320] = 12'h222;
rom[124321] = 12'h444;
rom[124322] = 12'h444;
rom[124323] = 12'h333;
rom[124324] = 12'h222;
rom[124325] = 12'h111;
rom[124326] = 12'h  0;
rom[124327] = 12'h  0;
rom[124328] = 12'h  0;
rom[124329] = 12'h  0;
rom[124330] = 12'h  0;
rom[124331] = 12'h  0;
rom[124332] = 12'h  0;
rom[124333] = 12'h  0;
rom[124334] = 12'h  0;
rom[124335] = 12'h  0;
rom[124336] = 12'h  0;
rom[124337] = 12'h  0;
rom[124338] = 12'h  0;
rom[124339] = 12'h  0;
rom[124340] = 12'h  0;
rom[124341] = 12'h  0;
rom[124342] = 12'h  0;
rom[124343] = 12'h  0;
rom[124344] = 12'h  0;
rom[124345] = 12'h  0;
rom[124346] = 12'h  0;
rom[124347] = 12'h  0;
rom[124348] = 12'h  0;
rom[124349] = 12'h  0;
rom[124350] = 12'h  0;
rom[124351] = 12'h  0;
rom[124352] = 12'h  0;
rom[124353] = 12'h  0;
rom[124354] = 12'h  0;
rom[124355] = 12'h  0;
rom[124356] = 12'h  0;
rom[124357] = 12'h  0;
rom[124358] = 12'h  0;
rom[124359] = 12'h  0;
rom[124360] = 12'h  0;
rom[124361] = 12'h  0;
rom[124362] = 12'h  0;
rom[124363] = 12'h  0;
rom[124364] = 12'h  0;
rom[124365] = 12'h  0;
rom[124366] = 12'h  0;
rom[124367] = 12'h  0;
rom[124368] = 12'h  0;
rom[124369] = 12'h  0;
rom[124370] = 12'h  0;
rom[124371] = 12'h  0;
rom[124372] = 12'h  0;
rom[124373] = 12'h  0;
rom[124374] = 12'h  0;
rom[124375] = 12'h  0;
rom[124376] = 12'h  0;
rom[124377] = 12'h111;
rom[124378] = 12'h222;
rom[124379] = 12'h444;
rom[124380] = 12'h555;
rom[124381] = 12'h555;
rom[124382] = 12'h333;
rom[124383] = 12'h111;
rom[124384] = 12'h  0;
rom[124385] = 12'h  0;
rom[124386] = 12'h  0;
rom[124387] = 12'h  0;
rom[124388] = 12'h  0;
rom[124389] = 12'h  0;
rom[124390] = 12'h  0;
rom[124391] = 12'h  0;
rom[124392] = 12'h  0;
rom[124393] = 12'h  0;
rom[124394] = 12'h  0;
rom[124395] = 12'h  0;
rom[124396] = 12'h  0;
rom[124397] = 12'h  0;
rom[124398] = 12'h  0;
rom[124399] = 12'h  0;
rom[124400] = 12'hddd;
rom[124401] = 12'hddd;
rom[124402] = 12'hddd;
rom[124403] = 12'hddd;
rom[124404] = 12'hddd;
rom[124405] = 12'hccc;
rom[124406] = 12'hccc;
rom[124407] = 12'hccc;
rom[124408] = 12'hccc;
rom[124409] = 12'hccc;
rom[124410] = 12'hccc;
rom[124411] = 12'hccc;
rom[124412] = 12'hccc;
rom[124413] = 12'hbbb;
rom[124414] = 12'hbbb;
rom[124415] = 12'hbbb;
rom[124416] = 12'hbbb;
rom[124417] = 12'hbbb;
rom[124418] = 12'hbbb;
rom[124419] = 12'hbbb;
rom[124420] = 12'hbbb;
rom[124421] = 12'hbbb;
rom[124422] = 12'hbbb;
rom[124423] = 12'hbbb;
rom[124424] = 12'haaa;
rom[124425] = 12'haaa;
rom[124426] = 12'haaa;
rom[124427] = 12'haaa;
rom[124428] = 12'haaa;
rom[124429] = 12'haaa;
rom[124430] = 12'h999;
rom[124431] = 12'h999;
rom[124432] = 12'h999;
rom[124433] = 12'h999;
rom[124434] = 12'h999;
rom[124435] = 12'h999;
rom[124436] = 12'h999;
rom[124437] = 12'h999;
rom[124438] = 12'h999;
rom[124439] = 12'h888;
rom[124440] = 12'h888;
rom[124441] = 12'h888;
rom[124442] = 12'h888;
rom[124443] = 12'h888;
rom[124444] = 12'h888;
rom[124445] = 12'h777;
rom[124446] = 12'h777;
rom[124447] = 12'h777;
rom[124448] = 12'h777;
rom[124449] = 12'h777;
rom[124450] = 12'h777;
rom[124451] = 12'h777;
rom[124452] = 12'h777;
rom[124453] = 12'h777;
rom[124454] = 12'h777;
rom[124455] = 12'h777;
rom[124456] = 12'h777;
rom[124457] = 12'h777;
rom[124458] = 12'h777;
rom[124459] = 12'h888;
rom[124460] = 12'h888;
rom[124461] = 12'h888;
rom[124462] = 12'h999;
rom[124463] = 12'haaa;
rom[124464] = 12'heee;
rom[124465] = 12'hfff;
rom[124466] = 12'hfff;
rom[124467] = 12'hccc;
rom[124468] = 12'h999;
rom[124469] = 12'h888;
rom[124470] = 12'h777;
rom[124471] = 12'h666;
rom[124472] = 12'h555;
rom[124473] = 12'h666;
rom[124474] = 12'h666;
rom[124475] = 12'h555;
rom[124476] = 12'h555;
rom[124477] = 12'h666;
rom[124478] = 12'h555;
rom[124479] = 12'h555;
rom[124480] = 12'h555;
rom[124481] = 12'h555;
rom[124482] = 12'h666;
rom[124483] = 12'h666;
rom[124484] = 12'h888;
rom[124485] = 12'h999;
rom[124486] = 12'h888;
rom[124487] = 12'h666;
rom[124488] = 12'h555;
rom[124489] = 12'h555;
rom[124490] = 12'h555;
rom[124491] = 12'h555;
rom[124492] = 12'h444;
rom[124493] = 12'h444;
rom[124494] = 12'h444;
rom[124495] = 12'h444;
rom[124496] = 12'h444;
rom[124497] = 12'h555;
rom[124498] = 12'h555;
rom[124499] = 12'h555;
rom[124500] = 12'h555;
rom[124501] = 12'h444;
rom[124502] = 12'h444;
rom[124503] = 12'h444;
rom[124504] = 12'h555;
rom[124505] = 12'h444;
rom[124506] = 12'h555;
rom[124507] = 12'h555;
rom[124508] = 12'h666;
rom[124509] = 12'h555;
rom[124510] = 12'h555;
rom[124511] = 12'h555;
rom[124512] = 12'h555;
rom[124513] = 12'h555;
rom[124514] = 12'h555;
rom[124515] = 12'h444;
rom[124516] = 12'h444;
rom[124517] = 12'h555;
rom[124518] = 12'h555;
rom[124519] = 12'h444;
rom[124520] = 12'h444;
rom[124521] = 12'h444;
rom[124522] = 12'h444;
rom[124523] = 12'h444;
rom[124524] = 12'h444;
rom[124525] = 12'h444;
rom[124526] = 12'h333;
rom[124527] = 12'h333;
rom[124528] = 12'h444;
rom[124529] = 12'h444;
rom[124530] = 12'h444;
rom[124531] = 12'h444;
rom[124532] = 12'h555;
rom[124533] = 12'h555;
rom[124534] = 12'h444;
rom[124535] = 12'h333;
rom[124536] = 12'h333;
rom[124537] = 12'h333;
rom[124538] = 12'h333;
rom[124539] = 12'h333;
rom[124540] = 12'h333;
rom[124541] = 12'h333;
rom[124542] = 12'h222;
rom[124543] = 12'h222;
rom[124544] = 12'h222;
rom[124545] = 12'h222;
rom[124546] = 12'h333;
rom[124547] = 12'h333;
rom[124548] = 12'h333;
rom[124549] = 12'h333;
rom[124550] = 12'h333;
rom[124551] = 12'h222;
rom[124552] = 12'h222;
rom[124553] = 12'h222;
rom[124554] = 12'h222;
rom[124555] = 12'h222;
rom[124556] = 12'h222;
rom[124557] = 12'h222;
rom[124558] = 12'h222;
rom[124559] = 12'h222;
rom[124560] = 12'h222;
rom[124561] = 12'h222;
rom[124562] = 12'h222;
rom[124563] = 12'h111;
rom[124564] = 12'h111;
rom[124565] = 12'h111;
rom[124566] = 12'h111;
rom[124567] = 12'h111;
rom[124568] = 12'h111;
rom[124569] = 12'h111;
rom[124570] = 12'h  0;
rom[124571] = 12'h111;
rom[124572] = 12'h111;
rom[124573] = 12'h111;
rom[124574] = 12'h111;
rom[124575] = 12'h111;
rom[124576] = 12'h111;
rom[124577] = 12'h  0;
rom[124578] = 12'h  0;
rom[124579] = 12'h  0;
rom[124580] = 12'h  0;
rom[124581] = 12'h111;
rom[124582] = 12'h111;
rom[124583] = 12'h111;
rom[124584] = 12'h111;
rom[124585] = 12'h111;
rom[124586] = 12'h111;
rom[124587] = 12'h111;
rom[124588] = 12'h111;
rom[124589] = 12'h111;
rom[124590] = 12'h111;
rom[124591] = 12'h111;
rom[124592] = 12'h  0;
rom[124593] = 12'h  0;
rom[124594] = 12'h  0;
rom[124595] = 12'h  0;
rom[124596] = 12'h111;
rom[124597] = 12'h111;
rom[124598] = 12'h111;
rom[124599] = 12'h  0;
rom[124600] = 12'h  0;
rom[124601] = 12'h  0;
rom[124602] = 12'h  0;
rom[124603] = 12'h  0;
rom[124604] = 12'h  0;
rom[124605] = 12'h  0;
rom[124606] = 12'h  0;
rom[124607] = 12'h  0;
rom[124608] = 12'h  0;
rom[124609] = 12'h  0;
rom[124610] = 12'h  0;
rom[124611] = 12'h  0;
rom[124612] = 12'h  0;
rom[124613] = 12'h  0;
rom[124614] = 12'h  0;
rom[124615] = 12'h  0;
rom[124616] = 12'h  0;
rom[124617] = 12'h  0;
rom[124618] = 12'h  0;
rom[124619] = 12'h  0;
rom[124620] = 12'h  0;
rom[124621] = 12'h  0;
rom[124622] = 12'h  0;
rom[124623] = 12'h  0;
rom[124624] = 12'h  0;
rom[124625] = 12'h  0;
rom[124626] = 12'h  0;
rom[124627] = 12'h  0;
rom[124628] = 12'h  0;
rom[124629] = 12'h  0;
rom[124630] = 12'h  0;
rom[124631] = 12'h  0;
rom[124632] = 12'h111;
rom[124633] = 12'h111;
rom[124634] = 12'h  0;
rom[124635] = 12'h  0;
rom[124636] = 12'h  0;
rom[124637] = 12'h  0;
rom[124638] = 12'h  0;
rom[124639] = 12'h  0;
rom[124640] = 12'h  0;
rom[124641] = 12'h  0;
rom[124642] = 12'h  0;
rom[124643] = 12'h  0;
rom[124644] = 12'h  0;
rom[124645] = 12'h  0;
rom[124646] = 12'h  0;
rom[124647] = 12'h  0;
rom[124648] = 12'h  0;
rom[124649] = 12'h  0;
rom[124650] = 12'h  0;
rom[124651] = 12'h  0;
rom[124652] = 12'h  0;
rom[124653] = 12'h  0;
rom[124654] = 12'h  0;
rom[124655] = 12'h  0;
rom[124656] = 12'h  0;
rom[124657] = 12'h  0;
rom[124658] = 12'h  0;
rom[124659] = 12'h  0;
rom[124660] = 12'h  0;
rom[124661] = 12'h222;
rom[124662] = 12'h777;
rom[124663] = 12'hccc;
rom[124664] = 12'hccc;
rom[124665] = 12'h777;
rom[124666] = 12'h222;
rom[124667] = 12'h111;
rom[124668] = 12'h  0;
rom[124669] = 12'h  0;
rom[124670] = 12'h  0;
rom[124671] = 12'h  0;
rom[124672] = 12'h  0;
rom[124673] = 12'h  0;
rom[124674] = 12'h  0;
rom[124675] = 12'h  0;
rom[124676] = 12'h  0;
rom[124677] = 12'h  0;
rom[124678] = 12'h222;
rom[124679] = 12'h555;
rom[124680] = 12'haaa;
rom[124681] = 12'h777;
rom[124682] = 12'h333;
rom[124683] = 12'h  0;
rom[124684] = 12'h111;
rom[124685] = 12'h  0;
rom[124686] = 12'h  0;
rom[124687] = 12'h  0;
rom[124688] = 12'h  0;
rom[124689] = 12'h  0;
rom[124690] = 12'h  0;
rom[124691] = 12'h  0;
rom[124692] = 12'h  0;
rom[124693] = 12'h111;
rom[124694] = 12'h222;
rom[124695] = 12'h111;
rom[124696] = 12'h  0;
rom[124697] = 12'h  0;
rom[124698] = 12'h  0;
rom[124699] = 12'h  0;
rom[124700] = 12'h  0;
rom[124701] = 12'h  0;
rom[124702] = 12'h  0;
rom[124703] = 12'h  0;
rom[124704] = 12'h  0;
rom[124705] = 12'h111;
rom[124706] = 12'h111;
rom[124707] = 12'h  0;
rom[124708] = 12'h  0;
rom[124709] = 12'h  0;
rom[124710] = 12'h  0;
rom[124711] = 12'h  0;
rom[124712] = 12'h  0;
rom[124713] = 12'h  0;
rom[124714] = 12'h  0;
rom[124715] = 12'h  0;
rom[124716] = 12'h  0;
rom[124717] = 12'h  0;
rom[124718] = 12'h  0;
rom[124719] = 12'h  0;
rom[124720] = 12'h222;
rom[124721] = 12'h333;
rom[124722] = 12'h444;
rom[124723] = 12'h333;
rom[124724] = 12'h222;
rom[124725] = 12'h111;
rom[124726] = 12'h  0;
rom[124727] = 12'h  0;
rom[124728] = 12'h  0;
rom[124729] = 12'h  0;
rom[124730] = 12'h  0;
rom[124731] = 12'h  0;
rom[124732] = 12'h  0;
rom[124733] = 12'h  0;
rom[124734] = 12'h  0;
rom[124735] = 12'h  0;
rom[124736] = 12'h  0;
rom[124737] = 12'h  0;
rom[124738] = 12'h  0;
rom[124739] = 12'h  0;
rom[124740] = 12'h  0;
rom[124741] = 12'h  0;
rom[124742] = 12'h  0;
rom[124743] = 12'h  0;
rom[124744] = 12'h  0;
rom[124745] = 12'h  0;
rom[124746] = 12'h  0;
rom[124747] = 12'h  0;
rom[124748] = 12'h  0;
rom[124749] = 12'h  0;
rom[124750] = 12'h  0;
rom[124751] = 12'h  0;
rom[124752] = 12'h  0;
rom[124753] = 12'h  0;
rom[124754] = 12'h  0;
rom[124755] = 12'h  0;
rom[124756] = 12'h  0;
rom[124757] = 12'h  0;
rom[124758] = 12'h  0;
rom[124759] = 12'h  0;
rom[124760] = 12'h  0;
rom[124761] = 12'h  0;
rom[124762] = 12'h  0;
rom[124763] = 12'h  0;
rom[124764] = 12'h  0;
rom[124765] = 12'h  0;
rom[124766] = 12'h  0;
rom[124767] = 12'h  0;
rom[124768] = 12'h  0;
rom[124769] = 12'h  0;
rom[124770] = 12'h  0;
rom[124771] = 12'h  0;
rom[124772] = 12'h  0;
rom[124773] = 12'h  0;
rom[124774] = 12'h  0;
rom[124775] = 12'h  0;
rom[124776] = 12'h  0;
rom[124777] = 12'h  0;
rom[124778] = 12'h222;
rom[124779] = 12'h444;
rom[124780] = 12'h555;
rom[124781] = 12'h555;
rom[124782] = 12'h333;
rom[124783] = 12'h111;
rom[124784] = 12'h  0;
rom[124785] = 12'h  0;
rom[124786] = 12'h  0;
rom[124787] = 12'h  0;
rom[124788] = 12'h  0;
rom[124789] = 12'h  0;
rom[124790] = 12'h  0;
rom[124791] = 12'h  0;
rom[124792] = 12'h  0;
rom[124793] = 12'h  0;
rom[124794] = 12'h  0;
rom[124795] = 12'h  0;
rom[124796] = 12'h  0;
rom[124797] = 12'h  0;
rom[124798] = 12'h  0;
rom[124799] = 12'h  0;
rom[124800] = 12'hddd;
rom[124801] = 12'hddd;
rom[124802] = 12'hddd;
rom[124803] = 12'hccc;
rom[124804] = 12'hccc;
rom[124805] = 12'hccc;
rom[124806] = 12'hccc;
rom[124807] = 12'hccc;
rom[124808] = 12'hccc;
rom[124809] = 12'hccc;
rom[124810] = 12'hccc;
rom[124811] = 12'hbbb;
rom[124812] = 12'hbbb;
rom[124813] = 12'hbbb;
rom[124814] = 12'hbbb;
rom[124815] = 12'hbbb;
rom[124816] = 12'hbbb;
rom[124817] = 12'hbbb;
rom[124818] = 12'hbbb;
rom[124819] = 12'hbbb;
rom[124820] = 12'hbbb;
rom[124821] = 12'haaa;
rom[124822] = 12'haaa;
rom[124823] = 12'haaa;
rom[124824] = 12'haaa;
rom[124825] = 12'haaa;
rom[124826] = 12'haaa;
rom[124827] = 12'h999;
rom[124828] = 12'h999;
rom[124829] = 12'h999;
rom[124830] = 12'h999;
rom[124831] = 12'h999;
rom[124832] = 12'h999;
rom[124833] = 12'h999;
rom[124834] = 12'h999;
rom[124835] = 12'h999;
rom[124836] = 12'h999;
rom[124837] = 12'h999;
rom[124838] = 12'h888;
rom[124839] = 12'h888;
rom[124840] = 12'h888;
rom[124841] = 12'h888;
rom[124842] = 12'h888;
rom[124843] = 12'h888;
rom[124844] = 12'h777;
rom[124845] = 12'h777;
rom[124846] = 12'h777;
rom[124847] = 12'h777;
rom[124848] = 12'h777;
rom[124849] = 12'h777;
rom[124850] = 12'h777;
rom[124851] = 12'h777;
rom[124852] = 12'h777;
rom[124853] = 12'h777;
rom[124854] = 12'h666;
rom[124855] = 12'h666;
rom[124856] = 12'h666;
rom[124857] = 12'h666;
rom[124858] = 12'h777;
rom[124859] = 12'h888;
rom[124860] = 12'h888;
rom[124861] = 12'h888;
rom[124862] = 12'haaa;
rom[124863] = 12'hccc;
rom[124864] = 12'hfff;
rom[124865] = 12'heee;
rom[124866] = 12'hddd;
rom[124867] = 12'haaa;
rom[124868] = 12'h888;
rom[124869] = 12'h777;
rom[124870] = 12'h666;
rom[124871] = 12'h666;
rom[124872] = 12'h555;
rom[124873] = 12'h555;
rom[124874] = 12'h555;
rom[124875] = 12'h555;
rom[124876] = 12'h555;
rom[124877] = 12'h555;
rom[124878] = 12'h555;
rom[124879] = 12'h555;
rom[124880] = 12'h444;
rom[124881] = 12'h555;
rom[124882] = 12'h666;
rom[124883] = 12'h888;
rom[124884] = 12'h999;
rom[124885] = 12'h888;
rom[124886] = 12'h777;
rom[124887] = 12'h666;
rom[124888] = 12'h555;
rom[124889] = 12'h555;
rom[124890] = 12'h555;
rom[124891] = 12'h555;
rom[124892] = 12'h444;
rom[124893] = 12'h444;
rom[124894] = 12'h444;
rom[124895] = 12'h444;
rom[124896] = 12'h444;
rom[124897] = 12'h444;
rom[124898] = 12'h555;
rom[124899] = 12'h555;
rom[124900] = 12'h444;
rom[124901] = 12'h444;
rom[124902] = 12'h444;
rom[124903] = 12'h444;
rom[124904] = 12'h444;
rom[124905] = 12'h444;
rom[124906] = 12'h444;
rom[124907] = 12'h444;
rom[124908] = 12'h555;
rom[124909] = 12'h555;
rom[124910] = 12'h666;
rom[124911] = 12'h666;
rom[124912] = 12'h555;
rom[124913] = 12'h555;
rom[124914] = 12'h444;
rom[124915] = 12'h444;
rom[124916] = 12'h444;
rom[124917] = 12'h555;
rom[124918] = 12'h555;
rom[124919] = 12'h444;
rom[124920] = 12'h444;
rom[124921] = 12'h444;
rom[124922] = 12'h444;
rom[124923] = 12'h444;
rom[124924] = 12'h444;
rom[124925] = 12'h444;
rom[124926] = 12'h333;
rom[124927] = 12'h333;
rom[124928] = 12'h333;
rom[124929] = 12'h333;
rom[124930] = 12'h333;
rom[124931] = 12'h444;
rom[124932] = 12'h444;
rom[124933] = 12'h555;
rom[124934] = 12'h444;
rom[124935] = 12'h444;
rom[124936] = 12'h333;
rom[124937] = 12'h333;
rom[124938] = 12'h333;
rom[124939] = 12'h222;
rom[124940] = 12'h222;
rom[124941] = 12'h222;
rom[124942] = 12'h222;
rom[124943] = 12'h222;
rom[124944] = 12'h222;
rom[124945] = 12'h222;
rom[124946] = 12'h333;
rom[124947] = 12'h333;
rom[124948] = 12'h333;
rom[124949] = 12'h222;
rom[124950] = 12'h222;
rom[124951] = 12'h222;
rom[124952] = 12'h222;
rom[124953] = 12'h222;
rom[124954] = 12'h222;
rom[124955] = 12'h222;
rom[124956] = 12'h222;
rom[124957] = 12'h222;
rom[124958] = 12'h222;
rom[124959] = 12'h222;
rom[124960] = 12'h222;
rom[124961] = 12'h222;
rom[124962] = 12'h111;
rom[124963] = 12'h111;
rom[124964] = 12'h111;
rom[124965] = 12'h111;
rom[124966] = 12'h111;
rom[124967] = 12'h  0;
rom[124968] = 12'h  0;
rom[124969] = 12'h  0;
rom[124970] = 12'h  0;
rom[124971] = 12'h  0;
rom[124972] = 12'h111;
rom[124973] = 12'h111;
rom[124974] = 12'h  0;
rom[124975] = 12'h  0;
rom[124976] = 12'h  0;
rom[124977] = 12'h  0;
rom[124978] = 12'h  0;
rom[124979] = 12'h  0;
rom[124980] = 12'h  0;
rom[124981] = 12'h  0;
rom[124982] = 12'h111;
rom[124983] = 12'h111;
rom[124984] = 12'h111;
rom[124985] = 12'h111;
rom[124986] = 12'h111;
rom[124987] = 12'h111;
rom[124988] = 12'h111;
rom[124989] = 12'h111;
rom[124990] = 12'h111;
rom[124991] = 12'h111;
rom[124992] = 12'h  0;
rom[124993] = 12'h  0;
rom[124994] = 12'h  0;
rom[124995] = 12'h  0;
rom[124996] = 12'h  0;
rom[124997] = 12'h  0;
rom[124998] = 12'h  0;
rom[124999] = 12'h  0;
rom[125000] = 12'h  0;
rom[125001] = 12'h  0;
rom[125002] = 12'h  0;
rom[125003] = 12'h  0;
rom[125004] = 12'h  0;
rom[125005] = 12'h  0;
rom[125006] = 12'h  0;
rom[125007] = 12'h  0;
rom[125008] = 12'h  0;
rom[125009] = 12'h  0;
rom[125010] = 12'h  0;
rom[125011] = 12'h  0;
rom[125012] = 12'h  0;
rom[125013] = 12'h  0;
rom[125014] = 12'h  0;
rom[125015] = 12'h  0;
rom[125016] = 12'h  0;
rom[125017] = 12'h  0;
rom[125018] = 12'h  0;
rom[125019] = 12'h  0;
rom[125020] = 12'h  0;
rom[125021] = 12'h  0;
rom[125022] = 12'h  0;
rom[125023] = 12'h  0;
rom[125024] = 12'h  0;
rom[125025] = 12'h  0;
rom[125026] = 12'h  0;
rom[125027] = 12'h  0;
rom[125028] = 12'h  0;
rom[125029] = 12'h  0;
rom[125030] = 12'h  0;
rom[125031] = 12'h  0;
rom[125032] = 12'h  0;
rom[125033] = 12'h  0;
rom[125034] = 12'h  0;
rom[125035] = 12'h  0;
rom[125036] = 12'h  0;
rom[125037] = 12'h  0;
rom[125038] = 12'h  0;
rom[125039] = 12'h  0;
rom[125040] = 12'h  0;
rom[125041] = 12'h  0;
rom[125042] = 12'h  0;
rom[125043] = 12'h  0;
rom[125044] = 12'h  0;
rom[125045] = 12'h  0;
rom[125046] = 12'h  0;
rom[125047] = 12'h  0;
rom[125048] = 12'h  0;
rom[125049] = 12'h  0;
rom[125050] = 12'h  0;
rom[125051] = 12'h  0;
rom[125052] = 12'h  0;
rom[125053] = 12'h  0;
rom[125054] = 12'h  0;
rom[125055] = 12'h  0;
rom[125056] = 12'h  0;
rom[125057] = 12'h  0;
rom[125058] = 12'h  0;
rom[125059] = 12'h  0;
rom[125060] = 12'h111;
rom[125061] = 12'h333;
rom[125062] = 12'h777;
rom[125063] = 12'hccc;
rom[125064] = 12'hbbb;
rom[125065] = 12'h666;
rom[125066] = 12'h222;
rom[125067] = 12'h111;
rom[125068] = 12'h  0;
rom[125069] = 12'h  0;
rom[125070] = 12'h  0;
rom[125071] = 12'h  0;
rom[125072] = 12'h  0;
rom[125073] = 12'h  0;
rom[125074] = 12'h  0;
rom[125075] = 12'h  0;
rom[125076] = 12'h  0;
rom[125077] = 12'h  0;
rom[125078] = 12'h222;
rom[125079] = 12'h444;
rom[125080] = 12'h888;
rom[125081] = 12'h777;
rom[125082] = 12'h333;
rom[125083] = 12'h  0;
rom[125084] = 12'h  0;
rom[125085] = 12'h  0;
rom[125086] = 12'h  0;
rom[125087] = 12'h  0;
rom[125088] = 12'h  0;
rom[125089] = 12'h  0;
rom[125090] = 12'h  0;
rom[125091] = 12'h  0;
rom[125092] = 12'h  0;
rom[125093] = 12'h111;
rom[125094] = 12'h111;
rom[125095] = 12'h111;
rom[125096] = 12'h  0;
rom[125097] = 12'h  0;
rom[125098] = 12'h  0;
rom[125099] = 12'h  0;
rom[125100] = 12'h  0;
rom[125101] = 12'h  0;
rom[125102] = 12'h  0;
rom[125103] = 12'h  0;
rom[125104] = 12'h  0;
rom[125105] = 12'h  0;
rom[125106] = 12'h  0;
rom[125107] = 12'h  0;
rom[125108] = 12'h  0;
rom[125109] = 12'h  0;
rom[125110] = 12'h  0;
rom[125111] = 12'h  0;
rom[125112] = 12'h  0;
rom[125113] = 12'h  0;
rom[125114] = 12'h  0;
rom[125115] = 12'h  0;
rom[125116] = 12'h  0;
rom[125117] = 12'h  0;
rom[125118] = 12'h  0;
rom[125119] = 12'h  0;
rom[125120] = 12'h222;
rom[125121] = 12'h333;
rom[125122] = 12'h444;
rom[125123] = 12'h333;
rom[125124] = 12'h222;
rom[125125] = 12'h  0;
rom[125126] = 12'h  0;
rom[125127] = 12'h  0;
rom[125128] = 12'h  0;
rom[125129] = 12'h  0;
rom[125130] = 12'h  0;
rom[125131] = 12'h  0;
rom[125132] = 12'h  0;
rom[125133] = 12'h  0;
rom[125134] = 12'h  0;
rom[125135] = 12'h  0;
rom[125136] = 12'h  0;
rom[125137] = 12'h  0;
rom[125138] = 12'h  0;
rom[125139] = 12'h  0;
rom[125140] = 12'h  0;
rom[125141] = 12'h  0;
rom[125142] = 12'h  0;
rom[125143] = 12'h  0;
rom[125144] = 12'h  0;
rom[125145] = 12'h  0;
rom[125146] = 12'h  0;
rom[125147] = 12'h  0;
rom[125148] = 12'h  0;
rom[125149] = 12'h  0;
rom[125150] = 12'h  0;
rom[125151] = 12'h  0;
rom[125152] = 12'h  0;
rom[125153] = 12'h  0;
rom[125154] = 12'h  0;
rom[125155] = 12'h  0;
rom[125156] = 12'h  0;
rom[125157] = 12'h  0;
rom[125158] = 12'h  0;
rom[125159] = 12'h  0;
rom[125160] = 12'h  0;
rom[125161] = 12'h  0;
rom[125162] = 12'h  0;
rom[125163] = 12'h  0;
rom[125164] = 12'h  0;
rom[125165] = 12'h  0;
rom[125166] = 12'h  0;
rom[125167] = 12'h  0;
rom[125168] = 12'h  0;
rom[125169] = 12'h  0;
rom[125170] = 12'h  0;
rom[125171] = 12'h  0;
rom[125172] = 12'h  0;
rom[125173] = 12'h  0;
rom[125174] = 12'h  0;
rom[125175] = 12'h  0;
rom[125176] = 12'h  0;
rom[125177] = 12'h  0;
rom[125178] = 12'h111;
rom[125179] = 12'h222;
rom[125180] = 12'h444;
rom[125181] = 12'h555;
rom[125182] = 12'h444;
rom[125183] = 12'h111;
rom[125184] = 12'h111;
rom[125185] = 12'h  0;
rom[125186] = 12'h  0;
rom[125187] = 12'h  0;
rom[125188] = 12'h  0;
rom[125189] = 12'h  0;
rom[125190] = 12'h  0;
rom[125191] = 12'h  0;
rom[125192] = 12'h  0;
rom[125193] = 12'h  0;
rom[125194] = 12'h  0;
rom[125195] = 12'h  0;
rom[125196] = 12'h  0;
rom[125197] = 12'h  0;
rom[125198] = 12'h  0;
rom[125199] = 12'h  0;
rom[125200] = 12'hddd;
rom[125201] = 12'hddd;
rom[125202] = 12'hccc;
rom[125203] = 12'hccc;
rom[125204] = 12'hccc;
rom[125205] = 12'hccc;
rom[125206] = 12'hccc;
rom[125207] = 12'hccc;
rom[125208] = 12'hbbb;
rom[125209] = 12'hbbb;
rom[125210] = 12'hbbb;
rom[125211] = 12'hbbb;
rom[125212] = 12'hbbb;
rom[125213] = 12'hbbb;
rom[125214] = 12'hbbb;
rom[125215] = 12'haaa;
rom[125216] = 12'haaa;
rom[125217] = 12'haaa;
rom[125218] = 12'hbbb;
rom[125219] = 12'hbbb;
rom[125220] = 12'haaa;
rom[125221] = 12'haaa;
rom[125222] = 12'haaa;
rom[125223] = 12'haaa;
rom[125224] = 12'haaa;
rom[125225] = 12'haaa;
rom[125226] = 12'h999;
rom[125227] = 12'h999;
rom[125228] = 12'h999;
rom[125229] = 12'h999;
rom[125230] = 12'h999;
rom[125231] = 12'h999;
rom[125232] = 12'h999;
rom[125233] = 12'h999;
rom[125234] = 12'h999;
rom[125235] = 12'h999;
rom[125236] = 12'h999;
rom[125237] = 12'h888;
rom[125238] = 12'h888;
rom[125239] = 12'h888;
rom[125240] = 12'h888;
rom[125241] = 12'h888;
rom[125242] = 12'h888;
rom[125243] = 12'h888;
rom[125244] = 12'h777;
rom[125245] = 12'h777;
rom[125246] = 12'h777;
rom[125247] = 12'h777;
rom[125248] = 12'h777;
rom[125249] = 12'h777;
rom[125250] = 12'h777;
rom[125251] = 12'h777;
rom[125252] = 12'h777;
rom[125253] = 12'h777;
rom[125254] = 12'h666;
rom[125255] = 12'h666;
rom[125256] = 12'h666;
rom[125257] = 12'h666;
rom[125258] = 12'h777;
rom[125259] = 12'h777;
rom[125260] = 12'h888;
rom[125261] = 12'h999;
rom[125262] = 12'hbbb;
rom[125263] = 12'heee;
rom[125264] = 12'hfff;
rom[125265] = 12'heee;
rom[125266] = 12'hbbb;
rom[125267] = 12'h999;
rom[125268] = 12'h777;
rom[125269] = 12'h777;
rom[125270] = 12'h666;
rom[125271] = 12'h555;
rom[125272] = 12'h555;
rom[125273] = 12'h555;
rom[125274] = 12'h555;
rom[125275] = 12'h555;
rom[125276] = 12'h555;
rom[125277] = 12'h555;
rom[125278] = 12'h555;
rom[125279] = 12'h555;
rom[125280] = 12'h444;
rom[125281] = 12'h555;
rom[125282] = 12'h777;
rom[125283] = 12'h888;
rom[125284] = 12'h888;
rom[125285] = 12'h777;
rom[125286] = 12'h666;
rom[125287] = 12'h666;
rom[125288] = 12'h555;
rom[125289] = 12'h555;
rom[125290] = 12'h555;
rom[125291] = 12'h555;
rom[125292] = 12'h444;
rom[125293] = 12'h444;
rom[125294] = 12'h444;
rom[125295] = 12'h444;
rom[125296] = 12'h444;
rom[125297] = 12'h444;
rom[125298] = 12'h444;
rom[125299] = 12'h444;
rom[125300] = 12'h444;
rom[125301] = 12'h444;
rom[125302] = 12'h444;
rom[125303] = 12'h444;
rom[125304] = 12'h444;
rom[125305] = 12'h444;
rom[125306] = 12'h444;
rom[125307] = 12'h444;
rom[125308] = 12'h555;
rom[125309] = 12'h555;
rom[125310] = 12'h666;
rom[125311] = 12'h666;
rom[125312] = 12'h555;
rom[125313] = 12'h555;
rom[125314] = 12'h555;
rom[125315] = 12'h444;
rom[125316] = 12'h444;
rom[125317] = 12'h444;
rom[125318] = 12'h444;
rom[125319] = 12'h444;
rom[125320] = 12'h444;
rom[125321] = 12'h444;
rom[125322] = 12'h444;
rom[125323] = 12'h444;
rom[125324] = 12'h444;
rom[125325] = 12'h444;
rom[125326] = 12'h333;
rom[125327] = 12'h333;
rom[125328] = 12'h333;
rom[125329] = 12'h333;
rom[125330] = 12'h333;
rom[125331] = 12'h444;
rom[125332] = 12'h444;
rom[125333] = 12'h555;
rom[125334] = 12'h444;
rom[125335] = 12'h444;
rom[125336] = 12'h333;
rom[125337] = 12'h333;
rom[125338] = 12'h333;
rom[125339] = 12'h222;
rom[125340] = 12'h222;
rom[125341] = 12'h222;
rom[125342] = 12'h222;
rom[125343] = 12'h222;
rom[125344] = 12'h222;
rom[125345] = 12'h222;
rom[125346] = 12'h333;
rom[125347] = 12'h333;
rom[125348] = 12'h333;
rom[125349] = 12'h222;
rom[125350] = 12'h222;
rom[125351] = 12'h222;
rom[125352] = 12'h222;
rom[125353] = 12'h222;
rom[125354] = 12'h222;
rom[125355] = 12'h222;
rom[125356] = 12'h222;
rom[125357] = 12'h222;
rom[125358] = 12'h222;
rom[125359] = 12'h222;
rom[125360] = 12'h222;
rom[125361] = 12'h111;
rom[125362] = 12'h111;
rom[125363] = 12'h111;
rom[125364] = 12'h111;
rom[125365] = 12'h111;
rom[125366] = 12'h  0;
rom[125367] = 12'h  0;
rom[125368] = 12'h  0;
rom[125369] = 12'h  0;
rom[125370] = 12'h  0;
rom[125371] = 12'h  0;
rom[125372] = 12'h  0;
rom[125373] = 12'h  0;
rom[125374] = 12'h  0;
rom[125375] = 12'h  0;
rom[125376] = 12'h  0;
rom[125377] = 12'h  0;
rom[125378] = 12'h  0;
rom[125379] = 12'h  0;
rom[125380] = 12'h  0;
rom[125381] = 12'h  0;
rom[125382] = 12'h111;
rom[125383] = 12'h111;
rom[125384] = 12'h111;
rom[125385] = 12'h111;
rom[125386] = 12'h111;
rom[125387] = 12'h111;
rom[125388] = 12'h  0;
rom[125389] = 12'h  0;
rom[125390] = 12'h  0;
rom[125391] = 12'h  0;
rom[125392] = 12'h  0;
rom[125393] = 12'h  0;
rom[125394] = 12'h  0;
rom[125395] = 12'h  0;
rom[125396] = 12'h  0;
rom[125397] = 12'h  0;
rom[125398] = 12'h  0;
rom[125399] = 12'h  0;
rom[125400] = 12'h  0;
rom[125401] = 12'h  0;
rom[125402] = 12'h  0;
rom[125403] = 12'h  0;
rom[125404] = 12'h  0;
rom[125405] = 12'h  0;
rom[125406] = 12'h  0;
rom[125407] = 12'h  0;
rom[125408] = 12'h  0;
rom[125409] = 12'h  0;
rom[125410] = 12'h  0;
rom[125411] = 12'h  0;
rom[125412] = 12'h  0;
rom[125413] = 12'h  0;
rom[125414] = 12'h  0;
rom[125415] = 12'h  0;
rom[125416] = 12'h  0;
rom[125417] = 12'h  0;
rom[125418] = 12'h  0;
rom[125419] = 12'h  0;
rom[125420] = 12'h  0;
rom[125421] = 12'h  0;
rom[125422] = 12'h  0;
rom[125423] = 12'h  0;
rom[125424] = 12'h  0;
rom[125425] = 12'h  0;
rom[125426] = 12'h  0;
rom[125427] = 12'h  0;
rom[125428] = 12'h  0;
rom[125429] = 12'h  0;
rom[125430] = 12'h  0;
rom[125431] = 12'h  0;
rom[125432] = 12'h  0;
rom[125433] = 12'h  0;
rom[125434] = 12'h  0;
rom[125435] = 12'h  0;
rom[125436] = 12'h  0;
rom[125437] = 12'h  0;
rom[125438] = 12'h  0;
rom[125439] = 12'h  0;
rom[125440] = 12'h  0;
rom[125441] = 12'h  0;
rom[125442] = 12'h  0;
rom[125443] = 12'h  0;
rom[125444] = 12'h  0;
rom[125445] = 12'h  0;
rom[125446] = 12'h  0;
rom[125447] = 12'h  0;
rom[125448] = 12'h  0;
rom[125449] = 12'h  0;
rom[125450] = 12'h  0;
rom[125451] = 12'h  0;
rom[125452] = 12'h  0;
rom[125453] = 12'h  0;
rom[125454] = 12'h  0;
rom[125455] = 12'h  0;
rom[125456] = 12'h  0;
rom[125457] = 12'h  0;
rom[125458] = 12'h  0;
rom[125459] = 12'h  0;
rom[125460] = 12'h111;
rom[125461] = 12'h333;
rom[125462] = 12'h888;
rom[125463] = 12'hccc;
rom[125464] = 12'haaa;
rom[125465] = 12'h555;
rom[125466] = 12'h111;
rom[125467] = 12'h  0;
rom[125468] = 12'h  0;
rom[125469] = 12'h  0;
rom[125470] = 12'h  0;
rom[125471] = 12'h  0;
rom[125472] = 12'h  0;
rom[125473] = 12'h  0;
rom[125474] = 12'h  0;
rom[125475] = 12'h  0;
rom[125476] = 12'h  0;
rom[125477] = 12'h  0;
rom[125478] = 12'h111;
rom[125479] = 12'h444;
rom[125480] = 12'h888;
rom[125481] = 12'h777;
rom[125482] = 12'h444;
rom[125483] = 12'h111;
rom[125484] = 12'h  0;
rom[125485] = 12'h  0;
rom[125486] = 12'h  0;
rom[125487] = 12'h  0;
rom[125488] = 12'h  0;
rom[125489] = 12'h  0;
rom[125490] = 12'h  0;
rom[125491] = 12'h  0;
rom[125492] = 12'h  0;
rom[125493] = 12'h111;
rom[125494] = 12'h111;
rom[125495] = 12'h111;
rom[125496] = 12'h  0;
rom[125497] = 12'h  0;
rom[125498] = 12'h  0;
rom[125499] = 12'h  0;
rom[125500] = 12'h  0;
rom[125501] = 12'h  0;
rom[125502] = 12'h  0;
rom[125503] = 12'h  0;
rom[125504] = 12'h  0;
rom[125505] = 12'h  0;
rom[125506] = 12'h  0;
rom[125507] = 12'h  0;
rom[125508] = 12'h  0;
rom[125509] = 12'h  0;
rom[125510] = 12'h  0;
rom[125511] = 12'h  0;
rom[125512] = 12'h  0;
rom[125513] = 12'h  0;
rom[125514] = 12'h  0;
rom[125515] = 12'h  0;
rom[125516] = 12'h  0;
rom[125517] = 12'h  0;
rom[125518] = 12'h  0;
rom[125519] = 12'h  0;
rom[125520] = 12'h222;
rom[125521] = 12'h333;
rom[125522] = 12'h444;
rom[125523] = 12'h333;
rom[125524] = 12'h222;
rom[125525] = 12'h  0;
rom[125526] = 12'h  0;
rom[125527] = 12'h  0;
rom[125528] = 12'h  0;
rom[125529] = 12'h  0;
rom[125530] = 12'h  0;
rom[125531] = 12'h  0;
rom[125532] = 12'h  0;
rom[125533] = 12'h  0;
rom[125534] = 12'h  0;
rom[125535] = 12'h  0;
rom[125536] = 12'h  0;
rom[125537] = 12'h  0;
rom[125538] = 12'h  0;
rom[125539] = 12'h  0;
rom[125540] = 12'h  0;
rom[125541] = 12'h  0;
rom[125542] = 12'h  0;
rom[125543] = 12'h  0;
rom[125544] = 12'h  0;
rom[125545] = 12'h  0;
rom[125546] = 12'h  0;
rom[125547] = 12'h  0;
rom[125548] = 12'h  0;
rom[125549] = 12'h  0;
rom[125550] = 12'h  0;
rom[125551] = 12'h  0;
rom[125552] = 12'h  0;
rom[125553] = 12'h  0;
rom[125554] = 12'h  0;
rom[125555] = 12'h  0;
rom[125556] = 12'h  0;
rom[125557] = 12'h  0;
rom[125558] = 12'h  0;
rom[125559] = 12'h  0;
rom[125560] = 12'h  0;
rom[125561] = 12'h  0;
rom[125562] = 12'h  0;
rom[125563] = 12'h  0;
rom[125564] = 12'h  0;
rom[125565] = 12'h  0;
rom[125566] = 12'h  0;
rom[125567] = 12'h  0;
rom[125568] = 12'h  0;
rom[125569] = 12'h  0;
rom[125570] = 12'h  0;
rom[125571] = 12'h  0;
rom[125572] = 12'h  0;
rom[125573] = 12'h  0;
rom[125574] = 12'h  0;
rom[125575] = 12'h  0;
rom[125576] = 12'h  0;
rom[125577] = 12'h  0;
rom[125578] = 12'h111;
rom[125579] = 12'h222;
rom[125580] = 12'h444;
rom[125581] = 12'h555;
rom[125582] = 12'h444;
rom[125583] = 12'h222;
rom[125584] = 12'h111;
rom[125585] = 12'h  0;
rom[125586] = 12'h  0;
rom[125587] = 12'h  0;
rom[125588] = 12'h  0;
rom[125589] = 12'h  0;
rom[125590] = 12'h  0;
rom[125591] = 12'h  0;
rom[125592] = 12'h  0;
rom[125593] = 12'h  0;
rom[125594] = 12'h  0;
rom[125595] = 12'h  0;
rom[125596] = 12'h  0;
rom[125597] = 12'h  0;
rom[125598] = 12'h  0;
rom[125599] = 12'h  0;
rom[125600] = 12'hccc;
rom[125601] = 12'hccc;
rom[125602] = 12'hccc;
rom[125603] = 12'hccc;
rom[125604] = 12'hccc;
rom[125605] = 12'hccc;
rom[125606] = 12'hbbb;
rom[125607] = 12'hbbb;
rom[125608] = 12'hbbb;
rom[125609] = 12'hbbb;
rom[125610] = 12'hbbb;
rom[125611] = 12'hbbb;
rom[125612] = 12'hbbb;
rom[125613] = 12'haaa;
rom[125614] = 12'haaa;
rom[125615] = 12'haaa;
rom[125616] = 12'haaa;
rom[125617] = 12'haaa;
rom[125618] = 12'haaa;
rom[125619] = 12'haaa;
rom[125620] = 12'haaa;
rom[125621] = 12'haaa;
rom[125622] = 12'haaa;
rom[125623] = 12'haaa;
rom[125624] = 12'h999;
rom[125625] = 12'h999;
rom[125626] = 12'h999;
rom[125627] = 12'h999;
rom[125628] = 12'h999;
rom[125629] = 12'h999;
rom[125630] = 12'h999;
rom[125631] = 12'h999;
rom[125632] = 12'h888;
rom[125633] = 12'h888;
rom[125634] = 12'h888;
rom[125635] = 12'h888;
rom[125636] = 12'h888;
rom[125637] = 12'h888;
rom[125638] = 12'h888;
rom[125639] = 12'h888;
rom[125640] = 12'h888;
rom[125641] = 12'h888;
rom[125642] = 12'h888;
rom[125643] = 12'h777;
rom[125644] = 12'h777;
rom[125645] = 12'h777;
rom[125646] = 12'h777;
rom[125647] = 12'h777;
rom[125648] = 12'h777;
rom[125649] = 12'h777;
rom[125650] = 12'h777;
rom[125651] = 12'h777;
rom[125652] = 12'h777;
rom[125653] = 12'h666;
rom[125654] = 12'h666;
rom[125655] = 12'h666;
rom[125656] = 12'h666;
rom[125657] = 12'h666;
rom[125658] = 12'h666;
rom[125659] = 12'h777;
rom[125660] = 12'h888;
rom[125661] = 12'haaa;
rom[125662] = 12'hddd;
rom[125663] = 12'hfff;
rom[125664] = 12'heee;
rom[125665] = 12'hccc;
rom[125666] = 12'haaa;
rom[125667] = 12'h888;
rom[125668] = 12'h777;
rom[125669] = 12'h666;
rom[125670] = 12'h555;
rom[125671] = 12'h555;
rom[125672] = 12'h555;
rom[125673] = 12'h555;
rom[125674] = 12'h555;
rom[125675] = 12'h555;
rom[125676] = 12'h555;
rom[125677] = 12'h444;
rom[125678] = 12'h555;
rom[125679] = 12'h555;
rom[125680] = 12'h555;
rom[125681] = 12'h666;
rom[125682] = 12'h777;
rom[125683] = 12'h888;
rom[125684] = 12'h888;
rom[125685] = 12'h666;
rom[125686] = 12'h555;
rom[125687] = 12'h555;
rom[125688] = 12'h555;
rom[125689] = 12'h555;
rom[125690] = 12'h555;
rom[125691] = 12'h555;
rom[125692] = 12'h555;
rom[125693] = 12'h444;
rom[125694] = 12'h444;
rom[125695] = 12'h444;
rom[125696] = 12'h444;
rom[125697] = 12'h444;
rom[125698] = 12'h444;
rom[125699] = 12'h444;
rom[125700] = 12'h444;
rom[125701] = 12'h444;
rom[125702] = 12'h444;
rom[125703] = 12'h444;
rom[125704] = 12'h444;
rom[125705] = 12'h444;
rom[125706] = 12'h444;
rom[125707] = 12'h444;
rom[125708] = 12'h444;
rom[125709] = 12'h555;
rom[125710] = 12'h555;
rom[125711] = 12'h666;
rom[125712] = 12'h555;
rom[125713] = 12'h555;
rom[125714] = 12'h555;
rom[125715] = 12'h444;
rom[125716] = 12'h444;
rom[125717] = 12'h444;
rom[125718] = 12'h444;
rom[125719] = 12'h444;
rom[125720] = 12'h444;
rom[125721] = 12'h444;
rom[125722] = 12'h444;
rom[125723] = 12'h444;
rom[125724] = 12'h444;
rom[125725] = 12'h444;
rom[125726] = 12'h333;
rom[125727] = 12'h333;
rom[125728] = 12'h333;
rom[125729] = 12'h333;
rom[125730] = 12'h333;
rom[125731] = 12'h333;
rom[125732] = 12'h444;
rom[125733] = 12'h444;
rom[125734] = 12'h444;
rom[125735] = 12'h444;
rom[125736] = 12'h444;
rom[125737] = 12'h333;
rom[125738] = 12'h333;
rom[125739] = 12'h333;
rom[125740] = 12'h222;
rom[125741] = 12'h222;
rom[125742] = 12'h222;
rom[125743] = 12'h222;
rom[125744] = 12'h222;
rom[125745] = 12'h333;
rom[125746] = 12'h333;
rom[125747] = 12'h333;
rom[125748] = 12'h333;
rom[125749] = 12'h333;
rom[125750] = 12'h222;
rom[125751] = 12'h222;
rom[125752] = 12'h222;
rom[125753] = 12'h222;
rom[125754] = 12'h222;
rom[125755] = 12'h222;
rom[125756] = 12'h222;
rom[125757] = 12'h222;
rom[125758] = 12'h222;
rom[125759] = 12'h222;
rom[125760] = 12'h111;
rom[125761] = 12'h111;
rom[125762] = 12'h111;
rom[125763] = 12'h111;
rom[125764] = 12'h111;
rom[125765] = 12'h111;
rom[125766] = 12'h  0;
rom[125767] = 12'h  0;
rom[125768] = 12'h  0;
rom[125769] = 12'h  0;
rom[125770] = 12'h  0;
rom[125771] = 12'h  0;
rom[125772] = 12'h  0;
rom[125773] = 12'h  0;
rom[125774] = 12'h  0;
rom[125775] = 12'h  0;
rom[125776] = 12'h  0;
rom[125777] = 12'h  0;
rom[125778] = 12'h  0;
rom[125779] = 12'h  0;
rom[125780] = 12'h  0;
rom[125781] = 12'h  0;
rom[125782] = 12'h111;
rom[125783] = 12'h111;
rom[125784] = 12'h111;
rom[125785] = 12'h111;
rom[125786] = 12'h111;
rom[125787] = 12'h  0;
rom[125788] = 12'h  0;
rom[125789] = 12'h  0;
rom[125790] = 12'h  0;
rom[125791] = 12'h  0;
rom[125792] = 12'h  0;
rom[125793] = 12'h  0;
rom[125794] = 12'h  0;
rom[125795] = 12'h  0;
rom[125796] = 12'h  0;
rom[125797] = 12'h  0;
rom[125798] = 12'h  0;
rom[125799] = 12'h  0;
rom[125800] = 12'h  0;
rom[125801] = 12'h  0;
rom[125802] = 12'h  0;
rom[125803] = 12'h  0;
rom[125804] = 12'h  0;
rom[125805] = 12'h  0;
rom[125806] = 12'h  0;
rom[125807] = 12'h  0;
rom[125808] = 12'h  0;
rom[125809] = 12'h  0;
rom[125810] = 12'h  0;
rom[125811] = 12'h  0;
rom[125812] = 12'h  0;
rom[125813] = 12'h  0;
rom[125814] = 12'h  0;
rom[125815] = 12'h  0;
rom[125816] = 12'h  0;
rom[125817] = 12'h  0;
rom[125818] = 12'h  0;
rom[125819] = 12'h  0;
rom[125820] = 12'h  0;
rom[125821] = 12'h  0;
rom[125822] = 12'h  0;
rom[125823] = 12'h  0;
rom[125824] = 12'h  0;
rom[125825] = 12'h  0;
rom[125826] = 12'h  0;
rom[125827] = 12'h  0;
rom[125828] = 12'h  0;
rom[125829] = 12'h  0;
rom[125830] = 12'h  0;
rom[125831] = 12'h  0;
rom[125832] = 12'h  0;
rom[125833] = 12'h  0;
rom[125834] = 12'h  0;
rom[125835] = 12'h  0;
rom[125836] = 12'h  0;
rom[125837] = 12'h  0;
rom[125838] = 12'h  0;
rom[125839] = 12'h  0;
rom[125840] = 12'h  0;
rom[125841] = 12'h  0;
rom[125842] = 12'h  0;
rom[125843] = 12'h  0;
rom[125844] = 12'h  0;
rom[125845] = 12'h  0;
rom[125846] = 12'h  0;
rom[125847] = 12'h  0;
rom[125848] = 12'h  0;
rom[125849] = 12'h  0;
rom[125850] = 12'h  0;
rom[125851] = 12'h  0;
rom[125852] = 12'h  0;
rom[125853] = 12'h  0;
rom[125854] = 12'h  0;
rom[125855] = 12'h  0;
rom[125856] = 12'h  0;
rom[125857] = 12'h  0;
rom[125858] = 12'h  0;
rom[125859] = 12'h  0;
rom[125860] = 12'h111;
rom[125861] = 12'h444;
rom[125862] = 12'h888;
rom[125863] = 12'hbbb;
rom[125864] = 12'h999;
rom[125865] = 12'h444;
rom[125866] = 12'h111;
rom[125867] = 12'h  0;
rom[125868] = 12'h  0;
rom[125869] = 12'h  0;
rom[125870] = 12'h  0;
rom[125871] = 12'h  0;
rom[125872] = 12'h  0;
rom[125873] = 12'h  0;
rom[125874] = 12'h  0;
rom[125875] = 12'h  0;
rom[125876] = 12'h  0;
rom[125877] = 12'h  0;
rom[125878] = 12'h111;
rom[125879] = 12'h444;
rom[125880] = 12'h777;
rom[125881] = 12'h777;
rom[125882] = 12'h444;
rom[125883] = 12'h111;
rom[125884] = 12'h  0;
rom[125885] = 12'h  0;
rom[125886] = 12'h  0;
rom[125887] = 12'h  0;
rom[125888] = 12'h  0;
rom[125889] = 12'h  0;
rom[125890] = 12'h  0;
rom[125891] = 12'h  0;
rom[125892] = 12'h  0;
rom[125893] = 12'h  0;
rom[125894] = 12'h111;
rom[125895] = 12'h111;
rom[125896] = 12'h  0;
rom[125897] = 12'h  0;
rom[125898] = 12'h  0;
rom[125899] = 12'h  0;
rom[125900] = 12'h  0;
rom[125901] = 12'h  0;
rom[125902] = 12'h  0;
rom[125903] = 12'h  0;
rom[125904] = 12'h  0;
rom[125905] = 12'h  0;
rom[125906] = 12'h  0;
rom[125907] = 12'h  0;
rom[125908] = 12'h  0;
rom[125909] = 12'h  0;
rom[125910] = 12'h  0;
rom[125911] = 12'h  0;
rom[125912] = 12'h  0;
rom[125913] = 12'h  0;
rom[125914] = 12'h  0;
rom[125915] = 12'h  0;
rom[125916] = 12'h  0;
rom[125917] = 12'h  0;
rom[125918] = 12'h  0;
rom[125919] = 12'h  0;
rom[125920] = 12'h111;
rom[125921] = 12'h333;
rom[125922] = 12'h444;
rom[125923] = 12'h333;
rom[125924] = 12'h111;
rom[125925] = 12'h  0;
rom[125926] = 12'h  0;
rom[125927] = 12'h  0;
rom[125928] = 12'h  0;
rom[125929] = 12'h  0;
rom[125930] = 12'h  0;
rom[125931] = 12'h  0;
rom[125932] = 12'h  0;
rom[125933] = 12'h  0;
rom[125934] = 12'h  0;
rom[125935] = 12'h  0;
rom[125936] = 12'h  0;
rom[125937] = 12'h  0;
rom[125938] = 12'h  0;
rom[125939] = 12'h  0;
rom[125940] = 12'h  0;
rom[125941] = 12'h  0;
rom[125942] = 12'h  0;
rom[125943] = 12'h  0;
rom[125944] = 12'h  0;
rom[125945] = 12'h  0;
rom[125946] = 12'h  0;
rom[125947] = 12'h  0;
rom[125948] = 12'h  0;
rom[125949] = 12'h  0;
rom[125950] = 12'h  0;
rom[125951] = 12'h  0;
rom[125952] = 12'h  0;
rom[125953] = 12'h  0;
rom[125954] = 12'h  0;
rom[125955] = 12'h  0;
rom[125956] = 12'h  0;
rom[125957] = 12'h  0;
rom[125958] = 12'h  0;
rom[125959] = 12'h  0;
rom[125960] = 12'h  0;
rom[125961] = 12'h  0;
rom[125962] = 12'h  0;
rom[125963] = 12'h  0;
rom[125964] = 12'h  0;
rom[125965] = 12'h  0;
rom[125966] = 12'h  0;
rom[125967] = 12'h  0;
rom[125968] = 12'h  0;
rom[125969] = 12'h  0;
rom[125970] = 12'h  0;
rom[125971] = 12'h  0;
rom[125972] = 12'h  0;
rom[125973] = 12'h  0;
rom[125974] = 12'h  0;
rom[125975] = 12'h  0;
rom[125976] = 12'h  0;
rom[125977] = 12'h  0;
rom[125978] = 12'h111;
rom[125979] = 12'h111;
rom[125980] = 12'h333;
rom[125981] = 12'h555;
rom[125982] = 12'h444;
rom[125983] = 12'h333;
rom[125984] = 12'h111;
rom[125985] = 12'h  0;
rom[125986] = 12'h  0;
rom[125987] = 12'h  0;
rom[125988] = 12'h  0;
rom[125989] = 12'h  0;
rom[125990] = 12'h  0;
rom[125991] = 12'h  0;
rom[125992] = 12'h  0;
rom[125993] = 12'h  0;
rom[125994] = 12'h  0;
rom[125995] = 12'h  0;
rom[125996] = 12'h  0;
rom[125997] = 12'h  0;
rom[125998] = 12'h  0;
rom[125999] = 12'h  0;
rom[126000] = 12'hccc;
rom[126001] = 12'hccc;
rom[126002] = 12'hccc;
rom[126003] = 12'hbbb;
rom[126004] = 12'hbbb;
rom[126005] = 12'hbbb;
rom[126006] = 12'hbbb;
rom[126007] = 12'hbbb;
rom[126008] = 12'hbbb;
rom[126009] = 12'hbbb;
rom[126010] = 12'hbbb;
rom[126011] = 12'hbbb;
rom[126012] = 12'haaa;
rom[126013] = 12'haaa;
rom[126014] = 12'haaa;
rom[126015] = 12'haaa;
rom[126016] = 12'haaa;
rom[126017] = 12'haaa;
rom[126018] = 12'haaa;
rom[126019] = 12'haaa;
rom[126020] = 12'haaa;
rom[126021] = 12'haaa;
rom[126022] = 12'haaa;
rom[126023] = 12'h999;
rom[126024] = 12'h999;
rom[126025] = 12'h999;
rom[126026] = 12'h999;
rom[126027] = 12'h999;
rom[126028] = 12'h999;
rom[126029] = 12'h999;
rom[126030] = 12'h888;
rom[126031] = 12'h888;
rom[126032] = 12'h888;
rom[126033] = 12'h888;
rom[126034] = 12'h888;
rom[126035] = 12'h888;
rom[126036] = 12'h888;
rom[126037] = 12'h888;
rom[126038] = 12'h888;
rom[126039] = 12'h888;
rom[126040] = 12'h888;
rom[126041] = 12'h888;
rom[126042] = 12'h777;
rom[126043] = 12'h777;
rom[126044] = 12'h777;
rom[126045] = 12'h777;
rom[126046] = 12'h777;
rom[126047] = 12'h777;
rom[126048] = 12'h666;
rom[126049] = 12'h666;
rom[126050] = 12'h666;
rom[126051] = 12'h777;
rom[126052] = 12'h777;
rom[126053] = 12'h666;
rom[126054] = 12'h666;
rom[126055] = 12'h666;
rom[126056] = 12'h666;
rom[126057] = 12'h666;
rom[126058] = 12'h777;
rom[126059] = 12'h777;
rom[126060] = 12'h999;
rom[126061] = 12'hccc;
rom[126062] = 12'heee;
rom[126063] = 12'hfff;
rom[126064] = 12'hddd;
rom[126065] = 12'hbbb;
rom[126066] = 12'h888;
rom[126067] = 12'h777;
rom[126068] = 12'h777;
rom[126069] = 12'h666;
rom[126070] = 12'h555;
rom[126071] = 12'h555;
rom[126072] = 12'h555;
rom[126073] = 12'h555;
rom[126074] = 12'h555;
rom[126075] = 12'h555;
rom[126076] = 12'h444;
rom[126077] = 12'h444;
rom[126078] = 12'h444;
rom[126079] = 12'h555;
rom[126080] = 12'h555;
rom[126081] = 12'h666;
rom[126082] = 12'h888;
rom[126083] = 12'h888;
rom[126084] = 12'h666;
rom[126085] = 12'h555;
rom[126086] = 12'h555;
rom[126087] = 12'h555;
rom[126088] = 12'h555;
rom[126089] = 12'h555;
rom[126090] = 12'h555;
rom[126091] = 12'h444;
rom[126092] = 12'h444;
rom[126093] = 12'h444;
rom[126094] = 12'h444;
rom[126095] = 12'h444;
rom[126096] = 12'h444;
rom[126097] = 12'h444;
rom[126098] = 12'h444;
rom[126099] = 12'h444;
rom[126100] = 12'h444;
rom[126101] = 12'h444;
rom[126102] = 12'h444;
rom[126103] = 12'h444;
rom[126104] = 12'h444;
rom[126105] = 12'h444;
rom[126106] = 12'h444;
rom[126107] = 12'h444;
rom[126108] = 12'h444;
rom[126109] = 12'h444;
rom[126110] = 12'h555;
rom[126111] = 12'h555;
rom[126112] = 12'h666;
rom[126113] = 12'h555;
rom[126114] = 12'h555;
rom[126115] = 12'h444;
rom[126116] = 12'h444;
rom[126117] = 12'h444;
rom[126118] = 12'h444;
rom[126119] = 12'h444;
rom[126120] = 12'h444;
rom[126121] = 12'h444;
rom[126122] = 12'h444;
rom[126123] = 12'h444;
rom[126124] = 12'h444;
rom[126125] = 12'h333;
rom[126126] = 12'h333;
rom[126127] = 12'h333;
rom[126128] = 12'h333;
rom[126129] = 12'h333;
rom[126130] = 12'h333;
rom[126131] = 12'h333;
rom[126132] = 12'h444;
rom[126133] = 12'h444;
rom[126134] = 12'h444;
rom[126135] = 12'h555;
rom[126136] = 12'h444;
rom[126137] = 12'h333;
rom[126138] = 12'h333;
rom[126139] = 12'h333;
rom[126140] = 12'h333;
rom[126141] = 12'h222;
rom[126142] = 12'h222;
rom[126143] = 12'h222;
rom[126144] = 12'h333;
rom[126145] = 12'h333;
rom[126146] = 12'h333;
rom[126147] = 12'h333;
rom[126148] = 12'h333;
rom[126149] = 12'h333;
rom[126150] = 12'h222;
rom[126151] = 12'h222;
rom[126152] = 12'h222;
rom[126153] = 12'h222;
rom[126154] = 12'h222;
rom[126155] = 12'h222;
rom[126156] = 12'h222;
rom[126157] = 12'h222;
rom[126158] = 12'h111;
rom[126159] = 12'h111;
rom[126160] = 12'h111;
rom[126161] = 12'h111;
rom[126162] = 12'h111;
rom[126163] = 12'h111;
rom[126164] = 12'h111;
rom[126165] = 12'h  0;
rom[126166] = 12'h  0;
rom[126167] = 12'h  0;
rom[126168] = 12'h  0;
rom[126169] = 12'h  0;
rom[126170] = 12'h  0;
rom[126171] = 12'h  0;
rom[126172] = 12'h  0;
rom[126173] = 12'h  0;
rom[126174] = 12'h  0;
rom[126175] = 12'h  0;
rom[126176] = 12'h  0;
rom[126177] = 12'h  0;
rom[126178] = 12'h  0;
rom[126179] = 12'h  0;
rom[126180] = 12'h  0;
rom[126181] = 12'h  0;
rom[126182] = 12'h111;
rom[126183] = 12'h111;
rom[126184] = 12'h  0;
rom[126185] = 12'h  0;
rom[126186] = 12'h  0;
rom[126187] = 12'h  0;
rom[126188] = 12'h  0;
rom[126189] = 12'h  0;
rom[126190] = 12'h  0;
rom[126191] = 12'h  0;
rom[126192] = 12'h  0;
rom[126193] = 12'h  0;
rom[126194] = 12'h  0;
rom[126195] = 12'h  0;
rom[126196] = 12'h  0;
rom[126197] = 12'h  0;
rom[126198] = 12'h  0;
rom[126199] = 12'h  0;
rom[126200] = 12'h  0;
rom[126201] = 12'h  0;
rom[126202] = 12'h  0;
rom[126203] = 12'h  0;
rom[126204] = 12'h  0;
rom[126205] = 12'h  0;
rom[126206] = 12'h  0;
rom[126207] = 12'h  0;
rom[126208] = 12'h  0;
rom[126209] = 12'h  0;
rom[126210] = 12'h  0;
rom[126211] = 12'h  0;
rom[126212] = 12'h  0;
rom[126213] = 12'h  0;
rom[126214] = 12'h  0;
rom[126215] = 12'h  0;
rom[126216] = 12'h  0;
rom[126217] = 12'h  0;
rom[126218] = 12'h  0;
rom[126219] = 12'h  0;
rom[126220] = 12'h  0;
rom[126221] = 12'h  0;
rom[126222] = 12'h  0;
rom[126223] = 12'h  0;
rom[126224] = 12'h  0;
rom[126225] = 12'h  0;
rom[126226] = 12'h  0;
rom[126227] = 12'h  0;
rom[126228] = 12'h  0;
rom[126229] = 12'h  0;
rom[126230] = 12'h  0;
rom[126231] = 12'h  0;
rom[126232] = 12'h  0;
rom[126233] = 12'h  0;
rom[126234] = 12'h  0;
rom[126235] = 12'h  0;
rom[126236] = 12'h  0;
rom[126237] = 12'h  0;
rom[126238] = 12'h  0;
rom[126239] = 12'h  0;
rom[126240] = 12'h  0;
rom[126241] = 12'h  0;
rom[126242] = 12'h  0;
rom[126243] = 12'h  0;
rom[126244] = 12'h  0;
rom[126245] = 12'h  0;
rom[126246] = 12'h  0;
rom[126247] = 12'h  0;
rom[126248] = 12'h  0;
rom[126249] = 12'h  0;
rom[126250] = 12'h  0;
rom[126251] = 12'h  0;
rom[126252] = 12'h  0;
rom[126253] = 12'h  0;
rom[126254] = 12'h  0;
rom[126255] = 12'h  0;
rom[126256] = 12'h  0;
rom[126257] = 12'h  0;
rom[126258] = 12'h  0;
rom[126259] = 12'h  0;
rom[126260] = 12'h111;
rom[126261] = 12'h555;
rom[126262] = 12'h999;
rom[126263] = 12'haaa;
rom[126264] = 12'h777;
rom[126265] = 12'h444;
rom[126266] = 12'h111;
rom[126267] = 12'h  0;
rom[126268] = 12'h  0;
rom[126269] = 12'h  0;
rom[126270] = 12'h  0;
rom[126271] = 12'h  0;
rom[126272] = 12'h  0;
rom[126273] = 12'h  0;
rom[126274] = 12'h  0;
rom[126275] = 12'h  0;
rom[126276] = 12'h  0;
rom[126277] = 12'h  0;
rom[126278] = 12'h111;
rom[126279] = 12'h444;
rom[126280] = 12'h777;
rom[126281] = 12'h777;
rom[126282] = 12'h444;
rom[126283] = 12'h111;
rom[126284] = 12'h  0;
rom[126285] = 12'h  0;
rom[126286] = 12'h  0;
rom[126287] = 12'h  0;
rom[126288] = 12'h  0;
rom[126289] = 12'h  0;
rom[126290] = 12'h  0;
rom[126291] = 12'h  0;
rom[126292] = 12'h  0;
rom[126293] = 12'h  0;
rom[126294] = 12'h111;
rom[126295] = 12'h111;
rom[126296] = 12'h  0;
rom[126297] = 12'h  0;
rom[126298] = 12'h  0;
rom[126299] = 12'h  0;
rom[126300] = 12'h  0;
rom[126301] = 12'h  0;
rom[126302] = 12'h  0;
rom[126303] = 12'h  0;
rom[126304] = 12'h  0;
rom[126305] = 12'h  0;
rom[126306] = 12'h  0;
rom[126307] = 12'h  0;
rom[126308] = 12'h  0;
rom[126309] = 12'h  0;
rom[126310] = 12'h  0;
rom[126311] = 12'h  0;
rom[126312] = 12'h  0;
rom[126313] = 12'h  0;
rom[126314] = 12'h  0;
rom[126315] = 12'h  0;
rom[126316] = 12'h  0;
rom[126317] = 12'h  0;
rom[126318] = 12'h  0;
rom[126319] = 12'h  0;
rom[126320] = 12'h111;
rom[126321] = 12'h222;
rom[126322] = 12'h333;
rom[126323] = 12'h333;
rom[126324] = 12'h111;
rom[126325] = 12'h  0;
rom[126326] = 12'h  0;
rom[126327] = 12'h  0;
rom[126328] = 12'h  0;
rom[126329] = 12'h  0;
rom[126330] = 12'h  0;
rom[126331] = 12'h  0;
rom[126332] = 12'h  0;
rom[126333] = 12'h  0;
rom[126334] = 12'h  0;
rom[126335] = 12'h  0;
rom[126336] = 12'h  0;
rom[126337] = 12'h  0;
rom[126338] = 12'h  0;
rom[126339] = 12'h  0;
rom[126340] = 12'h  0;
rom[126341] = 12'h  0;
rom[126342] = 12'h  0;
rom[126343] = 12'h  0;
rom[126344] = 12'h  0;
rom[126345] = 12'h  0;
rom[126346] = 12'h  0;
rom[126347] = 12'h  0;
rom[126348] = 12'h  0;
rom[126349] = 12'h  0;
rom[126350] = 12'h  0;
rom[126351] = 12'h  0;
rom[126352] = 12'h  0;
rom[126353] = 12'h  0;
rom[126354] = 12'h  0;
rom[126355] = 12'h  0;
rom[126356] = 12'h  0;
rom[126357] = 12'h  0;
rom[126358] = 12'h  0;
rom[126359] = 12'h  0;
rom[126360] = 12'h  0;
rom[126361] = 12'h  0;
rom[126362] = 12'h  0;
rom[126363] = 12'h  0;
rom[126364] = 12'h  0;
rom[126365] = 12'h  0;
rom[126366] = 12'h  0;
rom[126367] = 12'h  0;
rom[126368] = 12'h  0;
rom[126369] = 12'h  0;
rom[126370] = 12'h  0;
rom[126371] = 12'h  0;
rom[126372] = 12'h  0;
rom[126373] = 12'h  0;
rom[126374] = 12'h  0;
rom[126375] = 12'h  0;
rom[126376] = 12'h  0;
rom[126377] = 12'h  0;
rom[126378] = 12'h  0;
rom[126379] = 12'h111;
rom[126380] = 12'h222;
rom[126381] = 12'h444;
rom[126382] = 12'h444;
rom[126383] = 12'h333;
rom[126384] = 12'h111;
rom[126385] = 12'h111;
rom[126386] = 12'h  0;
rom[126387] = 12'h  0;
rom[126388] = 12'h  0;
rom[126389] = 12'h  0;
rom[126390] = 12'h  0;
rom[126391] = 12'h  0;
rom[126392] = 12'h  0;
rom[126393] = 12'h  0;
rom[126394] = 12'h  0;
rom[126395] = 12'h  0;
rom[126396] = 12'h  0;
rom[126397] = 12'h  0;
rom[126398] = 12'h  0;
rom[126399] = 12'h  0;
rom[126400] = 12'hccc;
rom[126401] = 12'hccc;
rom[126402] = 12'hbbb;
rom[126403] = 12'hbbb;
rom[126404] = 12'hbbb;
rom[126405] = 12'hbbb;
rom[126406] = 12'hbbb;
rom[126407] = 12'hbbb;
rom[126408] = 12'haaa;
rom[126409] = 12'haaa;
rom[126410] = 12'haaa;
rom[126411] = 12'haaa;
rom[126412] = 12'haaa;
rom[126413] = 12'haaa;
rom[126414] = 12'haaa;
rom[126415] = 12'h999;
rom[126416] = 12'h999;
rom[126417] = 12'haaa;
rom[126418] = 12'haaa;
rom[126419] = 12'haaa;
rom[126420] = 12'haaa;
rom[126421] = 12'haaa;
rom[126422] = 12'h999;
rom[126423] = 12'h999;
rom[126424] = 12'h999;
rom[126425] = 12'h999;
rom[126426] = 12'h999;
rom[126427] = 12'h999;
rom[126428] = 12'h888;
rom[126429] = 12'h888;
rom[126430] = 12'h888;
rom[126431] = 12'h888;
rom[126432] = 12'h888;
rom[126433] = 12'h888;
rom[126434] = 12'h888;
rom[126435] = 12'h888;
rom[126436] = 12'h888;
rom[126437] = 12'h888;
rom[126438] = 12'h888;
rom[126439] = 12'h888;
rom[126440] = 12'h888;
rom[126441] = 12'h888;
rom[126442] = 12'h777;
rom[126443] = 12'h777;
rom[126444] = 12'h777;
rom[126445] = 12'h777;
rom[126446] = 12'h777;
rom[126447] = 12'h777;
rom[126448] = 12'h666;
rom[126449] = 12'h666;
rom[126450] = 12'h666;
rom[126451] = 12'h777;
rom[126452] = 12'h777;
rom[126453] = 12'h666;
rom[126454] = 12'h666;
rom[126455] = 12'h666;
rom[126456] = 12'h666;
rom[126457] = 12'h666;
rom[126458] = 12'h777;
rom[126459] = 12'h888;
rom[126460] = 12'hbbb;
rom[126461] = 12'hddd;
rom[126462] = 12'heee;
rom[126463] = 12'heee;
rom[126464] = 12'hccc;
rom[126465] = 12'h999;
rom[126466] = 12'h777;
rom[126467] = 12'h777;
rom[126468] = 12'h777;
rom[126469] = 12'h666;
rom[126470] = 12'h555;
rom[126471] = 12'h555;
rom[126472] = 12'h555;
rom[126473] = 12'h555;
rom[126474] = 12'h555;
rom[126475] = 12'h555;
rom[126476] = 12'h444;
rom[126477] = 12'h444;
rom[126478] = 12'h444;
rom[126479] = 12'h555;
rom[126480] = 12'h666;
rom[126481] = 12'h777;
rom[126482] = 12'h777;
rom[126483] = 12'h777;
rom[126484] = 12'h555;
rom[126485] = 12'h444;
rom[126486] = 12'h555;
rom[126487] = 12'h555;
rom[126488] = 12'h555;
rom[126489] = 12'h555;
rom[126490] = 12'h444;
rom[126491] = 12'h444;
rom[126492] = 12'h444;
rom[126493] = 12'h444;
rom[126494] = 12'h444;
rom[126495] = 12'h444;
rom[126496] = 12'h444;
rom[126497] = 12'h444;
rom[126498] = 12'h444;
rom[126499] = 12'h444;
rom[126500] = 12'h444;
rom[126501] = 12'h444;
rom[126502] = 12'h444;
rom[126503] = 12'h444;
rom[126504] = 12'h444;
rom[126505] = 12'h444;
rom[126506] = 12'h444;
rom[126507] = 12'h444;
rom[126508] = 12'h444;
rom[126509] = 12'h444;
rom[126510] = 12'h444;
rom[126511] = 12'h555;
rom[126512] = 12'h555;
rom[126513] = 12'h666;
rom[126514] = 12'h555;
rom[126515] = 12'h555;
rom[126516] = 12'h444;
rom[126517] = 12'h444;
rom[126518] = 12'h444;
rom[126519] = 12'h444;
rom[126520] = 12'h444;
rom[126521] = 12'h444;
rom[126522] = 12'h444;
rom[126523] = 12'h444;
rom[126524] = 12'h444;
rom[126525] = 12'h333;
rom[126526] = 12'h333;
rom[126527] = 12'h333;
rom[126528] = 12'h333;
rom[126529] = 12'h333;
rom[126530] = 12'h333;
rom[126531] = 12'h333;
rom[126532] = 12'h333;
rom[126533] = 12'h444;
rom[126534] = 12'h444;
rom[126535] = 12'h444;
rom[126536] = 12'h444;
rom[126537] = 12'h444;
rom[126538] = 12'h333;
rom[126539] = 12'h333;
rom[126540] = 12'h333;
rom[126541] = 12'h222;
rom[126542] = 12'h222;
rom[126543] = 12'h222;
rom[126544] = 12'h333;
rom[126545] = 12'h333;
rom[126546] = 12'h333;
rom[126547] = 12'h333;
rom[126548] = 12'h333;
rom[126549] = 12'h333;
rom[126550] = 12'h222;
rom[126551] = 12'h222;
rom[126552] = 12'h222;
rom[126553] = 12'h222;
rom[126554] = 12'h222;
rom[126555] = 12'h222;
rom[126556] = 12'h222;
rom[126557] = 12'h222;
rom[126558] = 12'h111;
rom[126559] = 12'h111;
rom[126560] = 12'h111;
rom[126561] = 12'h111;
rom[126562] = 12'h111;
rom[126563] = 12'h111;
rom[126564] = 12'h111;
rom[126565] = 12'h  0;
rom[126566] = 12'h  0;
rom[126567] = 12'h  0;
rom[126568] = 12'h  0;
rom[126569] = 12'h  0;
rom[126570] = 12'h  0;
rom[126571] = 12'h  0;
rom[126572] = 12'h  0;
rom[126573] = 12'h  0;
rom[126574] = 12'h  0;
rom[126575] = 12'h  0;
rom[126576] = 12'h  0;
rom[126577] = 12'h  0;
rom[126578] = 12'h  0;
rom[126579] = 12'h  0;
rom[126580] = 12'h  0;
rom[126581] = 12'h  0;
rom[126582] = 12'h  0;
rom[126583] = 12'h111;
rom[126584] = 12'h  0;
rom[126585] = 12'h  0;
rom[126586] = 12'h  0;
rom[126587] = 12'h  0;
rom[126588] = 12'h  0;
rom[126589] = 12'h  0;
rom[126590] = 12'h  0;
rom[126591] = 12'h  0;
rom[126592] = 12'h  0;
rom[126593] = 12'h  0;
rom[126594] = 12'h  0;
rom[126595] = 12'h  0;
rom[126596] = 12'h  0;
rom[126597] = 12'h  0;
rom[126598] = 12'h  0;
rom[126599] = 12'h  0;
rom[126600] = 12'h  0;
rom[126601] = 12'h  0;
rom[126602] = 12'h  0;
rom[126603] = 12'h  0;
rom[126604] = 12'h  0;
rom[126605] = 12'h  0;
rom[126606] = 12'h  0;
rom[126607] = 12'h  0;
rom[126608] = 12'h  0;
rom[126609] = 12'h  0;
rom[126610] = 12'h  0;
rom[126611] = 12'h  0;
rom[126612] = 12'h  0;
rom[126613] = 12'h  0;
rom[126614] = 12'h  0;
rom[126615] = 12'h  0;
rom[126616] = 12'h  0;
rom[126617] = 12'h  0;
rom[126618] = 12'h  0;
rom[126619] = 12'h  0;
rom[126620] = 12'h  0;
rom[126621] = 12'h  0;
rom[126622] = 12'h  0;
rom[126623] = 12'h  0;
rom[126624] = 12'h  0;
rom[126625] = 12'h  0;
rom[126626] = 12'h  0;
rom[126627] = 12'h  0;
rom[126628] = 12'h  0;
rom[126629] = 12'h  0;
rom[126630] = 12'h  0;
rom[126631] = 12'h  0;
rom[126632] = 12'h  0;
rom[126633] = 12'h  0;
rom[126634] = 12'h  0;
rom[126635] = 12'h  0;
rom[126636] = 12'h  0;
rom[126637] = 12'h  0;
rom[126638] = 12'h  0;
rom[126639] = 12'h  0;
rom[126640] = 12'h  0;
rom[126641] = 12'h  0;
rom[126642] = 12'h  0;
rom[126643] = 12'h  0;
rom[126644] = 12'h  0;
rom[126645] = 12'h  0;
rom[126646] = 12'h  0;
rom[126647] = 12'h  0;
rom[126648] = 12'h  0;
rom[126649] = 12'h  0;
rom[126650] = 12'h  0;
rom[126651] = 12'h  0;
rom[126652] = 12'h  0;
rom[126653] = 12'h  0;
rom[126654] = 12'h  0;
rom[126655] = 12'h  0;
rom[126656] = 12'h  0;
rom[126657] = 12'h  0;
rom[126658] = 12'h  0;
rom[126659] = 12'h  0;
rom[126660] = 12'h222;
rom[126661] = 12'h666;
rom[126662] = 12'h999;
rom[126663] = 12'haaa;
rom[126664] = 12'h777;
rom[126665] = 12'h333;
rom[126666] = 12'h111;
rom[126667] = 12'h  0;
rom[126668] = 12'h  0;
rom[126669] = 12'h  0;
rom[126670] = 12'h  0;
rom[126671] = 12'h  0;
rom[126672] = 12'h  0;
rom[126673] = 12'h  0;
rom[126674] = 12'h  0;
rom[126675] = 12'h  0;
rom[126676] = 12'h  0;
rom[126677] = 12'h  0;
rom[126678] = 12'h111;
rom[126679] = 12'h333;
rom[126680] = 12'h666;
rom[126681] = 12'h666;
rom[126682] = 12'h444;
rom[126683] = 12'h111;
rom[126684] = 12'h  0;
rom[126685] = 12'h  0;
rom[126686] = 12'h  0;
rom[126687] = 12'h  0;
rom[126688] = 12'h  0;
rom[126689] = 12'h  0;
rom[126690] = 12'h  0;
rom[126691] = 12'h  0;
rom[126692] = 12'h  0;
rom[126693] = 12'h  0;
rom[126694] = 12'h  0;
rom[126695] = 12'h111;
rom[126696] = 12'h  0;
rom[126697] = 12'h  0;
rom[126698] = 12'h  0;
rom[126699] = 12'h  0;
rom[126700] = 12'h  0;
rom[126701] = 12'h  0;
rom[126702] = 12'h  0;
rom[126703] = 12'h  0;
rom[126704] = 12'h  0;
rom[126705] = 12'h  0;
rom[126706] = 12'h  0;
rom[126707] = 12'h  0;
rom[126708] = 12'h  0;
rom[126709] = 12'h  0;
rom[126710] = 12'h  0;
rom[126711] = 12'h  0;
rom[126712] = 12'h  0;
rom[126713] = 12'h  0;
rom[126714] = 12'h  0;
rom[126715] = 12'h  0;
rom[126716] = 12'h  0;
rom[126717] = 12'h  0;
rom[126718] = 12'h  0;
rom[126719] = 12'h  0;
rom[126720] = 12'h111;
rom[126721] = 12'h222;
rom[126722] = 12'h333;
rom[126723] = 12'h222;
rom[126724] = 12'h111;
rom[126725] = 12'h  0;
rom[126726] = 12'h  0;
rom[126727] = 12'h  0;
rom[126728] = 12'h  0;
rom[126729] = 12'h  0;
rom[126730] = 12'h  0;
rom[126731] = 12'h  0;
rom[126732] = 12'h  0;
rom[126733] = 12'h  0;
rom[126734] = 12'h  0;
rom[126735] = 12'h  0;
rom[126736] = 12'h  0;
rom[126737] = 12'h  0;
rom[126738] = 12'h  0;
rom[126739] = 12'h  0;
rom[126740] = 12'h  0;
rom[126741] = 12'h  0;
rom[126742] = 12'h  0;
rom[126743] = 12'h  0;
rom[126744] = 12'h  0;
rom[126745] = 12'h  0;
rom[126746] = 12'h  0;
rom[126747] = 12'h  0;
rom[126748] = 12'h  0;
rom[126749] = 12'h  0;
rom[126750] = 12'h  0;
rom[126751] = 12'h  0;
rom[126752] = 12'h  0;
rom[126753] = 12'h  0;
rom[126754] = 12'h  0;
rom[126755] = 12'h  0;
rom[126756] = 12'h  0;
rom[126757] = 12'h  0;
rom[126758] = 12'h  0;
rom[126759] = 12'h  0;
rom[126760] = 12'h  0;
rom[126761] = 12'h  0;
rom[126762] = 12'h  0;
rom[126763] = 12'h  0;
rom[126764] = 12'h  0;
rom[126765] = 12'h  0;
rom[126766] = 12'h  0;
rom[126767] = 12'h  0;
rom[126768] = 12'h  0;
rom[126769] = 12'h  0;
rom[126770] = 12'h  0;
rom[126771] = 12'h  0;
rom[126772] = 12'h  0;
rom[126773] = 12'h  0;
rom[126774] = 12'h  0;
rom[126775] = 12'h  0;
rom[126776] = 12'h  0;
rom[126777] = 12'h  0;
rom[126778] = 12'h  0;
rom[126779] = 12'h  0;
rom[126780] = 12'h222;
rom[126781] = 12'h333;
rom[126782] = 12'h444;
rom[126783] = 12'h444;
rom[126784] = 12'h111;
rom[126785] = 12'h111;
rom[126786] = 12'h  0;
rom[126787] = 12'h  0;
rom[126788] = 12'h  0;
rom[126789] = 12'h  0;
rom[126790] = 12'h  0;
rom[126791] = 12'h  0;
rom[126792] = 12'h  0;
rom[126793] = 12'h  0;
rom[126794] = 12'h  0;
rom[126795] = 12'h  0;
rom[126796] = 12'h  0;
rom[126797] = 12'h  0;
rom[126798] = 12'h  0;
rom[126799] = 12'h  0;
rom[126800] = 12'hccc;
rom[126801] = 12'hbbb;
rom[126802] = 12'hbbb;
rom[126803] = 12'hbbb;
rom[126804] = 12'hbbb;
rom[126805] = 12'haaa;
rom[126806] = 12'haaa;
rom[126807] = 12'haaa;
rom[126808] = 12'haaa;
rom[126809] = 12'haaa;
rom[126810] = 12'haaa;
rom[126811] = 12'haaa;
rom[126812] = 12'haaa;
rom[126813] = 12'haaa;
rom[126814] = 12'h999;
rom[126815] = 12'h999;
rom[126816] = 12'h999;
rom[126817] = 12'h999;
rom[126818] = 12'haaa;
rom[126819] = 12'haaa;
rom[126820] = 12'haaa;
rom[126821] = 12'haaa;
rom[126822] = 12'h999;
rom[126823] = 12'h999;
rom[126824] = 12'h999;
rom[126825] = 12'h999;
rom[126826] = 12'h999;
rom[126827] = 12'h888;
rom[126828] = 12'h888;
rom[126829] = 12'h888;
rom[126830] = 12'h888;
rom[126831] = 12'h888;
rom[126832] = 12'h888;
rom[126833] = 12'h888;
rom[126834] = 12'h777;
rom[126835] = 12'h777;
rom[126836] = 12'h777;
rom[126837] = 12'h777;
rom[126838] = 12'h777;
rom[126839] = 12'h888;
rom[126840] = 12'h888;
rom[126841] = 12'h777;
rom[126842] = 12'h777;
rom[126843] = 12'h777;
rom[126844] = 12'h777;
rom[126845] = 12'h777;
rom[126846] = 12'h777;
rom[126847] = 12'h777;
rom[126848] = 12'h666;
rom[126849] = 12'h666;
rom[126850] = 12'h777;
rom[126851] = 12'h777;
rom[126852] = 12'h777;
rom[126853] = 12'h777;
rom[126854] = 12'h666;
rom[126855] = 12'h666;
rom[126856] = 12'h666;
rom[126857] = 12'h777;
rom[126858] = 12'h888;
rom[126859] = 12'h999;
rom[126860] = 12'hccc;
rom[126861] = 12'heee;
rom[126862] = 12'heee;
rom[126863] = 12'hddd;
rom[126864] = 12'h999;
rom[126865] = 12'h888;
rom[126866] = 12'h777;
rom[126867] = 12'h777;
rom[126868] = 12'h777;
rom[126869] = 12'h666;
rom[126870] = 12'h555;
rom[126871] = 12'h555;
rom[126872] = 12'h555;
rom[126873] = 12'h555;
rom[126874] = 12'h555;
rom[126875] = 12'h555;
rom[126876] = 12'h555;
rom[126877] = 12'h444;
rom[126878] = 12'h555;
rom[126879] = 12'h555;
rom[126880] = 12'h777;
rom[126881] = 12'h777;
rom[126882] = 12'h777;
rom[126883] = 12'h666;
rom[126884] = 12'h444;
rom[126885] = 12'h444;
rom[126886] = 12'h444;
rom[126887] = 12'h555;
rom[126888] = 12'h555;
rom[126889] = 12'h444;
rom[126890] = 12'h444;
rom[126891] = 12'h444;
rom[126892] = 12'h444;
rom[126893] = 12'h444;
rom[126894] = 12'h444;
rom[126895] = 12'h444;
rom[126896] = 12'h444;
rom[126897] = 12'h444;
rom[126898] = 12'h444;
rom[126899] = 12'h444;
rom[126900] = 12'h444;
rom[126901] = 12'h444;
rom[126902] = 12'h444;
rom[126903] = 12'h444;
rom[126904] = 12'h444;
rom[126905] = 12'h444;
rom[126906] = 12'h444;
rom[126907] = 12'h444;
rom[126908] = 12'h444;
rom[126909] = 12'h444;
rom[126910] = 12'h444;
rom[126911] = 12'h444;
rom[126912] = 12'h555;
rom[126913] = 12'h555;
rom[126914] = 12'h555;
rom[126915] = 12'h555;
rom[126916] = 12'h444;
rom[126917] = 12'h444;
rom[126918] = 12'h444;
rom[126919] = 12'h444;
rom[126920] = 12'h444;
rom[126921] = 12'h444;
rom[126922] = 12'h444;
rom[126923] = 12'h444;
rom[126924] = 12'h444;
rom[126925] = 12'h333;
rom[126926] = 12'h333;
rom[126927] = 12'h333;
rom[126928] = 12'h333;
rom[126929] = 12'h333;
rom[126930] = 12'h333;
rom[126931] = 12'h333;
rom[126932] = 12'h333;
rom[126933] = 12'h333;
rom[126934] = 12'h444;
rom[126935] = 12'h444;
rom[126936] = 12'h444;
rom[126937] = 12'h444;
rom[126938] = 12'h333;
rom[126939] = 12'h333;
rom[126940] = 12'h333;
rom[126941] = 12'h333;
rom[126942] = 12'h222;
rom[126943] = 12'h222;
rom[126944] = 12'h333;
rom[126945] = 12'h333;
rom[126946] = 12'h333;
rom[126947] = 12'h333;
rom[126948] = 12'h333;
rom[126949] = 12'h333;
rom[126950] = 12'h222;
rom[126951] = 12'h222;
rom[126952] = 12'h222;
rom[126953] = 12'h222;
rom[126954] = 12'h222;
rom[126955] = 12'h222;
rom[126956] = 12'h222;
rom[126957] = 12'h111;
rom[126958] = 12'h111;
rom[126959] = 12'h111;
rom[126960] = 12'h111;
rom[126961] = 12'h111;
rom[126962] = 12'h111;
rom[126963] = 12'h111;
rom[126964] = 12'h111;
rom[126965] = 12'h  0;
rom[126966] = 12'h  0;
rom[126967] = 12'h  0;
rom[126968] = 12'h  0;
rom[126969] = 12'h  0;
rom[126970] = 12'h  0;
rom[126971] = 12'h  0;
rom[126972] = 12'h  0;
rom[126973] = 12'h  0;
rom[126974] = 12'h  0;
rom[126975] = 12'h  0;
rom[126976] = 12'h  0;
rom[126977] = 12'h  0;
rom[126978] = 12'h  0;
rom[126979] = 12'h  0;
rom[126980] = 12'h  0;
rom[126981] = 12'h  0;
rom[126982] = 12'h  0;
rom[126983] = 12'h111;
rom[126984] = 12'h  0;
rom[126985] = 12'h  0;
rom[126986] = 12'h  0;
rom[126987] = 12'h  0;
rom[126988] = 12'h  0;
rom[126989] = 12'h  0;
rom[126990] = 12'h  0;
rom[126991] = 12'h  0;
rom[126992] = 12'h  0;
rom[126993] = 12'h  0;
rom[126994] = 12'h  0;
rom[126995] = 12'h  0;
rom[126996] = 12'h  0;
rom[126997] = 12'h  0;
rom[126998] = 12'h  0;
rom[126999] = 12'h  0;
rom[127000] = 12'h  0;
rom[127001] = 12'h  0;
rom[127002] = 12'h  0;
rom[127003] = 12'h  0;
rom[127004] = 12'h  0;
rom[127005] = 12'h  0;
rom[127006] = 12'h  0;
rom[127007] = 12'h  0;
rom[127008] = 12'h  0;
rom[127009] = 12'h  0;
rom[127010] = 12'h  0;
rom[127011] = 12'h  0;
rom[127012] = 12'h  0;
rom[127013] = 12'h  0;
rom[127014] = 12'h  0;
rom[127015] = 12'h  0;
rom[127016] = 12'h  0;
rom[127017] = 12'h  0;
rom[127018] = 12'h  0;
rom[127019] = 12'h  0;
rom[127020] = 12'h  0;
rom[127021] = 12'h  0;
rom[127022] = 12'h  0;
rom[127023] = 12'h  0;
rom[127024] = 12'h  0;
rom[127025] = 12'h  0;
rom[127026] = 12'h  0;
rom[127027] = 12'h  0;
rom[127028] = 12'h  0;
rom[127029] = 12'h  0;
rom[127030] = 12'h  0;
rom[127031] = 12'h  0;
rom[127032] = 12'h  0;
rom[127033] = 12'h  0;
rom[127034] = 12'h  0;
rom[127035] = 12'h  0;
rom[127036] = 12'h  0;
rom[127037] = 12'h  0;
rom[127038] = 12'h  0;
rom[127039] = 12'h  0;
rom[127040] = 12'h  0;
rom[127041] = 12'h  0;
rom[127042] = 12'h  0;
rom[127043] = 12'h  0;
rom[127044] = 12'h  0;
rom[127045] = 12'h  0;
rom[127046] = 12'h  0;
rom[127047] = 12'h  0;
rom[127048] = 12'h  0;
rom[127049] = 12'h  0;
rom[127050] = 12'h  0;
rom[127051] = 12'h  0;
rom[127052] = 12'h  0;
rom[127053] = 12'h  0;
rom[127054] = 12'h  0;
rom[127055] = 12'h  0;
rom[127056] = 12'h  0;
rom[127057] = 12'h  0;
rom[127058] = 12'h  0;
rom[127059] = 12'h  0;
rom[127060] = 12'h222;
rom[127061] = 12'h777;
rom[127062] = 12'haaa;
rom[127063] = 12'h999;
rom[127064] = 12'h666;
rom[127065] = 12'h333;
rom[127066] = 12'h111;
rom[127067] = 12'h111;
rom[127068] = 12'h  0;
rom[127069] = 12'h  0;
rom[127070] = 12'h  0;
rom[127071] = 12'h  0;
rom[127072] = 12'h  0;
rom[127073] = 12'h  0;
rom[127074] = 12'h  0;
rom[127075] = 12'h  0;
rom[127076] = 12'h  0;
rom[127077] = 12'h  0;
rom[127078] = 12'h111;
rom[127079] = 12'h333;
rom[127080] = 12'h555;
rom[127081] = 12'h666;
rom[127082] = 12'h444;
rom[127083] = 12'h111;
rom[127084] = 12'h  0;
rom[127085] = 12'h  0;
rom[127086] = 12'h  0;
rom[127087] = 12'h  0;
rom[127088] = 12'h  0;
rom[127089] = 12'h  0;
rom[127090] = 12'h  0;
rom[127091] = 12'h  0;
rom[127092] = 12'h  0;
rom[127093] = 12'h  0;
rom[127094] = 12'h  0;
rom[127095] = 12'h111;
rom[127096] = 12'h  0;
rom[127097] = 12'h  0;
rom[127098] = 12'h  0;
rom[127099] = 12'h  0;
rom[127100] = 12'h  0;
rom[127101] = 12'h  0;
rom[127102] = 12'h  0;
rom[127103] = 12'h  0;
rom[127104] = 12'h  0;
rom[127105] = 12'h  0;
rom[127106] = 12'h  0;
rom[127107] = 12'h  0;
rom[127108] = 12'h  0;
rom[127109] = 12'h  0;
rom[127110] = 12'h  0;
rom[127111] = 12'h  0;
rom[127112] = 12'h  0;
rom[127113] = 12'h  0;
rom[127114] = 12'h  0;
rom[127115] = 12'h  0;
rom[127116] = 12'h  0;
rom[127117] = 12'h  0;
rom[127118] = 12'h  0;
rom[127119] = 12'h  0;
rom[127120] = 12'h111;
rom[127121] = 12'h222;
rom[127122] = 12'h333;
rom[127123] = 12'h222;
rom[127124] = 12'h111;
rom[127125] = 12'h  0;
rom[127126] = 12'h  0;
rom[127127] = 12'h  0;
rom[127128] = 12'h  0;
rom[127129] = 12'h  0;
rom[127130] = 12'h  0;
rom[127131] = 12'h  0;
rom[127132] = 12'h  0;
rom[127133] = 12'h  0;
rom[127134] = 12'h  0;
rom[127135] = 12'h  0;
rom[127136] = 12'h  0;
rom[127137] = 12'h  0;
rom[127138] = 12'h  0;
rom[127139] = 12'h  0;
rom[127140] = 12'h  0;
rom[127141] = 12'h  0;
rom[127142] = 12'h  0;
rom[127143] = 12'h  0;
rom[127144] = 12'h  0;
rom[127145] = 12'h  0;
rom[127146] = 12'h  0;
rom[127147] = 12'h  0;
rom[127148] = 12'h  0;
rom[127149] = 12'h  0;
rom[127150] = 12'h  0;
rom[127151] = 12'h  0;
rom[127152] = 12'h  0;
rom[127153] = 12'h  0;
rom[127154] = 12'h  0;
rom[127155] = 12'h  0;
rom[127156] = 12'h  0;
rom[127157] = 12'h  0;
rom[127158] = 12'h  0;
rom[127159] = 12'h  0;
rom[127160] = 12'h  0;
rom[127161] = 12'h  0;
rom[127162] = 12'h  0;
rom[127163] = 12'h  0;
rom[127164] = 12'h  0;
rom[127165] = 12'h  0;
rom[127166] = 12'h  0;
rom[127167] = 12'h  0;
rom[127168] = 12'h  0;
rom[127169] = 12'h  0;
rom[127170] = 12'h  0;
rom[127171] = 12'h  0;
rom[127172] = 12'h  0;
rom[127173] = 12'h  0;
rom[127174] = 12'h  0;
rom[127175] = 12'h  0;
rom[127176] = 12'h  0;
rom[127177] = 12'h  0;
rom[127178] = 12'h  0;
rom[127179] = 12'h  0;
rom[127180] = 12'h111;
rom[127181] = 12'h333;
rom[127182] = 12'h444;
rom[127183] = 12'h444;
rom[127184] = 12'h111;
rom[127185] = 12'h111;
rom[127186] = 12'h  0;
rom[127187] = 12'h  0;
rom[127188] = 12'h  0;
rom[127189] = 12'h  0;
rom[127190] = 12'h  0;
rom[127191] = 12'h  0;
rom[127192] = 12'h  0;
rom[127193] = 12'h  0;
rom[127194] = 12'h  0;
rom[127195] = 12'h  0;
rom[127196] = 12'h  0;
rom[127197] = 12'h  0;
rom[127198] = 12'h  0;
rom[127199] = 12'h111;
rom[127200] = 12'hbbb;
rom[127201] = 12'hbbb;
rom[127202] = 12'hbbb;
rom[127203] = 12'hbbb;
rom[127204] = 12'haaa;
rom[127205] = 12'haaa;
rom[127206] = 12'haaa;
rom[127207] = 12'haaa;
rom[127208] = 12'hbbb;
rom[127209] = 12'haaa;
rom[127210] = 12'haaa;
rom[127211] = 12'haaa;
rom[127212] = 12'haaa;
rom[127213] = 12'h999;
rom[127214] = 12'h999;
rom[127215] = 12'h999;
rom[127216] = 12'h999;
rom[127217] = 12'h999;
rom[127218] = 12'haaa;
rom[127219] = 12'haaa;
rom[127220] = 12'haaa;
rom[127221] = 12'haaa;
rom[127222] = 12'h999;
rom[127223] = 12'h999;
rom[127224] = 12'h999;
rom[127225] = 12'h999;
rom[127226] = 12'h888;
rom[127227] = 12'h888;
rom[127228] = 12'h888;
rom[127229] = 12'h888;
rom[127230] = 12'h888;
rom[127231] = 12'h888;
rom[127232] = 12'h888;
rom[127233] = 12'h888;
rom[127234] = 12'h777;
rom[127235] = 12'h777;
rom[127236] = 12'h777;
rom[127237] = 12'h777;
rom[127238] = 12'h777;
rom[127239] = 12'h888;
rom[127240] = 12'h888;
rom[127241] = 12'h777;
rom[127242] = 12'h777;
rom[127243] = 12'h777;
rom[127244] = 12'h777;
rom[127245] = 12'h777;
rom[127246] = 12'h777;
rom[127247] = 12'h777;
rom[127248] = 12'h666;
rom[127249] = 12'h666;
rom[127250] = 12'h777;
rom[127251] = 12'h777;
rom[127252] = 12'h777;
rom[127253] = 12'h777;
rom[127254] = 12'h666;
rom[127255] = 12'h666;
rom[127256] = 12'h777;
rom[127257] = 12'h888;
rom[127258] = 12'h999;
rom[127259] = 12'haaa;
rom[127260] = 12'hddd;
rom[127261] = 12'hfff;
rom[127262] = 12'heee;
rom[127263] = 12'hccc;
rom[127264] = 12'h888;
rom[127265] = 12'h777;
rom[127266] = 12'h777;
rom[127267] = 12'h777;
rom[127268] = 12'h777;
rom[127269] = 12'h666;
rom[127270] = 12'h555;
rom[127271] = 12'h555;
rom[127272] = 12'h666;
rom[127273] = 12'h555;
rom[127274] = 12'h555;
rom[127275] = 12'h555;
rom[127276] = 12'h555;
rom[127277] = 12'h444;
rom[127278] = 12'h555;
rom[127279] = 12'h666;
rom[127280] = 12'h777;
rom[127281] = 12'h777;
rom[127282] = 12'h666;
rom[127283] = 12'h555;
rom[127284] = 12'h444;
rom[127285] = 12'h555;
rom[127286] = 12'h555;
rom[127287] = 12'h444;
rom[127288] = 12'h444;
rom[127289] = 12'h444;
rom[127290] = 12'h555;
rom[127291] = 12'h444;
rom[127292] = 12'h444;
rom[127293] = 12'h444;
rom[127294] = 12'h444;
rom[127295] = 12'h444;
rom[127296] = 12'h444;
rom[127297] = 12'h444;
rom[127298] = 12'h444;
rom[127299] = 12'h444;
rom[127300] = 12'h444;
rom[127301] = 12'h444;
rom[127302] = 12'h444;
rom[127303] = 12'h444;
rom[127304] = 12'h444;
rom[127305] = 12'h444;
rom[127306] = 12'h444;
rom[127307] = 12'h444;
rom[127308] = 12'h444;
rom[127309] = 12'h444;
rom[127310] = 12'h444;
rom[127311] = 12'h444;
rom[127312] = 12'h555;
rom[127313] = 12'h555;
rom[127314] = 12'h555;
rom[127315] = 12'h555;
rom[127316] = 12'h555;
rom[127317] = 12'h555;
rom[127318] = 12'h444;
rom[127319] = 12'h444;
rom[127320] = 12'h444;
rom[127321] = 12'h444;
rom[127322] = 12'h444;
rom[127323] = 12'h444;
rom[127324] = 12'h444;
rom[127325] = 12'h444;
rom[127326] = 12'h333;
rom[127327] = 12'h333;
rom[127328] = 12'h333;
rom[127329] = 12'h333;
rom[127330] = 12'h333;
rom[127331] = 12'h333;
rom[127332] = 12'h333;
rom[127333] = 12'h333;
rom[127334] = 12'h444;
rom[127335] = 12'h444;
rom[127336] = 12'h444;
rom[127337] = 12'h444;
rom[127338] = 12'h333;
rom[127339] = 12'h333;
rom[127340] = 12'h333;
rom[127341] = 12'h333;
rom[127342] = 12'h333;
rom[127343] = 12'h222;
rom[127344] = 12'h333;
rom[127345] = 12'h333;
rom[127346] = 12'h333;
rom[127347] = 12'h333;
rom[127348] = 12'h333;
rom[127349] = 12'h333;
rom[127350] = 12'h222;
rom[127351] = 12'h222;
rom[127352] = 12'h222;
rom[127353] = 12'h222;
rom[127354] = 12'h222;
rom[127355] = 12'h222;
rom[127356] = 12'h222;
rom[127357] = 12'h111;
rom[127358] = 12'h111;
rom[127359] = 12'h111;
rom[127360] = 12'h111;
rom[127361] = 12'h111;
rom[127362] = 12'h111;
rom[127363] = 12'h111;
rom[127364] = 12'h111;
rom[127365] = 12'h  0;
rom[127366] = 12'h  0;
rom[127367] = 12'h  0;
rom[127368] = 12'h  0;
rom[127369] = 12'h  0;
rom[127370] = 12'h  0;
rom[127371] = 12'h  0;
rom[127372] = 12'h  0;
rom[127373] = 12'h  0;
rom[127374] = 12'h  0;
rom[127375] = 12'h  0;
rom[127376] = 12'h  0;
rom[127377] = 12'h  0;
rom[127378] = 12'h  0;
rom[127379] = 12'h  0;
rom[127380] = 12'h  0;
rom[127381] = 12'h  0;
rom[127382] = 12'h  0;
rom[127383] = 12'h  0;
rom[127384] = 12'h  0;
rom[127385] = 12'h  0;
rom[127386] = 12'h  0;
rom[127387] = 12'h  0;
rom[127388] = 12'h  0;
rom[127389] = 12'h  0;
rom[127390] = 12'h  0;
rom[127391] = 12'h  0;
rom[127392] = 12'h  0;
rom[127393] = 12'h  0;
rom[127394] = 12'h  0;
rom[127395] = 12'h  0;
rom[127396] = 12'h  0;
rom[127397] = 12'h  0;
rom[127398] = 12'h  0;
rom[127399] = 12'h  0;
rom[127400] = 12'h  0;
rom[127401] = 12'h  0;
rom[127402] = 12'h  0;
rom[127403] = 12'h  0;
rom[127404] = 12'h  0;
rom[127405] = 12'h  0;
rom[127406] = 12'h  0;
rom[127407] = 12'h  0;
rom[127408] = 12'h  0;
rom[127409] = 12'h  0;
rom[127410] = 12'h  0;
rom[127411] = 12'h  0;
rom[127412] = 12'h  0;
rom[127413] = 12'h  0;
rom[127414] = 12'h  0;
rom[127415] = 12'h  0;
rom[127416] = 12'h  0;
rom[127417] = 12'h  0;
rom[127418] = 12'h  0;
rom[127419] = 12'h  0;
rom[127420] = 12'h  0;
rom[127421] = 12'h  0;
rom[127422] = 12'h  0;
rom[127423] = 12'h  0;
rom[127424] = 12'h  0;
rom[127425] = 12'h  0;
rom[127426] = 12'h  0;
rom[127427] = 12'h  0;
rom[127428] = 12'h  0;
rom[127429] = 12'h  0;
rom[127430] = 12'h  0;
rom[127431] = 12'h  0;
rom[127432] = 12'h  0;
rom[127433] = 12'h  0;
rom[127434] = 12'h  0;
rom[127435] = 12'h  0;
rom[127436] = 12'h  0;
rom[127437] = 12'h  0;
rom[127438] = 12'h  0;
rom[127439] = 12'h  0;
rom[127440] = 12'h  0;
rom[127441] = 12'h  0;
rom[127442] = 12'h  0;
rom[127443] = 12'h  0;
rom[127444] = 12'h  0;
rom[127445] = 12'h  0;
rom[127446] = 12'h  0;
rom[127447] = 12'h  0;
rom[127448] = 12'h  0;
rom[127449] = 12'h  0;
rom[127450] = 12'h  0;
rom[127451] = 12'h  0;
rom[127452] = 12'h  0;
rom[127453] = 12'h  0;
rom[127454] = 12'h  0;
rom[127455] = 12'h  0;
rom[127456] = 12'h  0;
rom[127457] = 12'h  0;
rom[127458] = 12'h  0;
rom[127459] = 12'h111;
rom[127460] = 12'h333;
rom[127461] = 12'h888;
rom[127462] = 12'hbbb;
rom[127463] = 12'h888;
rom[127464] = 12'h666;
rom[127465] = 12'h333;
rom[127466] = 12'h111;
rom[127467] = 12'h111;
rom[127468] = 12'h  0;
rom[127469] = 12'h  0;
rom[127470] = 12'h  0;
rom[127471] = 12'h  0;
rom[127472] = 12'h  0;
rom[127473] = 12'h  0;
rom[127474] = 12'h  0;
rom[127475] = 12'h  0;
rom[127476] = 12'h  0;
rom[127477] = 12'h  0;
rom[127478] = 12'h111;
rom[127479] = 12'h333;
rom[127480] = 12'h555;
rom[127481] = 12'h666;
rom[127482] = 12'h444;
rom[127483] = 12'h111;
rom[127484] = 12'h  0;
rom[127485] = 12'h  0;
rom[127486] = 12'h  0;
rom[127487] = 12'h  0;
rom[127488] = 12'h  0;
rom[127489] = 12'h  0;
rom[127490] = 12'h  0;
rom[127491] = 12'h  0;
rom[127492] = 12'h  0;
rom[127493] = 12'h  0;
rom[127494] = 12'h  0;
rom[127495] = 12'h111;
rom[127496] = 12'h  0;
rom[127497] = 12'h  0;
rom[127498] = 12'h  0;
rom[127499] = 12'h  0;
rom[127500] = 12'h  0;
rom[127501] = 12'h  0;
rom[127502] = 12'h  0;
rom[127503] = 12'h  0;
rom[127504] = 12'h  0;
rom[127505] = 12'h  0;
rom[127506] = 12'h  0;
rom[127507] = 12'h  0;
rom[127508] = 12'h  0;
rom[127509] = 12'h  0;
rom[127510] = 12'h  0;
rom[127511] = 12'h  0;
rom[127512] = 12'h  0;
rom[127513] = 12'h  0;
rom[127514] = 12'h  0;
rom[127515] = 12'h  0;
rom[127516] = 12'h  0;
rom[127517] = 12'h  0;
rom[127518] = 12'h  0;
rom[127519] = 12'h  0;
rom[127520] = 12'h222;
rom[127521] = 12'h333;
rom[127522] = 12'h333;
rom[127523] = 12'h222;
rom[127524] = 12'h  0;
rom[127525] = 12'h  0;
rom[127526] = 12'h  0;
rom[127527] = 12'h  0;
rom[127528] = 12'h  0;
rom[127529] = 12'h  0;
rom[127530] = 12'h  0;
rom[127531] = 12'h  0;
rom[127532] = 12'h  0;
rom[127533] = 12'h  0;
rom[127534] = 12'h  0;
rom[127535] = 12'h  0;
rom[127536] = 12'h  0;
rom[127537] = 12'h  0;
rom[127538] = 12'h  0;
rom[127539] = 12'h  0;
rom[127540] = 12'h  0;
rom[127541] = 12'h  0;
rom[127542] = 12'h  0;
rom[127543] = 12'h  0;
rom[127544] = 12'h  0;
rom[127545] = 12'h  0;
rom[127546] = 12'h  0;
rom[127547] = 12'h  0;
rom[127548] = 12'h  0;
rom[127549] = 12'h  0;
rom[127550] = 12'h  0;
rom[127551] = 12'h  0;
rom[127552] = 12'h  0;
rom[127553] = 12'h  0;
rom[127554] = 12'h  0;
rom[127555] = 12'h  0;
rom[127556] = 12'h  0;
rom[127557] = 12'h  0;
rom[127558] = 12'h  0;
rom[127559] = 12'h  0;
rom[127560] = 12'h  0;
rom[127561] = 12'h  0;
rom[127562] = 12'h  0;
rom[127563] = 12'h  0;
rom[127564] = 12'h  0;
rom[127565] = 12'h  0;
rom[127566] = 12'h  0;
rom[127567] = 12'h  0;
rom[127568] = 12'h  0;
rom[127569] = 12'h  0;
rom[127570] = 12'h  0;
rom[127571] = 12'h  0;
rom[127572] = 12'h  0;
rom[127573] = 12'h  0;
rom[127574] = 12'h  0;
rom[127575] = 12'h  0;
rom[127576] = 12'h  0;
rom[127577] = 12'h  0;
rom[127578] = 12'h  0;
rom[127579] = 12'h  0;
rom[127580] = 12'h111;
rom[127581] = 12'h222;
rom[127582] = 12'h333;
rom[127583] = 12'h444;
rom[127584] = 12'h222;
rom[127585] = 12'h111;
rom[127586] = 12'h  0;
rom[127587] = 12'h  0;
rom[127588] = 12'h  0;
rom[127589] = 12'h  0;
rom[127590] = 12'h  0;
rom[127591] = 12'h  0;
rom[127592] = 12'h  0;
rom[127593] = 12'h  0;
rom[127594] = 12'h  0;
rom[127595] = 12'h  0;
rom[127596] = 12'h  0;
rom[127597] = 12'h  0;
rom[127598] = 12'h  0;
rom[127599] = 12'h111;
rom[127600] = 12'hbbb;
rom[127601] = 12'hbbb;
rom[127602] = 12'hbbb;
rom[127603] = 12'haaa;
rom[127604] = 12'haaa;
rom[127605] = 12'haaa;
rom[127606] = 12'haaa;
rom[127607] = 12'haaa;
rom[127608] = 12'hbbb;
rom[127609] = 12'hbbb;
rom[127610] = 12'haaa;
rom[127611] = 12'haaa;
rom[127612] = 12'haaa;
rom[127613] = 12'h999;
rom[127614] = 12'h999;
rom[127615] = 12'h999;
rom[127616] = 12'h999;
rom[127617] = 12'h999;
rom[127618] = 12'haaa;
rom[127619] = 12'haaa;
rom[127620] = 12'haaa;
rom[127621] = 12'haaa;
rom[127622] = 12'h999;
rom[127623] = 12'h999;
rom[127624] = 12'h999;
rom[127625] = 12'h999;
rom[127626] = 12'h888;
rom[127627] = 12'h888;
rom[127628] = 12'h888;
rom[127629] = 12'h888;
rom[127630] = 12'h888;
rom[127631] = 12'h888;
rom[127632] = 12'h888;
rom[127633] = 12'h777;
rom[127634] = 12'h777;
rom[127635] = 12'h777;
rom[127636] = 12'h777;
rom[127637] = 12'h777;
rom[127638] = 12'h777;
rom[127639] = 12'h888;
rom[127640] = 12'h888;
rom[127641] = 12'h777;
rom[127642] = 12'h777;
rom[127643] = 12'h777;
rom[127644] = 12'h777;
rom[127645] = 12'h777;
rom[127646] = 12'h777;
rom[127647] = 12'h777;
rom[127648] = 12'h666;
rom[127649] = 12'h777;
rom[127650] = 12'h777;
rom[127651] = 12'h777;
rom[127652] = 12'h777;
rom[127653] = 12'h777;
rom[127654] = 12'h666;
rom[127655] = 12'h666;
rom[127656] = 12'h777;
rom[127657] = 12'h888;
rom[127658] = 12'h999;
rom[127659] = 12'hbbb;
rom[127660] = 12'heee;
rom[127661] = 12'hfff;
rom[127662] = 12'heee;
rom[127663] = 12'hccc;
rom[127664] = 12'h888;
rom[127665] = 12'h777;
rom[127666] = 12'h777;
rom[127667] = 12'h777;
rom[127668] = 12'h666;
rom[127669] = 12'h666;
rom[127670] = 12'h666;
rom[127671] = 12'h666;
rom[127672] = 12'h666;
rom[127673] = 12'h555;
rom[127674] = 12'h555;
rom[127675] = 12'h555;
rom[127676] = 12'h555;
rom[127677] = 12'h555;
rom[127678] = 12'h555;
rom[127679] = 12'h666;
rom[127680] = 12'h777;
rom[127681] = 12'h777;
rom[127682] = 12'h555;
rom[127683] = 12'h444;
rom[127684] = 12'h444;
rom[127685] = 12'h555;
rom[127686] = 12'h555;
rom[127687] = 12'h444;
rom[127688] = 12'h444;
rom[127689] = 12'h555;
rom[127690] = 12'h555;
rom[127691] = 12'h444;
rom[127692] = 12'h444;
rom[127693] = 12'h444;
rom[127694] = 12'h444;
rom[127695] = 12'h444;
rom[127696] = 12'h444;
rom[127697] = 12'h444;
rom[127698] = 12'h444;
rom[127699] = 12'h444;
rom[127700] = 12'h444;
rom[127701] = 12'h444;
rom[127702] = 12'h444;
rom[127703] = 12'h444;
rom[127704] = 12'h444;
rom[127705] = 12'h444;
rom[127706] = 12'h444;
rom[127707] = 12'h444;
rom[127708] = 12'h444;
rom[127709] = 12'h444;
rom[127710] = 12'h444;
rom[127711] = 12'h444;
rom[127712] = 12'h555;
rom[127713] = 12'h555;
rom[127714] = 12'h555;
rom[127715] = 12'h555;
rom[127716] = 12'h555;
rom[127717] = 12'h555;
rom[127718] = 12'h444;
rom[127719] = 12'h444;
rom[127720] = 12'h444;
rom[127721] = 12'h555;
rom[127722] = 12'h555;
rom[127723] = 12'h444;
rom[127724] = 12'h444;
rom[127725] = 12'h444;
rom[127726] = 12'h333;
rom[127727] = 12'h333;
rom[127728] = 12'h333;
rom[127729] = 12'h333;
rom[127730] = 12'h333;
rom[127731] = 12'h333;
rom[127732] = 12'h333;
rom[127733] = 12'h444;
rom[127734] = 12'h444;
rom[127735] = 12'h555;
rom[127736] = 12'h444;
rom[127737] = 12'h444;
rom[127738] = 12'h333;
rom[127739] = 12'h333;
rom[127740] = 12'h333;
rom[127741] = 12'h333;
rom[127742] = 12'h333;
rom[127743] = 12'h222;
rom[127744] = 12'h333;
rom[127745] = 12'h333;
rom[127746] = 12'h333;
rom[127747] = 12'h333;
rom[127748] = 12'h333;
rom[127749] = 12'h333;
rom[127750] = 12'h222;
rom[127751] = 12'h222;
rom[127752] = 12'h222;
rom[127753] = 12'h222;
rom[127754] = 12'h222;
rom[127755] = 12'h222;
rom[127756] = 12'h222;
rom[127757] = 12'h111;
rom[127758] = 12'h111;
rom[127759] = 12'h111;
rom[127760] = 12'h111;
rom[127761] = 12'h111;
rom[127762] = 12'h111;
rom[127763] = 12'h111;
rom[127764] = 12'h111;
rom[127765] = 12'h111;
rom[127766] = 12'h  0;
rom[127767] = 12'h  0;
rom[127768] = 12'h  0;
rom[127769] = 12'h  0;
rom[127770] = 12'h  0;
rom[127771] = 12'h  0;
rom[127772] = 12'h  0;
rom[127773] = 12'h  0;
rom[127774] = 12'h  0;
rom[127775] = 12'h  0;
rom[127776] = 12'h  0;
rom[127777] = 12'h  0;
rom[127778] = 12'h  0;
rom[127779] = 12'h  0;
rom[127780] = 12'h  0;
rom[127781] = 12'h  0;
rom[127782] = 12'h  0;
rom[127783] = 12'h  0;
rom[127784] = 12'h  0;
rom[127785] = 12'h  0;
rom[127786] = 12'h  0;
rom[127787] = 12'h  0;
rom[127788] = 12'h  0;
rom[127789] = 12'h  0;
rom[127790] = 12'h  0;
rom[127791] = 12'h  0;
rom[127792] = 12'h  0;
rom[127793] = 12'h  0;
rom[127794] = 12'h  0;
rom[127795] = 12'h  0;
rom[127796] = 12'h  0;
rom[127797] = 12'h  0;
rom[127798] = 12'h  0;
rom[127799] = 12'h  0;
rom[127800] = 12'h  0;
rom[127801] = 12'h  0;
rom[127802] = 12'h  0;
rom[127803] = 12'h  0;
rom[127804] = 12'h  0;
rom[127805] = 12'h  0;
rom[127806] = 12'h  0;
rom[127807] = 12'h  0;
rom[127808] = 12'h  0;
rom[127809] = 12'h  0;
rom[127810] = 12'h  0;
rom[127811] = 12'h  0;
rom[127812] = 12'h  0;
rom[127813] = 12'h  0;
rom[127814] = 12'h  0;
rom[127815] = 12'h  0;
rom[127816] = 12'h  0;
rom[127817] = 12'h  0;
rom[127818] = 12'h  0;
rom[127819] = 12'h  0;
rom[127820] = 12'h  0;
rom[127821] = 12'h  0;
rom[127822] = 12'h  0;
rom[127823] = 12'h  0;
rom[127824] = 12'h  0;
rom[127825] = 12'h  0;
rom[127826] = 12'h  0;
rom[127827] = 12'h  0;
rom[127828] = 12'h  0;
rom[127829] = 12'h  0;
rom[127830] = 12'h  0;
rom[127831] = 12'h  0;
rom[127832] = 12'h  0;
rom[127833] = 12'h  0;
rom[127834] = 12'h  0;
rom[127835] = 12'h  0;
rom[127836] = 12'h  0;
rom[127837] = 12'h  0;
rom[127838] = 12'h  0;
rom[127839] = 12'h  0;
rom[127840] = 12'h  0;
rom[127841] = 12'h  0;
rom[127842] = 12'h  0;
rom[127843] = 12'h  0;
rom[127844] = 12'h  0;
rom[127845] = 12'h  0;
rom[127846] = 12'h  0;
rom[127847] = 12'h  0;
rom[127848] = 12'h  0;
rom[127849] = 12'h  0;
rom[127850] = 12'h  0;
rom[127851] = 12'h  0;
rom[127852] = 12'h  0;
rom[127853] = 12'h  0;
rom[127854] = 12'h  0;
rom[127855] = 12'h  0;
rom[127856] = 12'h  0;
rom[127857] = 12'h  0;
rom[127858] = 12'h  0;
rom[127859] = 12'h111;
rom[127860] = 12'h333;
rom[127861] = 12'h999;
rom[127862] = 12'hbbb;
rom[127863] = 12'h888;
rom[127864] = 12'h555;
rom[127865] = 12'h333;
rom[127866] = 12'h111;
rom[127867] = 12'h  0;
rom[127868] = 12'h  0;
rom[127869] = 12'h  0;
rom[127870] = 12'h  0;
rom[127871] = 12'h  0;
rom[127872] = 12'h  0;
rom[127873] = 12'h  0;
rom[127874] = 12'h  0;
rom[127875] = 12'h  0;
rom[127876] = 12'h  0;
rom[127877] = 12'h  0;
rom[127878] = 12'h111;
rom[127879] = 12'h333;
rom[127880] = 12'h555;
rom[127881] = 12'h666;
rom[127882] = 12'h444;
rom[127883] = 12'h  0;
rom[127884] = 12'h  0;
rom[127885] = 12'h  0;
rom[127886] = 12'h  0;
rom[127887] = 12'h  0;
rom[127888] = 12'h  0;
rom[127889] = 12'h  0;
rom[127890] = 12'h  0;
rom[127891] = 12'h  0;
rom[127892] = 12'h  0;
rom[127893] = 12'h  0;
rom[127894] = 12'h  0;
rom[127895] = 12'h111;
rom[127896] = 12'h  0;
rom[127897] = 12'h  0;
rom[127898] = 12'h  0;
rom[127899] = 12'h  0;
rom[127900] = 12'h  0;
rom[127901] = 12'h  0;
rom[127902] = 12'h  0;
rom[127903] = 12'h  0;
rom[127904] = 12'h  0;
rom[127905] = 12'h  0;
rom[127906] = 12'h  0;
rom[127907] = 12'h  0;
rom[127908] = 12'h  0;
rom[127909] = 12'h  0;
rom[127910] = 12'h  0;
rom[127911] = 12'h  0;
rom[127912] = 12'h  0;
rom[127913] = 12'h  0;
rom[127914] = 12'h  0;
rom[127915] = 12'h  0;
rom[127916] = 12'h  0;
rom[127917] = 12'h  0;
rom[127918] = 12'h  0;
rom[127919] = 12'h  0;
rom[127920] = 12'h222;
rom[127921] = 12'h333;
rom[127922] = 12'h333;
rom[127923] = 12'h222;
rom[127924] = 12'h  0;
rom[127925] = 12'h  0;
rom[127926] = 12'h  0;
rom[127927] = 12'h  0;
rom[127928] = 12'h  0;
rom[127929] = 12'h  0;
rom[127930] = 12'h  0;
rom[127931] = 12'h  0;
rom[127932] = 12'h  0;
rom[127933] = 12'h  0;
rom[127934] = 12'h  0;
rom[127935] = 12'h  0;
rom[127936] = 12'h  0;
rom[127937] = 12'h  0;
rom[127938] = 12'h  0;
rom[127939] = 12'h  0;
rom[127940] = 12'h  0;
rom[127941] = 12'h  0;
rom[127942] = 12'h  0;
rom[127943] = 12'h  0;
rom[127944] = 12'h  0;
rom[127945] = 12'h  0;
rom[127946] = 12'h  0;
rom[127947] = 12'h  0;
rom[127948] = 12'h  0;
rom[127949] = 12'h  0;
rom[127950] = 12'h  0;
rom[127951] = 12'h  0;
rom[127952] = 12'h  0;
rom[127953] = 12'h  0;
rom[127954] = 12'h  0;
rom[127955] = 12'h  0;
rom[127956] = 12'h  0;
rom[127957] = 12'h  0;
rom[127958] = 12'h  0;
rom[127959] = 12'h  0;
rom[127960] = 12'h  0;
rom[127961] = 12'h  0;
rom[127962] = 12'h  0;
rom[127963] = 12'h  0;
rom[127964] = 12'h  0;
rom[127965] = 12'h  0;
rom[127966] = 12'h  0;
rom[127967] = 12'h  0;
rom[127968] = 12'h  0;
rom[127969] = 12'h  0;
rom[127970] = 12'h  0;
rom[127971] = 12'h  0;
rom[127972] = 12'h  0;
rom[127973] = 12'h  0;
rom[127974] = 12'h  0;
rom[127975] = 12'h  0;
rom[127976] = 12'h  0;
rom[127977] = 12'h  0;
rom[127978] = 12'h  0;
rom[127979] = 12'h  0;
rom[127980] = 12'h111;
rom[127981] = 12'h222;
rom[127982] = 12'h333;
rom[127983] = 12'h444;
rom[127984] = 12'h222;
rom[127985] = 12'h111;
rom[127986] = 12'h  0;
rom[127987] = 12'h  0;
rom[127988] = 12'h  0;
rom[127989] = 12'h  0;
rom[127990] = 12'h  0;
rom[127991] = 12'h  0;
rom[127992] = 12'h  0;
rom[127993] = 12'h  0;
rom[127994] = 12'h  0;
rom[127995] = 12'h  0;
rom[127996] = 12'h  0;
rom[127997] = 12'h  0;
rom[127998] = 12'h111;
rom[127999] = 12'h111;
;end
endmodule
