module sber_logo_rom (
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);
  logic [11:0] rom [(128 * 128)];
  assign word = rom[addr];
  initial begin
rom[0] = 12'hfff;
rom[1] = 12'hfff;
rom[2] = 12'hfff;
rom[3] = 12'hfff;
rom[4] = 12'hfff;
rom[5] = 12'hfff;
rom[6] = 12'hfff;
rom[7] = 12'hfff;
rom[8] = 12'hfff;
rom[9] = 12'hfff;
rom[10] = 12'hfff;
rom[11] = 12'hfff;
rom[12] = 12'hfff;
rom[13] = 12'hfff;
rom[14] = 12'hfff;
rom[15] = 12'hfff;
rom[16] = 12'hfff;
rom[17] = 12'hfff;
rom[18] = 12'hfff;
rom[19] = 12'hfff;
rom[20] = 12'hfff;
rom[21] = 12'hfff;
rom[22] = 12'hfff;
rom[23] = 12'hfff;
rom[24] = 12'hfff;
rom[25] = 12'hfff;
rom[26] = 12'hfff;
rom[27] = 12'hfff;
rom[28] = 12'hfff;
rom[29] = 12'hfff;
rom[30] = 12'hfff;
rom[31] = 12'hfff;
rom[32] = 12'hfff;
rom[33] = 12'hfff;
rom[34] = 12'hfff;
rom[35] = 12'hfff;
rom[36] = 12'hfff;
rom[37] = 12'hfff;
rom[38] = 12'hfff;
rom[39] = 12'hfff;
rom[40] = 12'hfff;
rom[41] = 12'hfff;
rom[42] = 12'hfff;
rom[43] = 12'hfff;
rom[44] = 12'hfff;
rom[45] = 12'hfff;
rom[46] = 12'hfff;
rom[47] = 12'hfff;
rom[48] = 12'hfff;
rom[49] = 12'hfff;
rom[50] = 12'hfff;
rom[51] = 12'hfff;
rom[52] = 12'hfff;
rom[53] = 12'hfff;
rom[54] = 12'hfff;
rom[55] = 12'hfff;
rom[56] = 12'hfff;
rom[57] = 12'hfff;
rom[58] = 12'hfff;
rom[59] = 12'hfff;
rom[60] = 12'hfff;
rom[61] = 12'hfff;
rom[62] = 12'hfff;
rom[63] = 12'hfff;
rom[64] = 12'hfff;
rom[65] = 12'hfff;
rom[66] = 12'hfff;
rom[67] = 12'hfff;
rom[68] = 12'hfff;
rom[69] = 12'hfff;
rom[70] = 12'hfff;
rom[71] = 12'hfff;
rom[72] = 12'hfff;
rom[73] = 12'hfff;
rom[74] = 12'hfff;
rom[75] = 12'hfff;
rom[76] = 12'hfff;
rom[77] = 12'hfff;
rom[78] = 12'hfff;
rom[79] = 12'hfff;
rom[80] = 12'hfff;
rom[81] = 12'hfff;
rom[82] = 12'hfff;
rom[83] = 12'hfff;
rom[84] = 12'hfff;
rom[85] = 12'hfff;
rom[86] = 12'hfff;
rom[87] = 12'hfff;
rom[88] = 12'hfff;
rom[89] = 12'hfff;
rom[90] = 12'hfff;
rom[91] = 12'hfff;
rom[92] = 12'hfff;
rom[93] = 12'hfff;
rom[94] = 12'hfff;
rom[95] = 12'hfff;
rom[96] = 12'hfff;
rom[97] = 12'hfff;
rom[98] = 12'hfff;
rom[99] = 12'hfff;
rom[100] = 12'hfff;
rom[101] = 12'hfff;
rom[102] = 12'hfff;
rom[103] = 12'hfff;
rom[104] = 12'hfff;
rom[105] = 12'hfff;
rom[106] = 12'hfff;
rom[107] = 12'hfff;
rom[108] = 12'hfff;
rom[109] = 12'hfff;
rom[110] = 12'hfff;
rom[111] = 12'hfff;
rom[112] = 12'hfff;
rom[113] = 12'hfff;
rom[114] = 12'hfff;
rom[115] = 12'hfff;
rom[116] = 12'hfff;
rom[117] = 12'hfff;
rom[118] = 12'hfff;
rom[119] = 12'hfff;
rom[120] = 12'hfff;
rom[121] = 12'hfff;
rom[122] = 12'hfff;
rom[123] = 12'hfff;
rom[124] = 12'hfff;
rom[125] = 12'hfff;
rom[126] = 12'hfff;
rom[127] = 12'hfff;
rom[128] = 12'hfff;
rom[129] = 12'hfff;
rom[130] = 12'hfff;
rom[131] = 12'hfff;
rom[132] = 12'hfff;
rom[133] = 12'hfff;
rom[134] = 12'hfff;
rom[135] = 12'hfff;
rom[136] = 12'hfff;
rom[137] = 12'hfff;
rom[138] = 12'hfff;
rom[139] = 12'hfff;
rom[140] = 12'hfff;
rom[141] = 12'hfff;
rom[142] = 12'hfff;
rom[143] = 12'hfff;
rom[144] = 12'hfff;
rom[145] = 12'hfff;
rom[146] = 12'hfff;
rom[147] = 12'hfff;
rom[148] = 12'hfff;
rom[149] = 12'hfff;
rom[150] = 12'hfff;
rom[151] = 12'hfff;
rom[152] = 12'hfff;
rom[153] = 12'hfff;
rom[154] = 12'hfff;
rom[155] = 12'hfff;
rom[156] = 12'hfff;
rom[157] = 12'hfff;
rom[158] = 12'hfff;
rom[159] = 12'hfff;
rom[160] = 12'hfff;
rom[161] = 12'hfff;
rom[162] = 12'hfff;
rom[163] = 12'hfff;
rom[164] = 12'hfff;
rom[165] = 12'hfff;
rom[166] = 12'hfff;
rom[167] = 12'hfff;
rom[168] = 12'hfff;
rom[169] = 12'hfff;
rom[170] = 12'hfff;
rom[171] = 12'hfff;
rom[172] = 12'hfff;
rom[173] = 12'hfff;
rom[174] = 12'hfff;
rom[175] = 12'hfff;
rom[176] = 12'hfff;
rom[177] = 12'hfff;
rom[178] = 12'hfff;
rom[179] = 12'hfff;
rom[180] = 12'hfff;
rom[181] = 12'hfff;
rom[182] = 12'hfff;
rom[183] = 12'hfff;
rom[184] = 12'hfff;
rom[185] = 12'hfff;
rom[186] = 12'hfff;
rom[187] = 12'hfff;
rom[188] = 12'hfff;
rom[189] = 12'hfff;
rom[190] = 12'hfff;
rom[191] = 12'hfff;
rom[192] = 12'hfff;
rom[193] = 12'hfff;
rom[194] = 12'hfff;
rom[195] = 12'hfff;
rom[196] = 12'hfff;
rom[197] = 12'hfff;
rom[198] = 12'hfff;
rom[199] = 12'hfff;
rom[200] = 12'hfff;
rom[201] = 12'hfff;
rom[202] = 12'hfff;
rom[203] = 12'hfff;
rom[204] = 12'hfff;
rom[205] = 12'hfff;
rom[206] = 12'hfff;
rom[207] = 12'hfff;
rom[208] = 12'hfff;
rom[209] = 12'hfff;
rom[210] = 12'hfff;
rom[211] = 12'hfff;
rom[212] = 12'hfff;
rom[213] = 12'hfff;
rom[214] = 12'hfff;
rom[215] = 12'hfff;
rom[216] = 12'hfff;
rom[217] = 12'hfff;
rom[218] = 12'hfff;
rom[219] = 12'hfff;
rom[220] = 12'hfff;
rom[221] = 12'hfff;
rom[222] = 12'hfff;
rom[223] = 12'hfff;
rom[224] = 12'hfff;
rom[225] = 12'hfff;
rom[226] = 12'hfff;
rom[227] = 12'hfff;
rom[228] = 12'hfff;
rom[229] = 12'hfff;
rom[230] = 12'hfff;
rom[231] = 12'hfff;
rom[232] = 12'hfff;
rom[233] = 12'hfff;
rom[234] = 12'hfff;
rom[235] = 12'hfff;
rom[236] = 12'hfff;
rom[237] = 12'hfff;
rom[238] = 12'hfff;
rom[239] = 12'hfff;
rom[240] = 12'hfff;
rom[241] = 12'hfff;
rom[242] = 12'hfff;
rom[243] = 12'hfff;
rom[244] = 12'hfff;
rom[245] = 12'hfff;
rom[246] = 12'hfff;
rom[247] = 12'hfff;
rom[248] = 12'hfff;
rom[249] = 12'hfff;
rom[250] = 12'hfff;
rom[251] = 12'hfff;
rom[252] = 12'hfff;
rom[253] = 12'hfff;
rom[254] = 12'hfff;
rom[255] = 12'hfff;
rom[256] = 12'hfff;
rom[257] = 12'hfff;
rom[258] = 12'hfff;
rom[259] = 12'hfff;
rom[260] = 12'hfff;
rom[261] = 12'hfff;
rom[262] = 12'hfff;
rom[263] = 12'hfff;
rom[264] = 12'hfff;
rom[265] = 12'hfff;
rom[266] = 12'hfff;
rom[267] = 12'hfff;
rom[268] = 12'hfff;
rom[269] = 12'hfff;
rom[270] = 12'hfff;
rom[271] = 12'hfff;
rom[272] = 12'hfff;
rom[273] = 12'hfff;
rom[274] = 12'hfff;
rom[275] = 12'hfff;
rom[276] = 12'hfff;
rom[277] = 12'hfff;
rom[278] = 12'hfff;
rom[279] = 12'hfff;
rom[280] = 12'hfff;
rom[281] = 12'hfff;
rom[282] = 12'hfff;
rom[283] = 12'hfff;
rom[284] = 12'hfff;
rom[285] = 12'hfff;
rom[286] = 12'hfff;
rom[287] = 12'hfff;
rom[288] = 12'hfff;
rom[289] = 12'hfff;
rom[290] = 12'hfff;
rom[291] = 12'hfff;
rom[292] = 12'hfff;
rom[293] = 12'hfff;
rom[294] = 12'hfff;
rom[295] = 12'hfff;
rom[296] = 12'hfff;
rom[297] = 12'hfff;
rom[298] = 12'hfff;
rom[299] = 12'hfff;
rom[300] = 12'hfff;
rom[301] = 12'hfff;
rom[302] = 12'hfff;
rom[303] = 12'hfff;
rom[304] = 12'hfff;
rom[305] = 12'hfff;
rom[306] = 12'hfff;
rom[307] = 12'hfff;
rom[308] = 12'hfff;
rom[309] = 12'hfff;
rom[310] = 12'hfff;
rom[311] = 12'hfff;
rom[312] = 12'hfff;
rom[313] = 12'hfff;
rom[314] = 12'hfff;
rom[315] = 12'hfff;
rom[316] = 12'hfff;
rom[317] = 12'hfff;
rom[318] = 12'hfff;
rom[319] = 12'hfff;
rom[320] = 12'hfff;
rom[321] = 12'hfff;
rom[322] = 12'hfff;
rom[323] = 12'hfff;
rom[324] = 12'hfff;
rom[325] = 12'hfff;
rom[326] = 12'hfff;
rom[327] = 12'hfff;
rom[328] = 12'hfff;
rom[329] = 12'hfff;
rom[330] = 12'hfff;
rom[331] = 12'hfff;
rom[332] = 12'hfff;
rom[333] = 12'hfff;
rom[334] = 12'hfff;
rom[335] = 12'hfff;
rom[336] = 12'hfff;
rom[337] = 12'hfff;
rom[338] = 12'hfff;
rom[339] = 12'hfff;
rom[340] = 12'hfff;
rom[341] = 12'hfff;
rom[342] = 12'hfff;
rom[343] = 12'hfff;
rom[344] = 12'hfff;
rom[345] = 12'hfff;
rom[346] = 12'hfff;
rom[347] = 12'hfff;
rom[348] = 12'hfff;
rom[349] = 12'hfff;
rom[350] = 12'hfff;
rom[351] = 12'hfff;
rom[352] = 12'hfff;
rom[353] = 12'hfff;
rom[354] = 12'hfff;
rom[355] = 12'hfff;
rom[356] = 12'hfff;
rom[357] = 12'hfff;
rom[358] = 12'hfff;
rom[359] = 12'hfff;
rom[360] = 12'hfff;
rom[361] = 12'hfff;
rom[362] = 12'hfff;
rom[363] = 12'hfff;
rom[364] = 12'hfff;
rom[365] = 12'hfff;
rom[366] = 12'hfff;
rom[367] = 12'hfff;
rom[368] = 12'hfff;
rom[369] = 12'hfff;
rom[370] = 12'hfff;
rom[371] = 12'hfff;
rom[372] = 12'hfff;
rom[373] = 12'hfff;
rom[374] = 12'hfff;
rom[375] = 12'hfff;
rom[376] = 12'hfff;
rom[377] = 12'hfff;
rom[378] = 12'hfff;
rom[379] = 12'hfff;
rom[380] = 12'hfff;
rom[381] = 12'hfff;
rom[382] = 12'hfff;
rom[383] = 12'hfff;
rom[384] = 12'hfff;
rom[385] = 12'hfff;
rom[386] = 12'hfff;
rom[387] = 12'hfff;
rom[388] = 12'hfff;
rom[389] = 12'hfff;
rom[390] = 12'hfff;
rom[391] = 12'hfff;
rom[392] = 12'hfff;
rom[393] = 12'hfff;
rom[394] = 12'hfff;
rom[395] = 12'hfff;
rom[396] = 12'hfff;
rom[397] = 12'hfff;
rom[398] = 12'hfff;
rom[399] = 12'hfff;
rom[400] = 12'hfff;
rom[401] = 12'hfff;
rom[402] = 12'hfff;
rom[403] = 12'hfff;
rom[404] = 12'hfff;
rom[405] = 12'hfff;
rom[406] = 12'hfff;
rom[407] = 12'hfff;
rom[408] = 12'hfff;
rom[409] = 12'hfff;
rom[410] = 12'hfff;
rom[411] = 12'hfff;
rom[412] = 12'hfff;
rom[413] = 12'hfff;
rom[414] = 12'hfff;
rom[415] = 12'hfff;
rom[416] = 12'hfff;
rom[417] = 12'hfff;
rom[418] = 12'hfff;
rom[419] = 12'hfff;
rom[420] = 12'hfff;
rom[421] = 12'hfff;
rom[422] = 12'hfff;
rom[423] = 12'hfff;
rom[424] = 12'hfff;
rom[425] = 12'hfff;
rom[426] = 12'hfff;
rom[427] = 12'hfff;
rom[428] = 12'hfff;
rom[429] = 12'hfff;
rom[430] = 12'hfff;
rom[431] = 12'hfff;
rom[432] = 12'hfff;
rom[433] = 12'hfff;
rom[434] = 12'hfff;
rom[435] = 12'hfff;
rom[436] = 12'hfff;
rom[437] = 12'hfff;
rom[438] = 12'hfff;
rom[439] = 12'hfff;
rom[440] = 12'hfff;
rom[441] = 12'hfff;
rom[442] = 12'hfff;
rom[443] = 12'hfff;
rom[444] = 12'hfff;
rom[445] = 12'hfff;
rom[446] = 12'hfff;
rom[447] = 12'hfff;
rom[448] = 12'hfff;
rom[449] = 12'hfff;
rom[450] = 12'hfff;
rom[451] = 12'hfff;
rom[452] = 12'hfff;
rom[453] = 12'hfff;
rom[454] = 12'hfff;
rom[455] = 12'hfff;
rom[456] = 12'hfff;
rom[457] = 12'hfff;
rom[458] = 12'hfff;
rom[459] = 12'hfff;
rom[460] = 12'hfff;
rom[461] = 12'hfff;
rom[462] = 12'hfff;
rom[463] = 12'hfff;
rom[464] = 12'hfff;
rom[465] = 12'hfff;
rom[466] = 12'hfff;
rom[467] = 12'hfff;
rom[468] = 12'hfff;
rom[469] = 12'hfff;
rom[470] = 12'hfff;
rom[471] = 12'hfff;
rom[472] = 12'hfff;
rom[473] = 12'hfff;
rom[474] = 12'hfff;
rom[475] = 12'hfff;
rom[476] = 12'hfff;
rom[477] = 12'hfff;
rom[478] = 12'hfff;
rom[479] = 12'hfff;
rom[480] = 12'hfff;
rom[481] = 12'hfff;
rom[482] = 12'hfff;
rom[483] = 12'hfff;
rom[484] = 12'hfff;
rom[485] = 12'hfff;
rom[486] = 12'hfff;
rom[487] = 12'hfff;
rom[488] = 12'hfff;
rom[489] = 12'hfff;
rom[490] = 12'hfff;
rom[491] = 12'hfff;
rom[492] = 12'hfff;
rom[493] = 12'hfff;
rom[494] = 12'hfff;
rom[495] = 12'hfff;
rom[496] = 12'hfff;
rom[497] = 12'hfff;
rom[498] = 12'hfff;
rom[499] = 12'hfff;
rom[500] = 12'hfff;
rom[501] = 12'hfff;
rom[502] = 12'hfff;
rom[503] = 12'hfff;
rom[504] = 12'hfff;
rom[505] = 12'hfff;
rom[506] = 12'hfff;
rom[507] = 12'hfff;
rom[508] = 12'hfff;
rom[509] = 12'hfff;
rom[510] = 12'hfff;
rom[511] = 12'hfff;
rom[512] = 12'hfff;
rom[513] = 12'hfff;
rom[514] = 12'hfff;
rom[515] = 12'hfff;
rom[516] = 12'hfff;
rom[517] = 12'hfff;
rom[518] = 12'hfff;
rom[519] = 12'hfff;
rom[520] = 12'hfff;
rom[521] = 12'hfff;
rom[522] = 12'hfff;
rom[523] = 12'hfff;
rom[524] = 12'hfff;
rom[525] = 12'hfff;
rom[526] = 12'hfff;
rom[527] = 12'hfff;
rom[528] = 12'hfff;
rom[529] = 12'hfff;
rom[530] = 12'hfff;
rom[531] = 12'hfff;
rom[532] = 12'hfff;
rom[533] = 12'hfff;
rom[534] = 12'hfff;
rom[535] = 12'hfff;
rom[536] = 12'hfff;
rom[537] = 12'hfff;
rom[538] = 12'hfff;
rom[539] = 12'hfff;
rom[540] = 12'hfff;
rom[541] = 12'hfff;
rom[542] = 12'hfff;
rom[543] = 12'hfff;
rom[544] = 12'hfff;
rom[545] = 12'hfff;
rom[546] = 12'hfff;
rom[547] = 12'hfff;
rom[548] = 12'hfff;
rom[549] = 12'hfff;
rom[550] = 12'hfff;
rom[551] = 12'hfff;
rom[552] = 12'hfff;
rom[553] = 12'hfff;
rom[554] = 12'hfff;
rom[555] = 12'hfff;
rom[556] = 12'hfff;
rom[557] = 12'hfff;
rom[558] = 12'hfff;
rom[559] = 12'hfff;
rom[560] = 12'hfff;
rom[561] = 12'hfff;
rom[562] = 12'hfff;
rom[563] = 12'hfff;
rom[564] = 12'hfff;
rom[565] = 12'hfff;
rom[566] = 12'hfff;
rom[567] = 12'hfff;
rom[568] = 12'hfff;
rom[569] = 12'hfff;
rom[570] = 12'hfff;
rom[571] = 12'hfff;
rom[572] = 12'hfff;
rom[573] = 12'hfff;
rom[574] = 12'hfff;
rom[575] = 12'hfff;
rom[576] = 12'hfff;
rom[577] = 12'hfff;
rom[578] = 12'hfff;
rom[579] = 12'hfff;
rom[580] = 12'hfff;
rom[581] = 12'hfff;
rom[582] = 12'hfff;
rom[583] = 12'hfff;
rom[584] = 12'hfff;
rom[585] = 12'hfff;
rom[586] = 12'hfff;
rom[587] = 12'hfff;
rom[588] = 12'hfff;
rom[589] = 12'hfff;
rom[590] = 12'hfff;
rom[591] = 12'hfff;
rom[592] = 12'hfff;
rom[593] = 12'hfff;
rom[594] = 12'hfff;
rom[595] = 12'hfff;
rom[596] = 12'hfff;
rom[597] = 12'hfff;
rom[598] = 12'hfff;
rom[599] = 12'hfff;
rom[600] = 12'hfff;
rom[601] = 12'hfff;
rom[602] = 12'hfff;
rom[603] = 12'hfff;
rom[604] = 12'hfff;
rom[605] = 12'hfff;
rom[606] = 12'hfff;
rom[607] = 12'hfff;
rom[608] = 12'hfff;
rom[609] = 12'hfff;
rom[610] = 12'hfff;
rom[611] = 12'hfff;
rom[612] = 12'hfff;
rom[613] = 12'hfff;
rom[614] = 12'hfff;
rom[615] = 12'hfff;
rom[616] = 12'hfff;
rom[617] = 12'hfff;
rom[618] = 12'hfff;
rom[619] = 12'hfff;
rom[620] = 12'hfff;
rom[621] = 12'hfff;
rom[622] = 12'hfff;
rom[623] = 12'hfff;
rom[624] = 12'hfff;
rom[625] = 12'hfff;
rom[626] = 12'hfff;
rom[627] = 12'hfff;
rom[628] = 12'hfff;
rom[629] = 12'hfff;
rom[630] = 12'hfff;
rom[631] = 12'hfff;
rom[632] = 12'hfff;
rom[633] = 12'hfff;
rom[634] = 12'hfff;
rom[635] = 12'hfff;
rom[636] = 12'hfff;
rom[637] = 12'hfff;
rom[638] = 12'hfff;
rom[639] = 12'hfff;
rom[640] = 12'hfff;
rom[641] = 12'hfff;
rom[642] = 12'hfff;
rom[643] = 12'hfff;
rom[644] = 12'hfff;
rom[645] = 12'hfff;
rom[646] = 12'hfff;
rom[647] = 12'hfff;
rom[648] = 12'hfff;
rom[649] = 12'hfff;
rom[650] = 12'hfff;
rom[651] = 12'hfff;
rom[652] = 12'hfff;
rom[653] = 12'hfff;
rom[654] = 12'hfff;
rom[655] = 12'hfff;
rom[656] = 12'hfff;
rom[657] = 12'hfff;
rom[658] = 12'hfff;
rom[659] = 12'hfff;
rom[660] = 12'hfff;
rom[661] = 12'hfff;
rom[662] = 12'hfff;
rom[663] = 12'hfff;
rom[664] = 12'hfff;
rom[665] = 12'hfff;
rom[666] = 12'hfff;
rom[667] = 12'hfff;
rom[668] = 12'hfff;
rom[669] = 12'hfff;
rom[670] = 12'hfff;
rom[671] = 12'hfff;
rom[672] = 12'hfff;
rom[673] = 12'hfff;
rom[674] = 12'hfff;
rom[675] = 12'hfff;
rom[676] = 12'hfff;
rom[677] = 12'hfff;
rom[678] = 12'hfff;
rom[679] = 12'hfff;
rom[680] = 12'hfff;
rom[681] = 12'hfff;
rom[682] = 12'hfff;
rom[683] = 12'hfff;
rom[684] = 12'hfff;
rom[685] = 12'hfff;
rom[686] = 12'hfff;
rom[687] = 12'hfff;
rom[688] = 12'hfff;
rom[689] = 12'hfff;
rom[690] = 12'hfff;
rom[691] = 12'hfff;
rom[692] = 12'hfff;
rom[693] = 12'hfff;
rom[694] = 12'hfff;
rom[695] = 12'hfff;
rom[696] = 12'hfff;
rom[697] = 12'hfff;
rom[698] = 12'hfff;
rom[699] = 12'hfff;
rom[700] = 12'hfff;
rom[701] = 12'hfff;
rom[702] = 12'hfff;
rom[703] = 12'hfff;
rom[704] = 12'hfff;
rom[705] = 12'hfff;
rom[706] = 12'hfff;
rom[707] = 12'hfff;
rom[708] = 12'hfff;
rom[709] = 12'hfff;
rom[710] = 12'hfff;
rom[711] = 12'hfff;
rom[712] = 12'hfff;
rom[713] = 12'hfff;
rom[714] = 12'hfff;
rom[715] = 12'hfff;
rom[716] = 12'hfff;
rom[717] = 12'hfff;
rom[718] = 12'hfff;
rom[719] = 12'hfff;
rom[720] = 12'hfff;
rom[721] = 12'hfff;
rom[722] = 12'hfff;
rom[723] = 12'hfff;
rom[724] = 12'hfff;
rom[725] = 12'hfff;
rom[726] = 12'hfff;
rom[727] = 12'hfff;
rom[728] = 12'hfff;
rom[729] = 12'hfff;
rom[730] = 12'hfff;
rom[731] = 12'hfff;
rom[732] = 12'hfff;
rom[733] = 12'hfff;
rom[734] = 12'hfff;
rom[735] = 12'hfff;
rom[736] = 12'hfff;
rom[737] = 12'hfff;
rom[738] = 12'hfff;
rom[739] = 12'hfff;
rom[740] = 12'hfff;
rom[741] = 12'hfff;
rom[742] = 12'hfff;
rom[743] = 12'hfff;
rom[744] = 12'hfff;
rom[745] = 12'hfff;
rom[746] = 12'hfff;
rom[747] = 12'hfff;
rom[748] = 12'hfff;
rom[749] = 12'hfff;
rom[750] = 12'hfff;
rom[751] = 12'hfff;
rom[752] = 12'hfff;
rom[753] = 12'hfff;
rom[754] = 12'hfff;
rom[755] = 12'hfff;
rom[756] = 12'hfff;
rom[757] = 12'hfff;
rom[758] = 12'hfff;
rom[759] = 12'hfff;
rom[760] = 12'hfff;
rom[761] = 12'hfff;
rom[762] = 12'hfff;
rom[763] = 12'hfff;
rom[764] = 12'hfff;
rom[765] = 12'hfff;
rom[766] = 12'hfff;
rom[767] = 12'hfff;
rom[768] = 12'hfff;
rom[769] = 12'hfff;
rom[770] = 12'hfff;
rom[771] = 12'hfff;
rom[772] = 12'hfff;
rom[773] = 12'hfff;
rom[774] = 12'hfff;
rom[775] = 12'hfff;
rom[776] = 12'hfff;
rom[777] = 12'hfff;
rom[778] = 12'hfff;
rom[779] = 12'hfff;
rom[780] = 12'hfff;
rom[781] = 12'hfff;
rom[782] = 12'hfff;
rom[783] = 12'hfff;
rom[784] = 12'hfff;
rom[785] = 12'hfff;
rom[786] = 12'hfff;
rom[787] = 12'hfff;
rom[788] = 12'hfff;
rom[789] = 12'hfff;
rom[790] = 12'hfff;
rom[791] = 12'hfff;
rom[792] = 12'hfff;
rom[793] = 12'hfff;
rom[794] = 12'hfff;
rom[795] = 12'hfff;
rom[796] = 12'hfff;
rom[797] = 12'hfff;
rom[798] = 12'hfff;
rom[799] = 12'hfff;
rom[800] = 12'hfff;
rom[801] = 12'hfff;
rom[802] = 12'hfff;
rom[803] = 12'hfff;
rom[804] = 12'hfff;
rom[805] = 12'hfff;
rom[806] = 12'hfff;
rom[807] = 12'hfff;
rom[808] = 12'hfff;
rom[809] = 12'hfff;
rom[810] = 12'hfff;
rom[811] = 12'hfff;
rom[812] = 12'hfff;
rom[813] = 12'hfff;
rom[814] = 12'hfff;
rom[815] = 12'hfff;
rom[816] = 12'hfff;
rom[817] = 12'hfff;
rom[818] = 12'hfff;
rom[819] = 12'hfff;
rom[820] = 12'hfff;
rom[821] = 12'hfff;
rom[822] = 12'hfff;
rom[823] = 12'hfff;
rom[824] = 12'hfff;
rom[825] = 12'hfff;
rom[826] = 12'hfff;
rom[827] = 12'hfff;
rom[828] = 12'hfff;
rom[829] = 12'hfff;
rom[830] = 12'hfff;
rom[831] = 12'hfff;
rom[832] = 12'hfff;
rom[833] = 12'hfff;
rom[834] = 12'hfff;
rom[835] = 12'hfff;
rom[836] = 12'hfff;
rom[837] = 12'hfff;
rom[838] = 12'hfff;
rom[839] = 12'hfff;
rom[840] = 12'hfff;
rom[841] = 12'hfff;
rom[842] = 12'hfff;
rom[843] = 12'hfff;
rom[844] = 12'hfff;
rom[845] = 12'hfff;
rom[846] = 12'hfff;
rom[847] = 12'hfff;
rom[848] = 12'hfff;
rom[849] = 12'hfff;
rom[850] = 12'hfff;
rom[851] = 12'hfff;
rom[852] = 12'hfff;
rom[853] = 12'hfff;
rom[854] = 12'hfff;
rom[855] = 12'hfff;
rom[856] = 12'hfff;
rom[857] = 12'hfff;
rom[858] = 12'hfff;
rom[859] = 12'hfff;
rom[860] = 12'hfff;
rom[861] = 12'hfff;
rom[862] = 12'hfff;
rom[863] = 12'hfff;
rom[864] = 12'hfff;
rom[865] = 12'hfff;
rom[866] = 12'hfff;
rom[867] = 12'hfff;
rom[868] = 12'hfff;
rom[869] = 12'hfff;
rom[870] = 12'hfff;
rom[871] = 12'hfff;
rom[872] = 12'hfff;
rom[873] = 12'hfff;
rom[874] = 12'hfff;
rom[875] = 12'hfff;
rom[876] = 12'hfff;
rom[877] = 12'hfff;
rom[878] = 12'hfff;
rom[879] = 12'hfff;
rom[880] = 12'hfff;
rom[881] = 12'hfff;
rom[882] = 12'hfff;
rom[883] = 12'hfff;
rom[884] = 12'hfff;
rom[885] = 12'hfff;
rom[886] = 12'hfff;
rom[887] = 12'hfff;
rom[888] = 12'hfff;
rom[889] = 12'hfff;
rom[890] = 12'hfff;
rom[891] = 12'hfff;
rom[892] = 12'hfff;
rom[893] = 12'hfff;
rom[894] = 12'hfff;
rom[895] = 12'hfff;
rom[896] = 12'hfff;
rom[897] = 12'hfff;
rom[898] = 12'hfff;
rom[899] = 12'hfff;
rom[900] = 12'hfff;
rom[901] = 12'hfff;
rom[902] = 12'hfff;
rom[903] = 12'hfff;
rom[904] = 12'hfff;
rom[905] = 12'hfff;
rom[906] = 12'hfff;
rom[907] = 12'hfff;
rom[908] = 12'hfff;
rom[909] = 12'hfff;
rom[910] = 12'hfff;
rom[911] = 12'hfff;
rom[912] = 12'hfff;
rom[913] = 12'hfff;
rom[914] = 12'hfff;
rom[915] = 12'hfff;
rom[916] = 12'hfff;
rom[917] = 12'hfff;
rom[918] = 12'hfff;
rom[919] = 12'hfff;
rom[920] = 12'hfff;
rom[921] = 12'hfff;
rom[922] = 12'hfff;
rom[923] = 12'hfff;
rom[924] = 12'hfff;
rom[925] = 12'hfff;
rom[926] = 12'hfff;
rom[927] = 12'hfff;
rom[928] = 12'hfff;
rom[929] = 12'hfff;
rom[930] = 12'hfff;
rom[931] = 12'hfff;
rom[932] = 12'hfff;
rom[933] = 12'hfff;
rom[934] = 12'hfff;
rom[935] = 12'hfff;
rom[936] = 12'hfff;
rom[937] = 12'hfff;
rom[938] = 12'hfff;
rom[939] = 12'hfff;
rom[940] = 12'hfff;
rom[941] = 12'hfff;
rom[942] = 12'hfff;
rom[943] = 12'hfff;
rom[944] = 12'hfff;
rom[945] = 12'hfff;
rom[946] = 12'hfff;
rom[947] = 12'hfff;
rom[948] = 12'hfff;
rom[949] = 12'hfff;
rom[950] = 12'hfff;
rom[951] = 12'hfff;
rom[952] = 12'hfff;
rom[953] = 12'hfff;
rom[954] = 12'hfff;
rom[955] = 12'hfff;
rom[956] = 12'hfff;
rom[957] = 12'hfff;
rom[958] = 12'hfff;
rom[959] = 12'hfff;
rom[960] = 12'hfff;
rom[961] = 12'hfff;
rom[962] = 12'hfff;
rom[963] = 12'hfff;
rom[964] = 12'hfff;
rom[965] = 12'hfff;
rom[966] = 12'hfff;
rom[967] = 12'hfff;
rom[968] = 12'hfff;
rom[969] = 12'hfff;
rom[970] = 12'hfff;
rom[971] = 12'hfff;
rom[972] = 12'hfff;
rom[973] = 12'hfff;
rom[974] = 12'hfff;
rom[975] = 12'hfff;
rom[976] = 12'hfff;
rom[977] = 12'hfff;
rom[978] = 12'hfff;
rom[979] = 12'hfff;
rom[980] = 12'hfff;
rom[981] = 12'hfff;
rom[982] = 12'hfff;
rom[983] = 12'hfff;
rom[984] = 12'hfff;
rom[985] = 12'hfff;
rom[986] = 12'hfff;
rom[987] = 12'hfff;
rom[988] = 12'hfff;
rom[989] = 12'hfff;
rom[990] = 12'hfff;
rom[991] = 12'hfff;
rom[992] = 12'hfff;
rom[993] = 12'hfff;
rom[994] = 12'hfff;
rom[995] = 12'hfff;
rom[996] = 12'hfff;
rom[997] = 12'hfff;
rom[998] = 12'hfff;
rom[999] = 12'hfff;
rom[1000] = 12'hfff;
rom[1001] = 12'hfff;
rom[1002] = 12'hfff;
rom[1003] = 12'hfff;
rom[1004] = 12'hfff;
rom[1005] = 12'hfff;
rom[1006] = 12'hfff;
rom[1007] = 12'hfff;
rom[1008] = 12'hfff;
rom[1009] = 12'hfff;
rom[1010] = 12'hfff;
rom[1011] = 12'hfff;
rom[1012] = 12'hfff;
rom[1013] = 12'hfff;
rom[1014] = 12'hfff;
rom[1015] = 12'hfff;
rom[1016] = 12'hfff;
rom[1017] = 12'hfff;
rom[1018] = 12'hfff;
rom[1019] = 12'hfff;
rom[1020] = 12'hfff;
rom[1021] = 12'hfff;
rom[1022] = 12'hfff;
rom[1023] = 12'hfff;
rom[1024] = 12'hfff;
rom[1025] = 12'hfff;
rom[1026] = 12'hfff;
rom[1027] = 12'hfff;
rom[1028] = 12'hfff;
rom[1029] = 12'hfff;
rom[1030] = 12'hfff;
rom[1031] = 12'hfff;
rom[1032] = 12'hfff;
rom[1033] = 12'hfff;
rom[1034] = 12'hfff;
rom[1035] = 12'hfff;
rom[1036] = 12'hfff;
rom[1037] = 12'hfff;
rom[1038] = 12'hfff;
rom[1039] = 12'hfff;
rom[1040] = 12'hfff;
rom[1041] = 12'hfff;
rom[1042] = 12'hfff;
rom[1043] = 12'hfff;
rom[1044] = 12'hfff;
rom[1045] = 12'hfff;
rom[1046] = 12'hfff;
rom[1047] = 12'hfff;
rom[1048] = 12'hfff;
rom[1049] = 12'hfff;
rom[1050] = 12'hfff;
rom[1051] = 12'hfff;
rom[1052] = 12'hfff;
rom[1053] = 12'hfff;
rom[1054] = 12'hfff;
rom[1055] = 12'hfff;
rom[1056] = 12'hfff;
rom[1057] = 12'hfff;
rom[1058] = 12'hfff;
rom[1059] = 12'hfff;
rom[1060] = 12'hfff;
rom[1061] = 12'hfff;
rom[1062] = 12'hfff;
rom[1063] = 12'hfff;
rom[1064] = 12'hfff;
rom[1065] = 12'hfff;
rom[1066] = 12'hfff;
rom[1067] = 12'hfff;
rom[1068] = 12'hfff;
rom[1069] = 12'hfff;
rom[1070] = 12'hfff;
rom[1071] = 12'hfff;
rom[1072] = 12'hfff;
rom[1073] = 12'hfff;
rom[1074] = 12'hfff;
rom[1075] = 12'hfff;
rom[1076] = 12'hfff;
rom[1077] = 12'hfff;
rom[1078] = 12'hfff;
rom[1079] = 12'hfff;
rom[1080] = 12'hfff;
rom[1081] = 12'hfff;
rom[1082] = 12'hfff;
rom[1083] = 12'hfff;
rom[1084] = 12'hfff;
rom[1085] = 12'hfff;
rom[1086] = 12'hfff;
rom[1087] = 12'hfff;
rom[1088] = 12'hfff;
rom[1089] = 12'hfff;
rom[1090] = 12'hfff;
rom[1091] = 12'hfff;
rom[1092] = 12'hfff;
rom[1093] = 12'hfff;
rom[1094] = 12'hfff;
rom[1095] = 12'hfff;
rom[1096] = 12'hfff;
rom[1097] = 12'hfff;
rom[1098] = 12'hfff;
rom[1099] = 12'hfff;
rom[1100] = 12'hfff;
rom[1101] = 12'hfff;
rom[1102] = 12'hfff;
rom[1103] = 12'hfff;
rom[1104] = 12'hfff;
rom[1105] = 12'hfff;
rom[1106] = 12'hfff;
rom[1107] = 12'hfff;
rom[1108] = 12'hfff;
rom[1109] = 12'hfff;
rom[1110] = 12'hfff;
rom[1111] = 12'hfff;
rom[1112] = 12'hfff;
rom[1113] = 12'hfff;
rom[1114] = 12'hfff;
rom[1115] = 12'hfff;
rom[1116] = 12'hfff;
rom[1117] = 12'hfff;
rom[1118] = 12'hfff;
rom[1119] = 12'hfff;
rom[1120] = 12'hfff;
rom[1121] = 12'hfff;
rom[1122] = 12'hfff;
rom[1123] = 12'hfff;
rom[1124] = 12'hfff;
rom[1125] = 12'hfff;
rom[1126] = 12'hfff;
rom[1127] = 12'hfff;
rom[1128] = 12'hfff;
rom[1129] = 12'hfff;
rom[1130] = 12'hfff;
rom[1131] = 12'hfff;
rom[1132] = 12'hfff;
rom[1133] = 12'hfff;
rom[1134] = 12'hfff;
rom[1135] = 12'hfff;
rom[1136] = 12'hfff;
rom[1137] = 12'hfff;
rom[1138] = 12'hfff;
rom[1139] = 12'hfff;
rom[1140] = 12'hfff;
rom[1141] = 12'hfff;
rom[1142] = 12'hfff;
rom[1143] = 12'hfff;
rom[1144] = 12'hfff;
rom[1145] = 12'hfff;
rom[1146] = 12'hfff;
rom[1147] = 12'hfff;
rom[1148] = 12'hfff;
rom[1149] = 12'hfff;
rom[1150] = 12'hfff;
rom[1151] = 12'hfff;
rom[1152] = 12'hfff;
rom[1153] = 12'hfff;
rom[1154] = 12'hfff;
rom[1155] = 12'hfff;
rom[1156] = 12'hfff;
rom[1157] = 12'hfff;
rom[1158] = 12'hfff;
rom[1159] = 12'hfff;
rom[1160] = 12'hfff;
rom[1161] = 12'hfff;
rom[1162] = 12'hfff;
rom[1163] = 12'hfff;
rom[1164] = 12'hfff;
rom[1165] = 12'hfff;
rom[1166] = 12'hfff;
rom[1167] = 12'hfff;
rom[1168] = 12'hfff;
rom[1169] = 12'hfff;
rom[1170] = 12'hfff;
rom[1171] = 12'hfff;
rom[1172] = 12'hfff;
rom[1173] = 12'hfff;
rom[1174] = 12'hfff;
rom[1175] = 12'hfff;
rom[1176] = 12'hfff;
rom[1177] = 12'hfff;
rom[1178] = 12'hfff;
rom[1179] = 12'hfff;
rom[1180] = 12'hfff;
rom[1181] = 12'hfff;
rom[1182] = 12'hfff;
rom[1183] = 12'hfff;
rom[1184] = 12'hfff;
rom[1185] = 12'hfff;
rom[1186] = 12'hfff;
rom[1187] = 12'hfff;
rom[1188] = 12'hfff;
rom[1189] = 12'hfff;
rom[1190] = 12'hfff;
rom[1191] = 12'hfff;
rom[1192] = 12'hfff;
rom[1193] = 12'hfff;
rom[1194] = 12'hfff;
rom[1195] = 12'hfff;
rom[1196] = 12'hfff;
rom[1197] = 12'hfff;
rom[1198] = 12'hfff;
rom[1199] = 12'hfff;
rom[1200] = 12'hfff;
rom[1201] = 12'hfff;
rom[1202] = 12'hfff;
rom[1203] = 12'hfff;
rom[1204] = 12'hfff;
rom[1205] = 12'hfff;
rom[1206] = 12'hfff;
rom[1207] = 12'hfff;
rom[1208] = 12'hfff;
rom[1209] = 12'hfff;
rom[1210] = 12'hfff;
rom[1211] = 12'hfff;
rom[1212] = 12'hfff;
rom[1213] = 12'hfff;
rom[1214] = 12'hfff;
rom[1215] = 12'hfff;
rom[1216] = 12'hfff;
rom[1217] = 12'hfff;
rom[1218] = 12'hfff;
rom[1219] = 12'hfff;
rom[1220] = 12'hfff;
rom[1221] = 12'hfff;
rom[1222] = 12'hfff;
rom[1223] = 12'hfff;
rom[1224] = 12'hfff;
rom[1225] = 12'hfff;
rom[1226] = 12'hfff;
rom[1227] = 12'hfff;
rom[1228] = 12'hfff;
rom[1229] = 12'hfff;
rom[1230] = 12'hfff;
rom[1231] = 12'hfff;
rom[1232] = 12'hfff;
rom[1233] = 12'hfff;
rom[1234] = 12'hfff;
rom[1235] = 12'hfff;
rom[1236] = 12'hfff;
rom[1237] = 12'hfff;
rom[1238] = 12'hfff;
rom[1239] = 12'hfff;
rom[1240] = 12'hfff;
rom[1241] = 12'hfff;
rom[1242] = 12'hfff;
rom[1243] = 12'hfff;
rom[1244] = 12'hfff;
rom[1245] = 12'hfff;
rom[1246] = 12'hfff;
rom[1247] = 12'hfff;
rom[1248] = 12'hfff;
rom[1249] = 12'hfff;
rom[1250] = 12'hfff;
rom[1251] = 12'hfff;
rom[1252] = 12'hfff;
rom[1253] = 12'hfff;
rom[1254] = 12'hfff;
rom[1255] = 12'hfff;
rom[1256] = 12'hfff;
rom[1257] = 12'hfff;
rom[1258] = 12'hfff;
rom[1259] = 12'hfff;
rom[1260] = 12'hfff;
rom[1261] = 12'hfff;
rom[1262] = 12'hfff;
rom[1263] = 12'hfff;
rom[1264] = 12'hfff;
rom[1265] = 12'hfff;
rom[1266] = 12'hfff;
rom[1267] = 12'hfff;
rom[1268] = 12'hfff;
rom[1269] = 12'hfff;
rom[1270] = 12'hfff;
rom[1271] = 12'hfff;
rom[1272] = 12'hfff;
rom[1273] = 12'hfff;
rom[1274] = 12'hfff;
rom[1275] = 12'hfff;
rom[1276] = 12'hfff;
rom[1277] = 12'hfff;
rom[1278] = 12'hfff;
rom[1279] = 12'hfff;
rom[1280] = 12'hfff;
rom[1281] = 12'hfff;
rom[1282] = 12'hfff;
rom[1283] = 12'hfff;
rom[1284] = 12'hfff;
rom[1285] = 12'hfff;
rom[1286] = 12'hfff;
rom[1287] = 12'hfff;
rom[1288] = 12'hfff;
rom[1289] = 12'hfff;
rom[1290] = 12'hfff;
rom[1291] = 12'hfff;
rom[1292] = 12'hfff;
rom[1293] = 12'hfff;
rom[1294] = 12'hfff;
rom[1295] = 12'hfff;
rom[1296] = 12'hfff;
rom[1297] = 12'hfff;
rom[1298] = 12'hfff;
rom[1299] = 12'hfff;
rom[1300] = 12'hfff;
rom[1301] = 12'hfff;
rom[1302] = 12'hfff;
rom[1303] = 12'hfff;
rom[1304] = 12'hfff;
rom[1305] = 12'hfff;
rom[1306] = 12'hfff;
rom[1307] = 12'hfff;
rom[1308] = 12'hfff;
rom[1309] = 12'hfff;
rom[1310] = 12'hfff;
rom[1311] = 12'hfff;
rom[1312] = 12'hfff;
rom[1313] = 12'hfff;
rom[1314] = 12'hfff;
rom[1315] = 12'hfff;
rom[1316] = 12'hfff;
rom[1317] = 12'hfff;
rom[1318] = 12'hfff;
rom[1319] = 12'hfff;
rom[1320] = 12'hfff;
rom[1321] = 12'hfff;
rom[1322] = 12'hfff;
rom[1323] = 12'hfff;
rom[1324] = 12'hfff;
rom[1325] = 12'hfff;
rom[1326] = 12'hfff;
rom[1327] = 12'hfff;
rom[1328] = 12'hfff;
rom[1329] = 12'hfff;
rom[1330] = 12'hfff;
rom[1331] = 12'hfff;
rom[1332] = 12'hfff;
rom[1333] = 12'hfff;
rom[1334] = 12'hfff;
rom[1335] = 12'hfff;
rom[1336] = 12'hfff;
rom[1337] = 12'hfff;
rom[1338] = 12'hfff;
rom[1339] = 12'hfff;
rom[1340] = 12'hfff;
rom[1341] = 12'hfff;
rom[1342] = 12'hfff;
rom[1343] = 12'hfff;
rom[1344] = 12'hfff;
rom[1345] = 12'hfff;
rom[1346] = 12'hfff;
rom[1347] = 12'hfff;
rom[1348] = 12'hfff;
rom[1349] = 12'hfff;
rom[1350] = 12'hfff;
rom[1351] = 12'hfff;
rom[1352] = 12'hfff;
rom[1353] = 12'hfff;
rom[1354] = 12'hfff;
rom[1355] = 12'hfff;
rom[1356] = 12'hfff;
rom[1357] = 12'hfff;
rom[1358] = 12'hfff;
rom[1359] = 12'hfff;
rom[1360] = 12'hfff;
rom[1361] = 12'hfff;
rom[1362] = 12'hfff;
rom[1363] = 12'hfff;
rom[1364] = 12'hfff;
rom[1365] = 12'hfff;
rom[1366] = 12'hfff;
rom[1367] = 12'hfff;
rom[1368] = 12'hfff;
rom[1369] = 12'hfff;
rom[1370] = 12'hfff;
rom[1371] = 12'hfff;
rom[1372] = 12'hfff;
rom[1373] = 12'hfff;
rom[1374] = 12'hfff;
rom[1375] = 12'hfff;
rom[1376] = 12'hfff;
rom[1377] = 12'hfff;
rom[1378] = 12'hfff;
rom[1379] = 12'hfff;
rom[1380] = 12'hfff;
rom[1381] = 12'hfff;
rom[1382] = 12'hfff;
rom[1383] = 12'hfff;
rom[1384] = 12'hfff;
rom[1385] = 12'hfff;
rom[1386] = 12'hfff;
rom[1387] = 12'hfff;
rom[1388] = 12'hfff;
rom[1389] = 12'hfff;
rom[1390] = 12'hfff;
rom[1391] = 12'hfff;
rom[1392] = 12'hfff;
rom[1393] = 12'hfff;
rom[1394] = 12'hfff;
rom[1395] = 12'hfff;
rom[1396] = 12'hfff;
rom[1397] = 12'hfff;
rom[1398] = 12'hfff;
rom[1399] = 12'hfff;
rom[1400] = 12'hfff;
rom[1401] = 12'hfff;
rom[1402] = 12'hfff;
rom[1403] = 12'hfff;
rom[1404] = 12'hfff;
rom[1405] = 12'hfff;
rom[1406] = 12'hfff;
rom[1407] = 12'hfff;
rom[1408] = 12'hfff;
rom[1409] = 12'hfff;
rom[1410] = 12'hfff;
rom[1411] = 12'hfff;
rom[1412] = 12'hfff;
rom[1413] = 12'hfff;
rom[1414] = 12'hfff;
rom[1415] = 12'hfff;
rom[1416] = 12'hfff;
rom[1417] = 12'hfff;
rom[1418] = 12'hfff;
rom[1419] = 12'hfff;
rom[1420] = 12'hfff;
rom[1421] = 12'hfff;
rom[1422] = 12'hfff;
rom[1423] = 12'hfff;
rom[1424] = 12'hfff;
rom[1425] = 12'hfff;
rom[1426] = 12'hfff;
rom[1427] = 12'hfff;
rom[1428] = 12'hfff;
rom[1429] = 12'hfff;
rom[1430] = 12'hfff;
rom[1431] = 12'hfff;
rom[1432] = 12'hfff;
rom[1433] = 12'hfff;
rom[1434] = 12'hfff;
rom[1435] = 12'hfff;
rom[1436] = 12'hfff;
rom[1437] = 12'hfff;
rom[1438] = 12'hfff;
rom[1439] = 12'hfff;
rom[1440] = 12'hfff;
rom[1441] = 12'hfff;
rom[1442] = 12'hfff;
rom[1443] = 12'hfff;
rom[1444] = 12'hfff;
rom[1445] = 12'hfff;
rom[1446] = 12'hfff;
rom[1447] = 12'hfff;
rom[1448] = 12'hfff;
rom[1449] = 12'hfff;
rom[1450] = 12'hfff;
rom[1451] = 12'hfff;
rom[1452] = 12'hfff;
rom[1453] = 12'hfff;
rom[1454] = 12'hfff;
rom[1455] = 12'hfff;
rom[1456] = 12'hfff;
rom[1457] = 12'hfff;
rom[1458] = 12'hfff;
rom[1459] = 12'hfff;
rom[1460] = 12'hfff;
rom[1461] = 12'hfff;
rom[1462] = 12'hfff;
rom[1463] = 12'hfff;
rom[1464] = 12'hfff;
rom[1465] = 12'hfff;
rom[1466] = 12'hfff;
rom[1467] = 12'hfff;
rom[1468] = 12'hfff;
rom[1469] = 12'hfff;
rom[1470] = 12'hfff;
rom[1471] = 12'hfff;
rom[1472] = 12'hfff;
rom[1473] = 12'hfff;
rom[1474] = 12'hfff;
rom[1475] = 12'hfff;
rom[1476] = 12'hfff;
rom[1477] = 12'hfff;
rom[1478] = 12'hfff;
rom[1479] = 12'hfff;
rom[1480] = 12'hfff;
rom[1481] = 12'hfff;
rom[1482] = 12'hfff;
rom[1483] = 12'hfff;
rom[1484] = 12'hfff;
rom[1485] = 12'hfff;
rom[1486] = 12'hfff;
rom[1487] = 12'hfff;
rom[1488] = 12'hfff;
rom[1489] = 12'hfff;
rom[1490] = 12'hfff;
rom[1491] = 12'hfff;
rom[1492] = 12'hfff;
rom[1493] = 12'hfff;
rom[1494] = 12'hfff;
rom[1495] = 12'hfff;
rom[1496] = 12'hfff;
rom[1497] = 12'hfff;
rom[1498] = 12'hfff;
rom[1499] = 12'hfff;
rom[1500] = 12'hfff;
rom[1501] = 12'hfff;
rom[1502] = 12'hfff;
rom[1503] = 12'hfff;
rom[1504] = 12'hfff;
rom[1505] = 12'hfff;
rom[1506] = 12'hfff;
rom[1507] = 12'hfff;
rom[1508] = 12'hfff;
rom[1509] = 12'hfff;
rom[1510] = 12'hfff;
rom[1511] = 12'hfff;
rom[1512] = 12'hfff;
rom[1513] = 12'hfff;
rom[1514] = 12'hfff;
rom[1515] = 12'hfff;
rom[1516] = 12'hfff;
rom[1517] = 12'hfff;
rom[1518] = 12'hfff;
rom[1519] = 12'hfff;
rom[1520] = 12'hfff;
rom[1521] = 12'hfff;
rom[1522] = 12'hfff;
rom[1523] = 12'hfff;
rom[1524] = 12'hfff;
rom[1525] = 12'hfff;
rom[1526] = 12'hfff;
rom[1527] = 12'hfff;
rom[1528] = 12'hfff;
rom[1529] = 12'hfff;
rom[1530] = 12'hfff;
rom[1531] = 12'hfff;
rom[1532] = 12'hfff;
rom[1533] = 12'hfff;
rom[1534] = 12'hfff;
rom[1535] = 12'hfff;
rom[1536] = 12'hfff;
rom[1537] = 12'hfff;
rom[1538] = 12'hfff;
rom[1539] = 12'hfff;
rom[1540] = 12'hfff;
rom[1541] = 12'hfff;
rom[1542] = 12'hfff;
rom[1543] = 12'hfff;
rom[1544] = 12'hfff;
rom[1545] = 12'hfff;
rom[1546] = 12'hfff;
rom[1547] = 12'hfff;
rom[1548] = 12'hfff;
rom[1549] = 12'hfff;
rom[1550] = 12'hfff;
rom[1551] = 12'hfff;
rom[1552] = 12'hfff;
rom[1553] = 12'hfff;
rom[1554] = 12'hfff;
rom[1555] = 12'hfff;
rom[1556] = 12'hfff;
rom[1557] = 12'hfff;
rom[1558] = 12'hfff;
rom[1559] = 12'hfff;
rom[1560] = 12'hfff;
rom[1561] = 12'hfff;
rom[1562] = 12'hfff;
rom[1563] = 12'hfff;
rom[1564] = 12'hfff;
rom[1565] = 12'hfff;
rom[1566] = 12'hfff;
rom[1567] = 12'hfff;
rom[1568] = 12'hfff;
rom[1569] = 12'hfff;
rom[1570] = 12'hfff;
rom[1571] = 12'hfff;
rom[1572] = 12'hfff;
rom[1573] = 12'hfff;
rom[1574] = 12'hfff;
rom[1575] = 12'hfff;
rom[1576] = 12'hfff;
rom[1577] = 12'hfff;
rom[1578] = 12'hfff;
rom[1579] = 12'hfff;
rom[1580] = 12'hfff;
rom[1581] = 12'hfff;
rom[1582] = 12'hfff;
rom[1583] = 12'hfff;
rom[1584] = 12'hfff;
rom[1585] = 12'hfff;
rom[1586] = 12'hfff;
rom[1587] = 12'hfff;
rom[1588] = 12'hfff;
rom[1589] = 12'hfff;
rom[1590] = 12'hfff;
rom[1591] = 12'hfff;
rom[1592] = 12'hfff;
rom[1593] = 12'hfff;
rom[1594] = 12'hfff;
rom[1595] = 12'hfff;
rom[1596] = 12'hfff;
rom[1597] = 12'hfff;
rom[1598] = 12'hfff;
rom[1599] = 12'hfff;
rom[1600] = 12'hfff;
rom[1601] = 12'hfff;
rom[1602] = 12'hfff;
rom[1603] = 12'hfff;
rom[1604] = 12'hfff;
rom[1605] = 12'hfff;
rom[1606] = 12'hfff;
rom[1607] = 12'hfff;
rom[1608] = 12'hfff;
rom[1609] = 12'hfff;
rom[1610] = 12'hfff;
rom[1611] = 12'hfff;
rom[1612] = 12'hfff;
rom[1613] = 12'hfff;
rom[1614] = 12'hfff;
rom[1615] = 12'hfff;
rom[1616] = 12'hfff;
rom[1617] = 12'hfff;
rom[1618] = 12'hfff;
rom[1619] = 12'hfff;
rom[1620] = 12'hfff;
rom[1621] = 12'hfff;
rom[1622] = 12'hfff;
rom[1623] = 12'hfff;
rom[1624] = 12'hfff;
rom[1625] = 12'hfff;
rom[1626] = 12'hfff;
rom[1627] = 12'hfff;
rom[1628] = 12'hfff;
rom[1629] = 12'hfff;
rom[1630] = 12'hfff;
rom[1631] = 12'hfff;
rom[1632] = 12'hfff;
rom[1633] = 12'hfff;
rom[1634] = 12'hfff;
rom[1635] = 12'hfff;
rom[1636] = 12'hfff;
rom[1637] = 12'hfff;
rom[1638] = 12'hfff;
rom[1639] = 12'hfff;
rom[1640] = 12'hfff;
rom[1641] = 12'hfff;
rom[1642] = 12'hfff;
rom[1643] = 12'hfff;
rom[1644] = 12'hfff;
rom[1645] = 12'hfff;
rom[1646] = 12'hfff;
rom[1647] = 12'hfff;
rom[1648] = 12'hfff;
rom[1649] = 12'hfff;
rom[1650] = 12'hfff;
rom[1651] = 12'hfff;
rom[1652] = 12'hfff;
rom[1653] = 12'hfff;
rom[1654] = 12'hfff;
rom[1655] = 12'hfff;
rom[1656] = 12'hfff;
rom[1657] = 12'hfff;
rom[1658] = 12'hfff;
rom[1659] = 12'hfff;
rom[1660] = 12'hfff;
rom[1661] = 12'hfff;
rom[1662] = 12'hfff;
rom[1663] = 12'hfff;
rom[1664] = 12'hfff;
rom[1665] = 12'hfff;
rom[1666] = 12'hfff;
rom[1667] = 12'hfff;
rom[1668] = 12'hfff;
rom[1669] = 12'hfff;
rom[1670] = 12'hfff;
rom[1671] = 12'hfff;
rom[1672] = 12'hfff;
rom[1673] = 12'hfff;
rom[1674] = 12'hfff;
rom[1675] = 12'hfff;
rom[1676] = 12'hfff;
rom[1677] = 12'hfff;
rom[1678] = 12'hfff;
rom[1679] = 12'hfff;
rom[1680] = 12'hfff;
rom[1681] = 12'hfff;
rom[1682] = 12'hfff;
rom[1683] = 12'hfff;
rom[1684] = 12'hfff;
rom[1685] = 12'hfff;
rom[1686] = 12'hfff;
rom[1687] = 12'hfff;
rom[1688] = 12'hfff;
rom[1689] = 12'hfff;
rom[1690] = 12'hfff;
rom[1691] = 12'hfff;
rom[1692] = 12'hfff;
rom[1693] = 12'hfff;
rom[1694] = 12'hfff;
rom[1695] = 12'hfff;
rom[1696] = 12'hfff;
rom[1697] = 12'hfff;
rom[1698] = 12'hfff;
rom[1699] = 12'hfff;
rom[1700] = 12'hfff;
rom[1701] = 12'hfff;
rom[1702] = 12'hfff;
rom[1703] = 12'hfff;
rom[1704] = 12'hfff;
rom[1705] = 12'hfff;
rom[1706] = 12'hfff;
rom[1707] = 12'hfff;
rom[1708] = 12'hfff;
rom[1709] = 12'hfff;
rom[1710] = 12'hfff;
rom[1711] = 12'hfff;
rom[1712] = 12'hfff;
rom[1713] = 12'hfff;
rom[1714] = 12'hfff;
rom[1715] = 12'hfff;
rom[1716] = 12'hfff;
rom[1717] = 12'hfff;
rom[1718] = 12'hfff;
rom[1719] = 12'hfff;
rom[1720] = 12'hfff;
rom[1721] = 12'hfff;
rom[1722] = 12'hfff;
rom[1723] = 12'hfff;
rom[1724] = 12'hfff;
rom[1725] = 12'hfff;
rom[1726] = 12'hfff;
rom[1727] = 12'hfff;
rom[1728] = 12'hfff;
rom[1729] = 12'hfff;
rom[1730] = 12'hfff;
rom[1731] = 12'hfff;
rom[1732] = 12'hfff;
rom[1733] = 12'hfff;
rom[1734] = 12'hfff;
rom[1735] = 12'hfff;
rom[1736] = 12'hfff;
rom[1737] = 12'hfff;
rom[1738] = 12'hfff;
rom[1739] = 12'hfff;
rom[1740] = 12'hfff;
rom[1741] = 12'hfff;
rom[1742] = 12'hfff;
rom[1743] = 12'hfff;
rom[1744] = 12'hfff;
rom[1745] = 12'hfff;
rom[1746] = 12'hfff;
rom[1747] = 12'hfff;
rom[1748] = 12'hfff;
rom[1749] = 12'hfff;
rom[1750] = 12'hfff;
rom[1751] = 12'hfff;
rom[1752] = 12'hfff;
rom[1753] = 12'hfff;
rom[1754] = 12'hfff;
rom[1755] = 12'hfff;
rom[1756] = 12'hfff;
rom[1757] = 12'hfff;
rom[1758] = 12'hfff;
rom[1759] = 12'hfff;
rom[1760] = 12'hfff;
rom[1761] = 12'hfff;
rom[1762] = 12'hfff;
rom[1763] = 12'hfff;
rom[1764] = 12'hfff;
rom[1765] = 12'hfff;
rom[1766] = 12'hfff;
rom[1767] = 12'hfff;
rom[1768] = 12'hfff;
rom[1769] = 12'hfff;
rom[1770] = 12'hfff;
rom[1771] = 12'hfff;
rom[1772] = 12'hfff;
rom[1773] = 12'hfff;
rom[1774] = 12'hfff;
rom[1775] = 12'hfff;
rom[1776] = 12'hfff;
rom[1777] = 12'hfff;
rom[1778] = 12'hfff;
rom[1779] = 12'hfff;
rom[1780] = 12'hfff;
rom[1781] = 12'hfff;
rom[1782] = 12'hfff;
rom[1783] = 12'hfff;
rom[1784] = 12'hfff;
rom[1785] = 12'hfff;
rom[1786] = 12'hfff;
rom[1787] = 12'hfff;
rom[1788] = 12'hfff;
rom[1789] = 12'hfff;
rom[1790] = 12'hfff;
rom[1791] = 12'hfff;
rom[1792] = 12'hfff;
rom[1793] = 12'hfff;
rom[1794] = 12'hfff;
rom[1795] = 12'hfff;
rom[1796] = 12'hfff;
rom[1797] = 12'hfff;
rom[1798] = 12'hfff;
rom[1799] = 12'hfff;
rom[1800] = 12'hfff;
rom[1801] = 12'hfff;
rom[1802] = 12'hfff;
rom[1803] = 12'hfff;
rom[1804] = 12'hfff;
rom[1805] = 12'hfff;
rom[1806] = 12'hfff;
rom[1807] = 12'hfff;
rom[1808] = 12'hfff;
rom[1809] = 12'hfff;
rom[1810] = 12'hfff;
rom[1811] = 12'hfff;
rom[1812] = 12'hfff;
rom[1813] = 12'hfff;
rom[1814] = 12'hfff;
rom[1815] = 12'hfff;
rom[1816] = 12'hfff;
rom[1817] = 12'hfff;
rom[1818] = 12'hfff;
rom[1819] = 12'hfff;
rom[1820] = 12'hfff;
rom[1821] = 12'hfff;
rom[1822] = 12'hfff;
rom[1823] = 12'hfff;
rom[1824] = 12'hfff;
rom[1825] = 12'hfff;
rom[1826] = 12'hfff;
rom[1827] = 12'hfff;
rom[1828] = 12'hfff;
rom[1829] = 12'hfff;
rom[1830] = 12'hfff;
rom[1831] = 12'hfff;
rom[1832] = 12'hfff;
rom[1833] = 12'hfff;
rom[1834] = 12'hfff;
rom[1835] = 12'hfff;
rom[1836] = 12'hfff;
rom[1837] = 12'hfff;
rom[1838] = 12'hfff;
rom[1839] = 12'hfff;
rom[1840] = 12'hfff;
rom[1841] = 12'hfff;
rom[1842] = 12'hfff;
rom[1843] = 12'hfff;
rom[1844] = 12'hfff;
rom[1845] = 12'hfff;
rom[1846] = 12'hfff;
rom[1847] = 12'hfff;
rom[1848] = 12'hfff;
rom[1849] = 12'hfff;
rom[1850] = 12'hfff;
rom[1851] = 12'hfff;
rom[1852] = 12'hfff;
rom[1853] = 12'hfff;
rom[1854] = 12'hfff;
rom[1855] = 12'hfff;
rom[1856] = 12'hfff;
rom[1857] = 12'hfff;
rom[1858] = 12'hfff;
rom[1859] = 12'hfff;
rom[1860] = 12'hfff;
rom[1861] = 12'hfff;
rom[1862] = 12'hfff;
rom[1863] = 12'hfff;
rom[1864] = 12'hfff;
rom[1865] = 12'hfff;
rom[1866] = 12'hfff;
rom[1867] = 12'hfff;
rom[1868] = 12'hfff;
rom[1869] = 12'hfff;
rom[1870] = 12'hfff;
rom[1871] = 12'hfff;
rom[1872] = 12'hfff;
rom[1873] = 12'hfff;
rom[1874] = 12'hfff;
rom[1875] = 12'hfff;
rom[1876] = 12'hfff;
rom[1877] = 12'hfff;
rom[1878] = 12'hfff;
rom[1879] = 12'hfff;
rom[1880] = 12'hfff;
rom[1881] = 12'hfff;
rom[1882] = 12'hfff;
rom[1883] = 12'hfff;
rom[1884] = 12'hfff;
rom[1885] = 12'hfff;
rom[1886] = 12'hfff;
rom[1887] = 12'hfff;
rom[1888] = 12'hfff;
rom[1889] = 12'hfff;
rom[1890] = 12'hfff;
rom[1891] = 12'hfff;
rom[1892] = 12'hfff;
rom[1893] = 12'hfff;
rom[1894] = 12'hfff;
rom[1895] = 12'hfff;
rom[1896] = 12'hfff;
rom[1897] = 12'hfff;
rom[1898] = 12'hfff;
rom[1899] = 12'hfff;
rom[1900] = 12'hfff;
rom[1901] = 12'hfff;
rom[1902] = 12'hfff;
rom[1903] = 12'hfff;
rom[1904] = 12'hfff;
rom[1905] = 12'hfff;
rom[1906] = 12'hfff;
rom[1907] = 12'hfff;
rom[1908] = 12'hfff;
rom[1909] = 12'hfff;
rom[1910] = 12'hfff;
rom[1911] = 12'hfff;
rom[1912] = 12'hfff;
rom[1913] = 12'hfff;
rom[1914] = 12'hfff;
rom[1915] = 12'hfff;
rom[1916] = 12'hfff;
rom[1917] = 12'hfff;
rom[1918] = 12'hfff;
rom[1919] = 12'hfff;
rom[1920] = 12'hfff;
rom[1921] = 12'hfff;
rom[1922] = 12'hfff;
rom[1923] = 12'hfff;
rom[1924] = 12'hfff;
rom[1925] = 12'hfff;
rom[1926] = 12'hfff;
rom[1927] = 12'hfff;
rom[1928] = 12'hfff;
rom[1929] = 12'hfff;
rom[1930] = 12'hfff;
rom[1931] = 12'hfff;
rom[1932] = 12'hfff;
rom[1933] = 12'hfff;
rom[1934] = 12'hfff;
rom[1935] = 12'hfff;
rom[1936] = 12'hfff;
rom[1937] = 12'hfff;
rom[1938] = 12'hfff;
rom[1939] = 12'hfff;
rom[1940] = 12'hfff;
rom[1941] = 12'hfff;
rom[1942] = 12'hfff;
rom[1943] = 12'hfff;
rom[1944] = 12'hfff;
rom[1945] = 12'hfff;
rom[1946] = 12'hfff;
rom[1947] = 12'hfff;
rom[1948] = 12'hfff;
rom[1949] = 12'hfff;
rom[1950] = 12'hfff;
rom[1951] = 12'hfff;
rom[1952] = 12'hfff;
rom[1953] = 12'hfff;
rom[1954] = 12'hfff;
rom[1955] = 12'hfff;
rom[1956] = 12'hfff;
rom[1957] = 12'hfff;
rom[1958] = 12'hfff;
rom[1959] = 12'hfff;
rom[1960] = 12'hfff;
rom[1961] = 12'hfff;
rom[1962] = 12'hfff;
rom[1963] = 12'hfff;
rom[1964] = 12'hfff;
rom[1965] = 12'hfff;
rom[1966] = 12'hfff;
rom[1967] = 12'hfff;
rom[1968] = 12'hfff;
rom[1969] = 12'hfff;
rom[1970] = 12'hfff;
rom[1971] = 12'hfff;
rom[1972] = 12'hfff;
rom[1973] = 12'hfff;
rom[1974] = 12'hfff;
rom[1975] = 12'hfff;
rom[1976] = 12'hfff;
rom[1977] = 12'hfff;
rom[1978] = 12'hfff;
rom[1979] = 12'hfff;
rom[1980] = 12'hfff;
rom[1981] = 12'hfff;
rom[1982] = 12'hfff;
rom[1983] = 12'hfff;
rom[1984] = 12'hfff;
rom[1985] = 12'hfff;
rom[1986] = 12'hfff;
rom[1987] = 12'hfff;
rom[1988] = 12'hfff;
rom[1989] = 12'hfff;
rom[1990] = 12'hfff;
rom[1991] = 12'hfff;
rom[1992] = 12'hfff;
rom[1993] = 12'hfff;
rom[1994] = 12'hfff;
rom[1995] = 12'hfff;
rom[1996] = 12'hfff;
rom[1997] = 12'hfff;
rom[1998] = 12'hfff;
rom[1999] = 12'hfff;
rom[2000] = 12'hfff;
rom[2001] = 12'hfff;
rom[2002] = 12'hfff;
rom[2003] = 12'hfff;
rom[2004] = 12'hfff;
rom[2005] = 12'hfff;
rom[2006] = 12'hfff;
rom[2007] = 12'hfff;
rom[2008] = 12'hfff;
rom[2009] = 12'hfff;
rom[2010] = 12'hfff;
rom[2011] = 12'hfff;
rom[2012] = 12'hfff;
rom[2013] = 12'hfff;
rom[2014] = 12'hfff;
rom[2015] = 12'hfff;
rom[2016] = 12'hfff;
rom[2017] = 12'hfff;
rom[2018] = 12'hfff;
rom[2019] = 12'hfff;
rom[2020] = 12'hfff;
rom[2021] = 12'hfff;
rom[2022] = 12'hfff;
rom[2023] = 12'hfff;
rom[2024] = 12'hfff;
rom[2025] = 12'hfff;
rom[2026] = 12'hfff;
rom[2027] = 12'hfff;
rom[2028] = 12'hfff;
rom[2029] = 12'hfff;
rom[2030] = 12'hfff;
rom[2031] = 12'hfff;
rom[2032] = 12'hfff;
rom[2033] = 12'hfff;
rom[2034] = 12'hfff;
rom[2035] = 12'hfff;
rom[2036] = 12'hfff;
rom[2037] = 12'hfff;
rom[2038] = 12'hfff;
rom[2039] = 12'hfff;
rom[2040] = 12'hfff;
rom[2041] = 12'hfff;
rom[2042] = 12'hfff;
rom[2043] = 12'hfff;
rom[2044] = 12'hfff;
rom[2045] = 12'hfff;
rom[2046] = 12'hfff;
rom[2047] = 12'hfff;
rom[2048] = 12'hfff;
rom[2049] = 12'hfff;
rom[2050] = 12'hfff;
rom[2051] = 12'hfff;
rom[2052] = 12'hfff;
rom[2053] = 12'hfff;
rom[2054] = 12'hfff;
rom[2055] = 12'hfff;
rom[2056] = 12'hfff;
rom[2057] = 12'hfff;
rom[2058] = 12'hfff;
rom[2059] = 12'hfff;
rom[2060] = 12'hfff;
rom[2061] = 12'hfff;
rom[2062] = 12'hfff;
rom[2063] = 12'hfff;
rom[2064] = 12'hfff;
rom[2065] = 12'hfff;
rom[2066] = 12'hfff;
rom[2067] = 12'hfff;
rom[2068] = 12'hfff;
rom[2069] = 12'hfff;
rom[2070] = 12'hfff;
rom[2071] = 12'hfff;
rom[2072] = 12'hfff;
rom[2073] = 12'hfff;
rom[2074] = 12'hfff;
rom[2075] = 12'hfff;
rom[2076] = 12'hfff;
rom[2077] = 12'hfff;
rom[2078] = 12'hfff;
rom[2079] = 12'hfff;
rom[2080] = 12'hfff;
rom[2081] = 12'hfff;
rom[2082] = 12'hfff;
rom[2083] = 12'hfff;
rom[2084] = 12'hfff;
rom[2085] = 12'hfff;
rom[2086] = 12'hfff;
rom[2087] = 12'hfff;
rom[2088] = 12'hfff;
rom[2089] = 12'hfff;
rom[2090] = 12'hfff;
rom[2091] = 12'hfff;
rom[2092] = 12'hfff;
rom[2093] = 12'hfff;
rom[2094] = 12'hfff;
rom[2095] = 12'hfff;
rom[2096] = 12'hfff;
rom[2097] = 12'hfff;
rom[2098] = 12'hfff;
rom[2099] = 12'hfff;
rom[2100] = 12'hfff;
rom[2101] = 12'hfff;
rom[2102] = 12'hfff;
rom[2103] = 12'hfff;
rom[2104] = 12'hfff;
rom[2105] = 12'hfff;
rom[2106] = 12'hfff;
rom[2107] = 12'hfff;
rom[2108] = 12'hfff;
rom[2109] = 12'hfff;
rom[2110] = 12'hfff;
rom[2111] = 12'hfff;
rom[2112] = 12'hfff;
rom[2113] = 12'hfff;
rom[2114] = 12'hfff;
rom[2115] = 12'hfff;
rom[2116] = 12'hfff;
rom[2117] = 12'hfff;
rom[2118] = 12'hfff;
rom[2119] = 12'hfff;
rom[2120] = 12'hfff;
rom[2121] = 12'hfff;
rom[2122] = 12'hfff;
rom[2123] = 12'hfff;
rom[2124] = 12'hfff;
rom[2125] = 12'hfff;
rom[2126] = 12'hfff;
rom[2127] = 12'hfff;
rom[2128] = 12'hfff;
rom[2129] = 12'hfff;
rom[2130] = 12'hfff;
rom[2131] = 12'hfff;
rom[2132] = 12'hfff;
rom[2133] = 12'hfff;
rom[2134] = 12'hfff;
rom[2135] = 12'hfff;
rom[2136] = 12'hfff;
rom[2137] = 12'hfff;
rom[2138] = 12'hfff;
rom[2139] = 12'hfff;
rom[2140] = 12'hfff;
rom[2141] = 12'hfff;
rom[2142] = 12'hfff;
rom[2143] = 12'hfff;
rom[2144] = 12'hfff;
rom[2145] = 12'hfff;
rom[2146] = 12'hfff;
rom[2147] = 12'hfff;
rom[2148] = 12'hfff;
rom[2149] = 12'hfff;
rom[2150] = 12'hfff;
rom[2151] = 12'hfff;
rom[2152] = 12'hfff;
rom[2153] = 12'hfff;
rom[2154] = 12'hfff;
rom[2155] = 12'hfff;
rom[2156] = 12'hfff;
rom[2157] = 12'hfff;
rom[2158] = 12'hfff;
rom[2159] = 12'hfff;
rom[2160] = 12'hfff;
rom[2161] = 12'hfff;
rom[2162] = 12'hfff;
rom[2163] = 12'hfff;
rom[2164] = 12'hfff;
rom[2165] = 12'hfff;
rom[2166] = 12'hfff;
rom[2167] = 12'hfff;
rom[2168] = 12'hfff;
rom[2169] = 12'hfff;
rom[2170] = 12'hfff;
rom[2171] = 12'hfff;
rom[2172] = 12'hfff;
rom[2173] = 12'hfff;
rom[2174] = 12'hfff;
rom[2175] = 12'hfff;
rom[2176] = 12'hfff;
rom[2177] = 12'hfff;
rom[2178] = 12'hfff;
rom[2179] = 12'hfff;
rom[2180] = 12'hfff;
rom[2181] = 12'hfff;
rom[2182] = 12'hfff;
rom[2183] = 12'hfff;
rom[2184] = 12'hfff;
rom[2185] = 12'hfff;
rom[2186] = 12'hfff;
rom[2187] = 12'hfff;
rom[2188] = 12'hfff;
rom[2189] = 12'hfff;
rom[2190] = 12'hfff;
rom[2191] = 12'hfff;
rom[2192] = 12'hfff;
rom[2193] = 12'hfff;
rom[2194] = 12'hfff;
rom[2195] = 12'hfff;
rom[2196] = 12'hfff;
rom[2197] = 12'hfff;
rom[2198] = 12'hfff;
rom[2199] = 12'hfff;
rom[2200] = 12'hfff;
rom[2201] = 12'hfff;
rom[2202] = 12'hfff;
rom[2203] = 12'hfff;
rom[2204] = 12'hfff;
rom[2205] = 12'hfff;
rom[2206] = 12'hfff;
rom[2207] = 12'hfff;
rom[2208] = 12'hfff;
rom[2209] = 12'hfff;
rom[2210] = 12'hfff;
rom[2211] = 12'hfff;
rom[2212] = 12'hfff;
rom[2213] = 12'hfff;
rom[2214] = 12'hfff;
rom[2215] = 12'hfff;
rom[2216] = 12'hfff;
rom[2217] = 12'hfff;
rom[2218] = 12'hfff;
rom[2219] = 12'hfff;
rom[2220] = 12'hfff;
rom[2221] = 12'hfff;
rom[2222] = 12'hfff;
rom[2223] = 12'hfff;
rom[2224] = 12'hfff;
rom[2225] = 12'hfff;
rom[2226] = 12'hfff;
rom[2227] = 12'hfff;
rom[2228] = 12'hfff;
rom[2229] = 12'hfff;
rom[2230] = 12'hfff;
rom[2231] = 12'hfff;
rom[2232] = 12'hfff;
rom[2233] = 12'hfff;
rom[2234] = 12'hfff;
rom[2235] = 12'hfff;
rom[2236] = 12'hfff;
rom[2237] = 12'hfff;
rom[2238] = 12'hfff;
rom[2239] = 12'hfff;
rom[2240] = 12'hfff;
rom[2241] = 12'hfff;
rom[2242] = 12'hfff;
rom[2243] = 12'hfff;
rom[2244] = 12'hfff;
rom[2245] = 12'hfff;
rom[2246] = 12'hfff;
rom[2247] = 12'hfff;
rom[2248] = 12'hfff;
rom[2249] = 12'hfff;
rom[2250] = 12'hfff;
rom[2251] = 12'hfff;
rom[2252] = 12'hfff;
rom[2253] = 12'hfff;
rom[2254] = 12'hfff;
rom[2255] = 12'hfff;
rom[2256] = 12'hfff;
rom[2257] = 12'hfff;
rom[2258] = 12'hfff;
rom[2259] = 12'hfff;
rom[2260] = 12'hfff;
rom[2261] = 12'hfff;
rom[2262] = 12'hfff;
rom[2263] = 12'hfff;
rom[2264] = 12'hfff;
rom[2265] = 12'hfff;
rom[2266] = 12'hfff;
rom[2267] = 12'hfff;
rom[2268] = 12'hfff;
rom[2269] = 12'hfff;
rom[2270] = 12'hfff;
rom[2271] = 12'hfff;
rom[2272] = 12'hfff;
rom[2273] = 12'hfff;
rom[2274] = 12'hfff;
rom[2275] = 12'hfff;
rom[2276] = 12'hfff;
rom[2277] = 12'hfff;
rom[2278] = 12'hfff;
rom[2279] = 12'hfff;
rom[2280] = 12'hfff;
rom[2281] = 12'hfff;
rom[2282] = 12'hfff;
rom[2283] = 12'hfff;
rom[2284] = 12'hfff;
rom[2285] = 12'hfff;
rom[2286] = 12'hfff;
rom[2287] = 12'hfff;
rom[2288] = 12'hfff;
rom[2289] = 12'hfff;
rom[2290] = 12'hfff;
rom[2291] = 12'hfff;
rom[2292] = 12'hfff;
rom[2293] = 12'hfff;
rom[2294] = 12'hfff;
rom[2295] = 12'hfff;
rom[2296] = 12'hfff;
rom[2297] = 12'hfff;
rom[2298] = 12'hfff;
rom[2299] = 12'hfff;
rom[2300] = 12'hfff;
rom[2301] = 12'hfff;
rom[2302] = 12'hfff;
rom[2303] = 12'hfff;
rom[2304] = 12'hfff;
rom[2305] = 12'hfff;
rom[2306] = 12'hfff;
rom[2307] = 12'hfff;
rom[2308] = 12'hfff;
rom[2309] = 12'hfff;
rom[2310] = 12'hfff;
rom[2311] = 12'hfff;
rom[2312] = 12'hfff;
rom[2313] = 12'hfff;
rom[2314] = 12'hfff;
rom[2315] = 12'hfff;
rom[2316] = 12'hfff;
rom[2317] = 12'hfff;
rom[2318] = 12'hfff;
rom[2319] = 12'hfff;
rom[2320] = 12'hfff;
rom[2321] = 12'hfff;
rom[2322] = 12'hfff;
rom[2323] = 12'hfff;
rom[2324] = 12'hfff;
rom[2325] = 12'hfff;
rom[2326] = 12'hfff;
rom[2327] = 12'hfff;
rom[2328] = 12'hfff;
rom[2329] = 12'hfff;
rom[2330] = 12'hfff;
rom[2331] = 12'hfff;
rom[2332] = 12'hfff;
rom[2333] = 12'hfff;
rom[2334] = 12'hfff;
rom[2335] = 12'hfff;
rom[2336] = 12'hfff;
rom[2337] = 12'hfff;
rom[2338] = 12'hfff;
rom[2339] = 12'hfff;
rom[2340] = 12'hfff;
rom[2341] = 12'hfff;
rom[2342] = 12'hfff;
rom[2343] = 12'hfff;
rom[2344] = 12'hfff;
rom[2345] = 12'hfff;
rom[2346] = 12'hfff;
rom[2347] = 12'hfff;
rom[2348] = 12'hfff;
rom[2349] = 12'hfff;
rom[2350] = 12'hfff;
rom[2351] = 12'hfff;
rom[2352] = 12'hfff;
rom[2353] = 12'hfff;
rom[2354] = 12'hfff;
rom[2355] = 12'hfff;
rom[2356] = 12'hfff;
rom[2357] = 12'hfff;
rom[2358] = 12'hfff;
rom[2359] = 12'hfff;
rom[2360] = 12'hfff;
rom[2361] = 12'hfff;
rom[2362] = 12'hfff;
rom[2363] = 12'hfff;
rom[2364] = 12'hfff;
rom[2365] = 12'hfff;
rom[2366] = 12'hfff;
rom[2367] = 12'hfff;
rom[2368] = 12'hfff;
rom[2369] = 12'hfff;
rom[2370] = 12'hfff;
rom[2371] = 12'hfff;
rom[2372] = 12'hfff;
rom[2373] = 12'hfff;
rom[2374] = 12'hfff;
rom[2375] = 12'hfff;
rom[2376] = 12'hfff;
rom[2377] = 12'hfff;
rom[2378] = 12'hfff;
rom[2379] = 12'hfff;
rom[2380] = 12'hfff;
rom[2381] = 12'hfff;
rom[2382] = 12'hfff;
rom[2383] = 12'hfff;
rom[2384] = 12'hfff;
rom[2385] = 12'hfff;
rom[2386] = 12'hfff;
rom[2387] = 12'hfff;
rom[2388] = 12'hfff;
rom[2389] = 12'hfff;
rom[2390] = 12'hfff;
rom[2391] = 12'hfff;
rom[2392] = 12'hfff;
rom[2393] = 12'hfff;
rom[2394] = 12'hfff;
rom[2395] = 12'hfff;
rom[2396] = 12'hfff;
rom[2397] = 12'hfff;
rom[2398] = 12'hfff;
rom[2399] = 12'hfff;
rom[2400] = 12'hfff;
rom[2401] = 12'hfff;
rom[2402] = 12'hfff;
rom[2403] = 12'hfff;
rom[2404] = 12'hfff;
rom[2405] = 12'hfff;
rom[2406] = 12'hfff;
rom[2407] = 12'hfff;
rom[2408] = 12'hfff;
rom[2409] = 12'hfff;
rom[2410] = 12'hfff;
rom[2411] = 12'hfff;
rom[2412] = 12'hfff;
rom[2413] = 12'hfff;
rom[2414] = 12'hfff;
rom[2415] = 12'hfff;
rom[2416] = 12'hfff;
rom[2417] = 12'hfff;
rom[2418] = 12'hfff;
rom[2419] = 12'hfff;
rom[2420] = 12'hfff;
rom[2421] = 12'hfff;
rom[2422] = 12'hfff;
rom[2423] = 12'hfff;
rom[2424] = 12'hfff;
rom[2425] = 12'hfff;
rom[2426] = 12'hfff;
rom[2427] = 12'hfff;
rom[2428] = 12'hfff;
rom[2429] = 12'hfff;
rom[2430] = 12'hfff;
rom[2431] = 12'hfff;
rom[2432] = 12'hfff;
rom[2433] = 12'hfff;
rom[2434] = 12'hfff;
rom[2435] = 12'hfff;
rom[2436] = 12'hfff;
rom[2437] = 12'hfff;
rom[2438] = 12'hfff;
rom[2439] = 12'hfff;
rom[2440] = 12'hfff;
rom[2441] = 12'hfff;
rom[2442] = 12'hfff;
rom[2443] = 12'hfff;
rom[2444] = 12'hfff;
rom[2445] = 12'hfff;
rom[2446] = 12'hfff;
rom[2447] = 12'hfff;
rom[2448] = 12'hfff;
rom[2449] = 12'hfff;
rom[2450] = 12'hfff;
rom[2451] = 12'hfff;
rom[2452] = 12'hfff;
rom[2453] = 12'hfff;
rom[2454] = 12'hfff;
rom[2455] = 12'hfff;
rom[2456] = 12'hfff;
rom[2457] = 12'hfff;
rom[2458] = 12'hfff;
rom[2459] = 12'hfff;
rom[2460] = 12'hfff;
rom[2461] = 12'hfff;
rom[2462] = 12'hfff;
rom[2463] = 12'hfff;
rom[2464] = 12'hfff;
rom[2465] = 12'hfff;
rom[2466] = 12'hfff;
rom[2467] = 12'hfff;
rom[2468] = 12'hfff;
rom[2469] = 12'hfff;
rom[2470] = 12'hfff;
rom[2471] = 12'hfff;
rom[2472] = 12'hfff;
rom[2473] = 12'hfff;
rom[2474] = 12'hfff;
rom[2475] = 12'hfff;
rom[2476] = 12'hfff;
rom[2477] = 12'hfff;
rom[2478] = 12'hfff;
rom[2479] = 12'hfff;
rom[2480] = 12'hfff;
rom[2481] = 12'hfff;
rom[2482] = 12'hfff;
rom[2483] = 12'hfff;
rom[2484] = 12'hfff;
rom[2485] = 12'hfff;
rom[2486] = 12'hfff;
rom[2487] = 12'hfff;
rom[2488] = 12'hfff;
rom[2489] = 12'hfff;
rom[2490] = 12'hfff;
rom[2491] = 12'hfff;
rom[2492] = 12'hfff;
rom[2493] = 12'hfff;
rom[2494] = 12'hfff;
rom[2495] = 12'hfff;
rom[2496] = 12'hfff;
rom[2497] = 12'hfff;
rom[2498] = 12'hfff;
rom[2499] = 12'hfff;
rom[2500] = 12'hfff;
rom[2501] = 12'hfff;
rom[2502] = 12'hfff;
rom[2503] = 12'hfff;
rom[2504] = 12'hfff;
rom[2505] = 12'hfff;
rom[2506] = 12'hfff;
rom[2507] = 12'hfff;
rom[2508] = 12'hfff;
rom[2509] = 12'hfff;
rom[2510] = 12'hfff;
rom[2511] = 12'hfff;
rom[2512] = 12'hfff;
rom[2513] = 12'hfff;
rom[2514] = 12'hfff;
rom[2515] = 12'hfff;
rom[2516] = 12'hfff;
rom[2517] = 12'hfff;
rom[2518] = 12'hfff;
rom[2519] = 12'hfff;
rom[2520] = 12'hfff;
rom[2521] = 12'hfff;
rom[2522] = 12'hfff;
rom[2523] = 12'hfff;
rom[2524] = 12'hfff;
rom[2525] = 12'hfff;
rom[2526] = 12'hfff;
rom[2527] = 12'hfff;
rom[2528] = 12'hfff;
rom[2529] = 12'hfff;
rom[2530] = 12'hfff;
rom[2531] = 12'hfff;
rom[2532] = 12'hfff;
rom[2533] = 12'hfff;
rom[2534] = 12'hfff;
rom[2535] = 12'hfff;
rom[2536] = 12'hfff;
rom[2537] = 12'hfff;
rom[2538] = 12'hfff;
rom[2539] = 12'hfff;
rom[2540] = 12'hfff;
rom[2541] = 12'hfff;
rom[2542] = 12'hfff;
rom[2543] = 12'hfff;
rom[2544] = 12'hfff;
rom[2545] = 12'hfff;
rom[2546] = 12'hfff;
rom[2547] = 12'hfff;
rom[2548] = 12'hfff;
rom[2549] = 12'hfff;
rom[2550] = 12'hfff;
rom[2551] = 12'hfff;
rom[2552] = 12'hfff;
rom[2553] = 12'hfff;
rom[2554] = 12'hfff;
rom[2555] = 12'hfff;
rom[2556] = 12'hfff;
rom[2557] = 12'hfff;
rom[2558] = 12'hfff;
rom[2559] = 12'hfff;
rom[2560] = 12'hfff;
rom[2561] = 12'hfff;
rom[2562] = 12'hfff;
rom[2563] = 12'hfff;
rom[2564] = 12'hfff;
rom[2565] = 12'hfff;
rom[2566] = 12'hfff;
rom[2567] = 12'hfff;
rom[2568] = 12'hfff;
rom[2569] = 12'hfff;
rom[2570] = 12'hfff;
rom[2571] = 12'hfff;
rom[2572] = 12'hfff;
rom[2573] = 12'hfff;
rom[2574] = 12'hfff;
rom[2575] = 12'hfff;
rom[2576] = 12'hfff;
rom[2577] = 12'hfff;
rom[2578] = 12'hfff;
rom[2579] = 12'hfff;
rom[2580] = 12'hfff;
rom[2581] = 12'hfff;
rom[2582] = 12'hfff;
rom[2583] = 12'hfff;
rom[2584] = 12'heef;
rom[2585] = 12'h99e;
rom[2586] = 12'h77e;
rom[2587] = 12'h66e;
rom[2588] = 12'h99e;
rom[2589] = 12'hccf;
rom[2590] = 12'heef;
rom[2591] = 12'hfff;
rom[2592] = 12'hfff;
rom[2593] = 12'hfff;
rom[2594] = 12'hfff;
rom[2595] = 12'hfff;
rom[2596] = 12'hfff;
rom[2597] = 12'hfff;
rom[2598] = 12'hfff;
rom[2599] = 12'hfff;
rom[2600] = 12'hfff;
rom[2601] = 12'hfff;
rom[2602] = 12'hfff;
rom[2603] = 12'hfff;
rom[2604] = 12'hfff;
rom[2605] = 12'hfff;
rom[2606] = 12'hfff;
rom[2607] = 12'hfff;
rom[2608] = 12'hfff;
rom[2609] = 12'hfff;
rom[2610] = 12'hfff;
rom[2611] = 12'hfff;
rom[2612] = 12'hfff;
rom[2613] = 12'hfff;
rom[2614] = 12'hfff;
rom[2615] = 12'hfff;
rom[2616] = 12'hfff;
rom[2617] = 12'hfff;
rom[2618] = 12'hfff;
rom[2619] = 12'hfff;
rom[2620] = 12'hfff;
rom[2621] = 12'hfff;
rom[2622] = 12'hfff;
rom[2623] = 12'hfff;
rom[2624] = 12'hfff;
rom[2625] = 12'hfff;
rom[2626] = 12'hfff;
rom[2627] = 12'hfff;
rom[2628] = 12'hfff;
rom[2629] = 12'hfff;
rom[2630] = 12'hfff;
rom[2631] = 12'hfff;
rom[2632] = 12'hfff;
rom[2633] = 12'hfff;
rom[2634] = 12'hfff;
rom[2635] = 12'hfff;
rom[2636] = 12'hfff;
rom[2637] = 12'hfff;
rom[2638] = 12'hfff;
rom[2639] = 12'hfff;
rom[2640] = 12'hfff;
rom[2641] = 12'hfff;
rom[2642] = 12'hfff;
rom[2643] = 12'hfff;
rom[2644] = 12'hfff;
rom[2645] = 12'hfff;
rom[2646] = 12'hfff;
rom[2647] = 12'hfff;
rom[2648] = 12'hfff;
rom[2649] = 12'hfff;
rom[2650] = 12'hfff;
rom[2651] = 12'hfff;
rom[2652] = 12'hfff;
rom[2653] = 12'hfff;
rom[2654] = 12'hfff;
rom[2655] = 12'hfff;
rom[2656] = 12'hfff;
rom[2657] = 12'hfff;
rom[2658] = 12'hfff;
rom[2659] = 12'hfff;
rom[2660] = 12'hfff;
rom[2661] = 12'hfff;
rom[2662] = 12'hfff;
rom[2663] = 12'hfff;
rom[2664] = 12'hfff;
rom[2665] = 12'hfff;
rom[2666] = 12'hfff;
rom[2667] = 12'hfff;
rom[2668] = 12'hfff;
rom[2669] = 12'hfff;
rom[2670] = 12'hfff;
rom[2671] = 12'hfff;
rom[2672] = 12'hfff;
rom[2673] = 12'hfff;
rom[2674] = 12'hfff;
rom[2675] = 12'hfff;
rom[2676] = 12'hfff;
rom[2677] = 12'hfff;
rom[2678] = 12'hfff;
rom[2679] = 12'hfff;
rom[2680] = 12'hfff;
rom[2681] = 12'hfff;
rom[2682] = 12'hfff;
rom[2683] = 12'hfff;
rom[2684] = 12'hfff;
rom[2685] = 12'hfff;
rom[2686] = 12'hfff;
rom[2687] = 12'hfff;
rom[2688] = 12'hfff;
rom[2689] = 12'hfff;
rom[2690] = 12'hfff;
rom[2691] = 12'hfff;
rom[2692] = 12'hfff;
rom[2693] = 12'hfff;
rom[2694] = 12'hfff;
rom[2695] = 12'hfff;
rom[2696] = 12'hfff;
rom[2697] = 12'hfff;
rom[2698] = 12'hfff;
rom[2699] = 12'hfff;
rom[2700] = 12'hfff;
rom[2701] = 12'hfff;
rom[2702] = 12'hfff;
rom[2703] = 12'hfff;
rom[2704] = 12'hfff;
rom[2705] = 12'hfff;
rom[2706] = 12'hfff;
rom[2707] = 12'hfff;
rom[2708] = 12'hfff;
rom[2709] = 12'hfff;
rom[2710] = 12'hfff;
rom[2711] = 12'heef;
rom[2712] = 12'h11d;
rom[2713] = 12'h  c;
rom[2714] = 12'h  c;
rom[2715] = 12'h  c;
rom[2716] = 12'h  c;
rom[2717] = 12'h  c;
rom[2718] = 12'h22d;
rom[2719] = 12'heef;
rom[2720] = 12'hfff;
rom[2721] = 12'hfff;
rom[2722] = 12'hfff;
rom[2723] = 12'hfff;
rom[2724] = 12'hfff;
rom[2725] = 12'hfff;
rom[2726] = 12'hfff;
rom[2727] = 12'hfff;
rom[2728] = 12'hfff;
rom[2729] = 12'hfff;
rom[2730] = 12'hfff;
rom[2731] = 12'hfff;
rom[2732] = 12'hfff;
rom[2733] = 12'hfff;
rom[2734] = 12'hfff;
rom[2735] = 12'hfff;
rom[2736] = 12'hfff;
rom[2737] = 12'hfff;
rom[2738] = 12'hfff;
rom[2739] = 12'hfff;
rom[2740] = 12'hfff;
rom[2741] = 12'hfff;
rom[2742] = 12'hfff;
rom[2743] = 12'hfff;
rom[2744] = 12'hfff;
rom[2745] = 12'hfff;
rom[2746] = 12'hfff;
rom[2747] = 12'hfff;
rom[2748] = 12'hfff;
rom[2749] = 12'hfff;
rom[2750] = 12'hfff;
rom[2751] = 12'hfff;
rom[2752] = 12'hfff;
rom[2753] = 12'hfff;
rom[2754] = 12'hfff;
rom[2755] = 12'hfff;
rom[2756] = 12'hfff;
rom[2757] = 12'hfff;
rom[2758] = 12'hfff;
rom[2759] = 12'hfff;
rom[2760] = 12'hfff;
rom[2761] = 12'hfff;
rom[2762] = 12'hfff;
rom[2763] = 12'hfff;
rom[2764] = 12'hfff;
rom[2765] = 12'hfff;
rom[2766] = 12'hfff;
rom[2767] = 12'hfff;
rom[2768] = 12'hfff;
rom[2769] = 12'hfff;
rom[2770] = 12'hfff;
rom[2771] = 12'hfff;
rom[2772] = 12'hfff;
rom[2773] = 12'hfff;
rom[2774] = 12'hfff;
rom[2775] = 12'hfff;
rom[2776] = 12'hfff;
rom[2777] = 12'hfff;
rom[2778] = 12'hfff;
rom[2779] = 12'hfff;
rom[2780] = 12'hfff;
rom[2781] = 12'hfff;
rom[2782] = 12'hfff;
rom[2783] = 12'hfff;
rom[2784] = 12'hfff;
rom[2785] = 12'hfff;
rom[2786] = 12'hfff;
rom[2787] = 12'hfff;
rom[2788] = 12'hfff;
rom[2789] = 12'hfff;
rom[2790] = 12'hfff;
rom[2791] = 12'hfff;
rom[2792] = 12'hfff;
rom[2793] = 12'hfff;
rom[2794] = 12'hfff;
rom[2795] = 12'hfff;
rom[2796] = 12'hfff;
rom[2797] = 12'hfff;
rom[2798] = 12'hfff;
rom[2799] = 12'hfff;
rom[2800] = 12'hfff;
rom[2801] = 12'hfff;
rom[2802] = 12'hfff;
rom[2803] = 12'hfff;
rom[2804] = 12'hfff;
rom[2805] = 12'hfff;
rom[2806] = 12'hfff;
rom[2807] = 12'hfff;
rom[2808] = 12'hfff;
rom[2809] = 12'hfff;
rom[2810] = 12'hfff;
rom[2811] = 12'hfff;
rom[2812] = 12'hfff;
rom[2813] = 12'hfff;
rom[2814] = 12'hfff;
rom[2815] = 12'hfff;
rom[2816] = 12'hfff;
rom[2817] = 12'hfff;
rom[2818] = 12'hfff;
rom[2819] = 12'hfff;
rom[2820] = 12'hfff;
rom[2821] = 12'hfff;
rom[2822] = 12'hfff;
rom[2823] = 12'hfff;
rom[2824] = 12'hfff;
rom[2825] = 12'hfff;
rom[2826] = 12'hfff;
rom[2827] = 12'hfff;
rom[2828] = 12'hfff;
rom[2829] = 12'hfff;
rom[2830] = 12'hfff;
rom[2831] = 12'hfff;
rom[2832] = 12'hfff;
rom[2833] = 12'hfff;
rom[2834] = 12'hfff;
rom[2835] = 12'hfff;
rom[2836] = 12'hfff;
rom[2837] = 12'hfff;
rom[2838] = 12'hfff;
rom[2839] = 12'h99e;
rom[2840] = 12'h  c;
rom[2841] = 12'h  c;
rom[2842] = 12'h  c;
rom[2843] = 12'h  c;
rom[2844] = 12'h  c;
rom[2845] = 12'h  c;
rom[2846] = 12'h  c;
rom[2847] = 12'h11d;
rom[2848] = 12'h88e;
rom[2849] = 12'h77e;
rom[2850] = 12'h77e;
rom[2851] = 12'haae;
rom[2852] = 12'heef;
rom[2853] = 12'hfff;
rom[2854] = 12'hfff;
rom[2855] = 12'hfff;
rom[2856] = 12'hfff;
rom[2857] = 12'hfff;
rom[2858] = 12'hfff;
rom[2859] = 12'hfff;
rom[2860] = 12'hfff;
rom[2861] = 12'hfff;
rom[2862] = 12'hfff;
rom[2863] = 12'hfff;
rom[2864] = 12'hfff;
rom[2865] = 12'hfff;
rom[2866] = 12'hfff;
rom[2867] = 12'hfff;
rom[2868] = 12'hfff;
rom[2869] = 12'hfff;
rom[2870] = 12'hfff;
rom[2871] = 12'hfff;
rom[2872] = 12'hfff;
rom[2873] = 12'hfff;
rom[2874] = 12'hfff;
rom[2875] = 12'hfff;
rom[2876] = 12'hfff;
rom[2877] = 12'hfff;
rom[2878] = 12'hfff;
rom[2879] = 12'hfff;
rom[2880] = 12'hfff;
rom[2881] = 12'hfff;
rom[2882] = 12'hfff;
rom[2883] = 12'hfff;
rom[2884] = 12'hfff;
rom[2885] = 12'hfff;
rom[2886] = 12'hfff;
rom[2887] = 12'hfff;
rom[2888] = 12'hfff;
rom[2889] = 12'hfff;
rom[2890] = 12'hfff;
rom[2891] = 12'hfff;
rom[2892] = 12'hfff;
rom[2893] = 12'hfff;
rom[2894] = 12'hfff;
rom[2895] = 12'hfff;
rom[2896] = 12'hfff;
rom[2897] = 12'hfff;
rom[2898] = 12'hfff;
rom[2899] = 12'hfff;
rom[2900] = 12'hfff;
rom[2901] = 12'hfff;
rom[2902] = 12'hfff;
rom[2903] = 12'hfff;
rom[2904] = 12'hfff;
rom[2905] = 12'hfff;
rom[2906] = 12'hfff;
rom[2907] = 12'hfff;
rom[2908] = 12'hfff;
rom[2909] = 12'hfff;
rom[2910] = 12'hfff;
rom[2911] = 12'hfff;
rom[2912] = 12'hfff;
rom[2913] = 12'hfff;
rom[2914] = 12'hfff;
rom[2915] = 12'hfff;
rom[2916] = 12'hfff;
rom[2917] = 12'hfff;
rom[2918] = 12'hfff;
rom[2919] = 12'hfff;
rom[2920] = 12'hfff;
rom[2921] = 12'hfff;
rom[2922] = 12'hfff;
rom[2923] = 12'hfff;
rom[2924] = 12'hfff;
rom[2925] = 12'hfff;
rom[2926] = 12'hfff;
rom[2927] = 12'hfff;
rom[2928] = 12'hfff;
rom[2929] = 12'hfff;
rom[2930] = 12'hfff;
rom[2931] = 12'hfff;
rom[2932] = 12'hfff;
rom[2933] = 12'hfff;
rom[2934] = 12'hfff;
rom[2935] = 12'hfff;
rom[2936] = 12'hfff;
rom[2937] = 12'hfff;
rom[2938] = 12'hfff;
rom[2939] = 12'hfff;
rom[2940] = 12'hfff;
rom[2941] = 12'hfff;
rom[2942] = 12'hfff;
rom[2943] = 12'hfff;
rom[2944] = 12'hfff;
rom[2945] = 12'hfff;
rom[2946] = 12'hfff;
rom[2947] = 12'hfff;
rom[2948] = 12'hfff;
rom[2949] = 12'hfff;
rom[2950] = 12'hfff;
rom[2951] = 12'hfff;
rom[2952] = 12'hfff;
rom[2953] = 12'hfff;
rom[2954] = 12'hfff;
rom[2955] = 12'hfff;
rom[2956] = 12'hfff;
rom[2957] = 12'hfff;
rom[2958] = 12'hfff;
rom[2959] = 12'hfff;
rom[2960] = 12'hfff;
rom[2961] = 12'hfff;
rom[2962] = 12'hfff;
rom[2963] = 12'hfff;
rom[2964] = 12'hfff;
rom[2965] = 12'hfff;
rom[2966] = 12'hfff;
rom[2967] = 12'h99e;
rom[2968] = 12'h  c;
rom[2969] = 12'h  c;
rom[2970] = 12'h  c;
rom[2971] = 12'h  c;
rom[2972] = 12'h  c;
rom[2973] = 12'h  c;
rom[2974] = 12'h  c;
rom[2975] = 12'h  c;
rom[2976] = 12'h11d;
rom[2977] = 12'h  c;
rom[2978] = 12'h  c;
rom[2979] = 12'h  c;
rom[2980] = 12'h22d;
rom[2981] = 12'heef;
rom[2982] = 12'hfff;
rom[2983] = 12'hfff;
rom[2984] = 12'hfff;
rom[2985] = 12'hfff;
rom[2986] = 12'hfff;
rom[2987] = 12'hfff;
rom[2988] = 12'hfff;
rom[2989] = 12'hfff;
rom[2990] = 12'hfff;
rom[2991] = 12'hfff;
rom[2992] = 12'hfff;
rom[2993] = 12'hfff;
rom[2994] = 12'hfff;
rom[2995] = 12'hfff;
rom[2996] = 12'hfff;
rom[2997] = 12'hfff;
rom[2998] = 12'hfff;
rom[2999] = 12'hfff;
rom[3000] = 12'hfff;
rom[3001] = 12'hfff;
rom[3002] = 12'hfff;
rom[3003] = 12'hfff;
rom[3004] = 12'hfff;
rom[3005] = 12'hfff;
rom[3006] = 12'hfff;
rom[3007] = 12'hfff;
rom[3008] = 12'hfff;
rom[3009] = 12'hfff;
rom[3010] = 12'hfff;
rom[3011] = 12'hfff;
rom[3012] = 12'hfff;
rom[3013] = 12'hfff;
rom[3014] = 12'hfff;
rom[3015] = 12'hfff;
rom[3016] = 12'hfff;
rom[3017] = 12'hfff;
rom[3018] = 12'hfff;
rom[3019] = 12'hfff;
rom[3020] = 12'hfff;
rom[3021] = 12'hfff;
rom[3022] = 12'hfff;
rom[3023] = 12'hfff;
rom[3024] = 12'hfff;
rom[3025] = 12'hfff;
rom[3026] = 12'hfff;
rom[3027] = 12'hfff;
rom[3028] = 12'hfff;
rom[3029] = 12'hfff;
rom[3030] = 12'hfff;
rom[3031] = 12'hfff;
rom[3032] = 12'hfff;
rom[3033] = 12'hfff;
rom[3034] = 12'hfff;
rom[3035] = 12'hfff;
rom[3036] = 12'heef;
rom[3037] = 12'h99e;
rom[3038] = 12'h77e;
rom[3039] = 12'h77e;
rom[3040] = 12'h66e;
rom[3041] = 12'h66d;
rom[3042] = 12'h55d;
rom[3043] = 12'h44d;
rom[3044] = 12'h44d;
rom[3045] = 12'h44d;
rom[3046] = 12'h44d;
rom[3047] = 12'h44d;
rom[3048] = 12'h44d;
rom[3049] = 12'h44d;
rom[3050] = 12'h44d;
rom[3051] = 12'h66e;
rom[3052] = 12'h99e;
rom[3053] = 12'hfff;
rom[3054] = 12'hfff;
rom[3055] = 12'hfff;
rom[3056] = 12'hfff;
rom[3057] = 12'hfff;
rom[3058] = 12'hfff;
rom[3059] = 12'hfff;
rom[3060] = 12'hfff;
rom[3061] = 12'hfff;
rom[3062] = 12'hfff;
rom[3063] = 12'hfff;
rom[3064] = 12'hfff;
rom[3065] = 12'hfff;
rom[3066] = 12'hfff;
rom[3067] = 12'hfff;
rom[3068] = 12'hfff;
rom[3069] = 12'hfff;
rom[3070] = 12'hfff;
rom[3071] = 12'hfff;
rom[3072] = 12'hfff;
rom[3073] = 12'hfff;
rom[3074] = 12'hfff;
rom[3075] = 12'hfff;
rom[3076] = 12'hfff;
rom[3077] = 12'hfff;
rom[3078] = 12'hfff;
rom[3079] = 12'hfff;
rom[3080] = 12'hfff;
rom[3081] = 12'hfff;
rom[3082] = 12'hfff;
rom[3083] = 12'hfff;
rom[3084] = 12'hfff;
rom[3085] = 12'hfff;
rom[3086] = 12'hfff;
rom[3087] = 12'hfff;
rom[3088] = 12'hfff;
rom[3089] = 12'hfff;
rom[3090] = 12'hfff;
rom[3091] = 12'hfff;
rom[3092] = 12'hfff;
rom[3093] = 12'hfff;
rom[3094] = 12'hfff;
rom[3095] = 12'heef;
rom[3096] = 12'h11d;
rom[3097] = 12'h  c;
rom[3098] = 12'h  c;
rom[3099] = 12'h  c;
rom[3100] = 12'h  c;
rom[3101] = 12'h  c;
rom[3102] = 12'h  c;
rom[3103] = 12'h  c;
rom[3104] = 12'h  c;
rom[3105] = 12'h  c;
rom[3106] = 12'h  c;
rom[3107] = 12'h  c;
rom[3108] = 12'h  c;
rom[3109] = 12'h11d;
rom[3110] = 12'hccf;
rom[3111] = 12'heef;
rom[3112] = 12'hfff;
rom[3113] = 12'hfff;
rom[3114] = 12'hfff;
rom[3115] = 12'hfff;
rom[3116] = 12'hfff;
rom[3117] = 12'hfff;
rom[3118] = 12'hfff;
rom[3119] = 12'hfff;
rom[3120] = 12'hfff;
rom[3121] = 12'hfff;
rom[3122] = 12'hfff;
rom[3123] = 12'hfff;
rom[3124] = 12'hfff;
rom[3125] = 12'hfff;
rom[3126] = 12'hfff;
rom[3127] = 12'hfff;
rom[3128] = 12'hfff;
rom[3129] = 12'hfff;
rom[3130] = 12'hfff;
rom[3131] = 12'hfff;
rom[3132] = 12'hfff;
rom[3133] = 12'hfff;
rom[3134] = 12'hfff;
rom[3135] = 12'hfff;
rom[3136] = 12'hfff;
rom[3137] = 12'hfff;
rom[3138] = 12'hfff;
rom[3139] = 12'hfff;
rom[3140] = 12'hfff;
rom[3141] = 12'hfff;
rom[3142] = 12'hfff;
rom[3143] = 12'hfff;
rom[3144] = 12'hfff;
rom[3145] = 12'hfff;
rom[3146] = 12'hfff;
rom[3147] = 12'hfff;
rom[3148] = 12'hfff;
rom[3149] = 12'hfff;
rom[3150] = 12'hfff;
rom[3151] = 12'hfff;
rom[3152] = 12'hfff;
rom[3153] = 12'hfff;
rom[3154] = 12'hfff;
rom[3155] = 12'hfff;
rom[3156] = 12'hfff;
rom[3157] = 12'hfff;
rom[3158] = 12'haae;
rom[3159] = 12'h88e;
rom[3160] = 12'h55d;
rom[3161] = 12'h55d;
rom[3162] = 12'h55d;
rom[3163] = 12'h55d;
rom[3164] = 12'h11d;
rom[3165] = 12'h  c;
rom[3166] = 12'h  c;
rom[3167] = 12'h  c;
rom[3168] = 12'h  c;
rom[3169] = 12'h  c;
rom[3170] = 12'h  c;
rom[3171] = 12'h  c;
rom[3172] = 12'h  c;
rom[3173] = 12'h  c;
rom[3174] = 12'h  c;
rom[3175] = 12'h  c;
rom[3176] = 12'h  c;
rom[3177] = 12'h  c;
rom[3178] = 12'h  c;
rom[3179] = 12'h  c;
rom[3180] = 12'h  c;
rom[3181] = 12'h22d;
rom[3182] = 12'h88e;
rom[3183] = 12'heef;
rom[3184] = 12'hfff;
rom[3185] = 12'hfff;
rom[3186] = 12'hfff;
rom[3187] = 12'hfff;
rom[3188] = 12'hfff;
rom[3189] = 12'hfff;
rom[3190] = 12'hfff;
rom[3191] = 12'hfff;
rom[3192] = 12'hfff;
rom[3193] = 12'hfff;
rom[3194] = 12'hfff;
rom[3195] = 12'hfff;
rom[3196] = 12'hfff;
rom[3197] = 12'hfff;
rom[3198] = 12'hfff;
rom[3199] = 12'hfff;
rom[3200] = 12'hfff;
rom[3201] = 12'hfff;
rom[3202] = 12'hfff;
rom[3203] = 12'hfff;
rom[3204] = 12'hfff;
rom[3205] = 12'hfff;
rom[3206] = 12'hfff;
rom[3207] = 12'hfff;
rom[3208] = 12'hfff;
rom[3209] = 12'hfff;
rom[3210] = 12'hfff;
rom[3211] = 12'hfff;
rom[3212] = 12'hfff;
rom[3213] = 12'hfff;
rom[3214] = 12'hfff;
rom[3215] = 12'hfff;
rom[3216] = 12'hfff;
rom[3217] = 12'hfff;
rom[3218] = 12'hfff;
rom[3219] = 12'hfff;
rom[3220] = 12'hfff;
rom[3221] = 12'hfff;
rom[3222] = 12'hfff;
rom[3223] = 12'hfff;
rom[3224] = 12'heef;
rom[3225] = 12'h99e;
rom[3226] = 12'h88e;
rom[3227] = 12'h99e;
rom[3228] = 12'h77e;
rom[3229] = 12'h22d;
rom[3230] = 12'h  c;
rom[3231] = 12'h  c;
rom[3232] = 12'h  c;
rom[3233] = 12'h  c;
rom[3234] = 12'h  c;
rom[3235] = 12'h  c;
rom[3236] = 12'h  c;
rom[3237] = 12'h  c;
rom[3238] = 12'h  c;
rom[3239] = 12'h22d;
rom[3240] = 12'heef;
rom[3241] = 12'hfff;
rom[3242] = 12'hfff;
rom[3243] = 12'hfff;
rom[3244] = 12'hfff;
rom[3245] = 12'hfff;
rom[3246] = 12'hfff;
rom[3247] = 12'hfff;
rom[3248] = 12'hfff;
rom[3249] = 12'hfff;
rom[3250] = 12'hfff;
rom[3251] = 12'hfff;
rom[3252] = 12'hfff;
rom[3253] = 12'hfff;
rom[3254] = 12'hfff;
rom[3255] = 12'hfff;
rom[3256] = 12'hfff;
rom[3257] = 12'hfff;
rom[3258] = 12'hfff;
rom[3259] = 12'hfff;
rom[3260] = 12'hfff;
rom[3261] = 12'hfff;
rom[3262] = 12'hfff;
rom[3263] = 12'hfff;
rom[3264] = 12'hfff;
rom[3265] = 12'hfff;
rom[3266] = 12'hfff;
rom[3267] = 12'hfff;
rom[3268] = 12'hfff;
rom[3269] = 12'hfff;
rom[3270] = 12'hfff;
rom[3271] = 12'hfff;
rom[3272] = 12'hfff;
rom[3273] = 12'hfff;
rom[3274] = 12'hfff;
rom[3275] = 12'hfff;
rom[3276] = 12'hfff;
rom[3277] = 12'hfff;
rom[3278] = 12'hfff;
rom[3279] = 12'hfff;
rom[3280] = 12'hfff;
rom[3281] = 12'hfff;
rom[3282] = 12'heef;
rom[3283] = 12'h99e;
rom[3284] = 12'h99e;
rom[3285] = 12'h33d;
rom[3286] = 12'h  c;
rom[3287] = 12'h  c;
rom[3288] = 12'h  c;
rom[3289] = 12'h  c;
rom[3290] = 12'h  c;
rom[3291] = 12'h  c;
rom[3292] = 12'h  c;
rom[3293] = 12'h  c;
rom[3294] = 12'h  c;
rom[3295] = 12'h  c;
rom[3296] = 12'h  c;
rom[3297] = 12'h  c;
rom[3298] = 12'h  c;
rom[3299] = 12'h  c;
rom[3300] = 12'h  c;
rom[3301] = 12'h  c;
rom[3302] = 12'h  c;
rom[3303] = 12'h  c;
rom[3304] = 12'h  c;
rom[3305] = 12'h  c;
rom[3306] = 12'h  c;
rom[3307] = 12'h  c;
rom[3308] = 12'h  c;
rom[3309] = 12'h  c;
rom[3310] = 12'h  c;
rom[3311] = 12'h22d;
rom[3312] = 12'h99e;
rom[3313] = 12'h88e;
rom[3314] = 12'h77e;
rom[3315] = 12'h99e;
rom[3316] = 12'heef;
rom[3317] = 12'hfff;
rom[3318] = 12'hfff;
rom[3319] = 12'hfff;
rom[3320] = 12'hfff;
rom[3321] = 12'hfff;
rom[3322] = 12'hfff;
rom[3323] = 12'hfff;
rom[3324] = 12'hfff;
rom[3325] = 12'hfff;
rom[3326] = 12'hfff;
rom[3327] = 12'hfff;
rom[3328] = 12'hfff;
rom[3329] = 12'hfff;
rom[3330] = 12'hfff;
rom[3331] = 12'hfff;
rom[3332] = 12'hfff;
rom[3333] = 12'hfff;
rom[3334] = 12'hfff;
rom[3335] = 12'hfff;
rom[3336] = 12'hfff;
rom[3337] = 12'hfff;
rom[3338] = 12'hfff;
rom[3339] = 12'hfff;
rom[3340] = 12'hfff;
rom[3341] = 12'hfff;
rom[3342] = 12'hfff;
rom[3343] = 12'hfff;
rom[3344] = 12'hfff;
rom[3345] = 12'hfff;
rom[3346] = 12'hfff;
rom[3347] = 12'hfff;
rom[3348] = 12'hfff;
rom[3349] = 12'hfff;
rom[3350] = 12'hfff;
rom[3351] = 12'hfff;
rom[3352] = 12'hfff;
rom[3353] = 12'hfff;
rom[3354] = 12'hfff;
rom[3355] = 12'hfff;
rom[3356] = 12'heef;
rom[3357] = 12'h66d;
rom[3358] = 12'h  c;
rom[3359] = 12'h  c;
rom[3360] = 12'h  c;
rom[3361] = 12'h  c;
rom[3362] = 12'h  c;
rom[3363] = 12'h  c;
rom[3364] = 12'h  c;
rom[3365] = 12'h  c;
rom[3366] = 12'h  c;
rom[3367] = 12'h  c;
rom[3368] = 12'h11d;
rom[3369] = 12'hbbf;
rom[3370] = 12'heef;
rom[3371] = 12'hfff;
rom[3372] = 12'hfff;
rom[3373] = 12'hfff;
rom[3374] = 12'hfff;
rom[3375] = 12'hfff;
rom[3376] = 12'hfff;
rom[3377] = 12'hfff;
rom[3378] = 12'hfff;
rom[3379] = 12'hfff;
rom[3380] = 12'hfff;
rom[3381] = 12'hfff;
rom[3382] = 12'hfff;
rom[3383] = 12'hfff;
rom[3384] = 12'hfff;
rom[3385] = 12'hfff;
rom[3386] = 12'hfff;
rom[3387] = 12'hfff;
rom[3388] = 12'hfff;
rom[3389] = 12'hfff;
rom[3390] = 12'hfff;
rom[3391] = 12'hfff;
rom[3392] = 12'hfff;
rom[3393] = 12'hfff;
rom[3394] = 12'hfff;
rom[3395] = 12'hfff;
rom[3396] = 12'hfff;
rom[3397] = 12'hfff;
rom[3398] = 12'hfff;
rom[3399] = 12'hfff;
rom[3400] = 12'hfff;
rom[3401] = 12'hfff;
rom[3402] = 12'hfff;
rom[3403] = 12'hfff;
rom[3404] = 12'hfff;
rom[3405] = 12'hfff;
rom[3406] = 12'hfff;
rom[3407] = 12'hfff;
rom[3408] = 12'hfff;
rom[3409] = 12'h99e;
rom[3410] = 12'h11d;
rom[3411] = 12'h  c;
rom[3412] = 12'h  c;
rom[3413] = 12'h  c;
rom[3414] = 12'h  c;
rom[3415] = 12'h  c;
rom[3416] = 12'h  c;
rom[3417] = 12'h  c;
rom[3418] = 12'h  c;
rom[3419] = 12'h  c;
rom[3420] = 12'h  c;
rom[3421] = 12'h  c;
rom[3422] = 12'h  c;
rom[3423] = 12'h  c;
rom[3424] = 12'h  c;
rom[3425] = 12'h  c;
rom[3426] = 12'h  c;
rom[3427] = 12'h  c;
rom[3428] = 12'h  c;
rom[3429] = 12'h  c;
rom[3430] = 12'h  c;
rom[3431] = 12'h  c;
rom[3432] = 12'h  c;
rom[3433] = 12'h  c;
rom[3434] = 12'h  c;
rom[3435] = 12'h  c;
rom[3436] = 12'h  c;
rom[3437] = 12'h  c;
rom[3438] = 12'h  c;
rom[3439] = 12'h  c;
rom[3440] = 12'h  c;
rom[3441] = 12'h  c;
rom[3442] = 12'h  c;
rom[3443] = 12'h  c;
rom[3444] = 12'h33d;
rom[3445] = 12'heef;
rom[3446] = 12'hfff;
rom[3447] = 12'hfff;
rom[3448] = 12'hfff;
rom[3449] = 12'hfff;
rom[3450] = 12'hfff;
rom[3451] = 12'hfff;
rom[3452] = 12'hfff;
rom[3453] = 12'hfff;
rom[3454] = 12'hfff;
rom[3455] = 12'hfff;
rom[3456] = 12'hfff;
rom[3457] = 12'hfff;
rom[3458] = 12'hfff;
rom[3459] = 12'hfff;
rom[3460] = 12'hfff;
rom[3461] = 12'hfff;
rom[3462] = 12'hfff;
rom[3463] = 12'hfff;
rom[3464] = 12'hfff;
rom[3465] = 12'hfff;
rom[3466] = 12'hfff;
rom[3467] = 12'hfff;
rom[3468] = 12'hfff;
rom[3469] = 12'hfff;
rom[3470] = 12'hfff;
rom[3471] = 12'hfff;
rom[3472] = 12'hfff;
rom[3473] = 12'hfff;
rom[3474] = 12'hfff;
rom[3475] = 12'hfff;
rom[3476] = 12'hfff;
rom[3477] = 12'hfff;
rom[3478] = 12'hfff;
rom[3479] = 12'hfff;
rom[3480] = 12'hfff;
rom[3481] = 12'hfff;
rom[3482] = 12'hfff;
rom[3483] = 12'hfff;
rom[3484] = 12'hfff;
rom[3485] = 12'heef;
rom[3486] = 12'h99e;
rom[3487] = 12'h77e;
rom[3488] = 12'h77e;
rom[3489] = 12'h88e;
rom[3490] = 12'h77e;
rom[3491] = 12'h22d;
rom[3492] = 12'h  c;
rom[3493] = 12'h  c;
rom[3494] = 12'h  c;
rom[3495] = 12'h  c;
rom[3496] = 12'h  c;
rom[3497] = 12'h  c;
rom[3498] = 12'h11d;
rom[3499] = 12'hccf;
rom[3500] = 12'hfff;
rom[3501] = 12'hfff;
rom[3502] = 12'hfff;
rom[3503] = 12'hfff;
rom[3504] = 12'hfff;
rom[3505] = 12'hfff;
rom[3506] = 12'hfff;
rom[3507] = 12'hfff;
rom[3508] = 12'hfff;
rom[3509] = 12'hfff;
rom[3510] = 12'hfff;
rom[3511] = 12'hfff;
rom[3512] = 12'hfff;
rom[3513] = 12'hfff;
rom[3514] = 12'hfff;
rom[3515] = 12'hfff;
rom[3516] = 12'hfff;
rom[3517] = 12'hfff;
rom[3518] = 12'hfff;
rom[3519] = 12'hfff;
rom[3520] = 12'hfff;
rom[3521] = 12'hfff;
rom[3522] = 12'hfff;
rom[3523] = 12'hfff;
rom[3524] = 12'hfff;
rom[3525] = 12'hfff;
rom[3526] = 12'hfff;
rom[3527] = 12'hfff;
rom[3528] = 12'hfff;
rom[3529] = 12'hfff;
rom[3530] = 12'hfff;
rom[3531] = 12'hfff;
rom[3532] = 12'hfff;
rom[3533] = 12'heef;
rom[3534] = 12'h99e;
rom[3535] = 12'hccf;
rom[3536] = 12'h44d;
rom[3537] = 12'h  c;
rom[3538] = 12'h  c;
rom[3539] = 12'h  c;
rom[3540] = 12'h  c;
rom[3541] = 12'h  c;
rom[3542] = 12'h  c;
rom[3543] = 12'h  c;
rom[3544] = 12'h  c;
rom[3545] = 12'h  c;
rom[3546] = 12'h  c;
rom[3547] = 12'h  c;
rom[3548] = 12'h  c;
rom[3549] = 12'h  c;
rom[3550] = 12'h  c;
rom[3551] = 12'h  c;
rom[3552] = 12'h  c;
rom[3553] = 12'h  c;
rom[3554] = 12'h  c;
rom[3555] = 12'h  c;
rom[3556] = 12'h  c;
rom[3557] = 12'h  c;
rom[3558] = 12'h  c;
rom[3559] = 12'h  c;
rom[3560] = 12'h  c;
rom[3561] = 12'h  c;
rom[3562] = 12'h  c;
rom[3563] = 12'h  c;
rom[3564] = 12'h  c;
rom[3565] = 12'h  c;
rom[3566] = 12'h  c;
rom[3567] = 12'h  c;
rom[3568] = 12'h  c;
rom[3569] = 12'h  c;
rom[3570] = 12'h  c;
rom[3571] = 12'h  c;
rom[3572] = 12'h  c;
rom[3573] = 12'h11d;
rom[3574] = 12'h99e;
rom[3575] = 12'hfff;
rom[3576] = 12'hfff;
rom[3577] = 12'hfff;
rom[3578] = 12'hfff;
rom[3579] = 12'hfff;
rom[3580] = 12'hfff;
rom[3581] = 12'hfff;
rom[3582] = 12'hfff;
rom[3583] = 12'hfff;
rom[3584] = 12'hfff;
rom[3585] = 12'hfff;
rom[3586] = 12'hfff;
rom[3587] = 12'hfff;
rom[3588] = 12'hfff;
rom[3589] = 12'hfff;
rom[3590] = 12'hfff;
rom[3591] = 12'hfff;
rom[3592] = 12'hfff;
rom[3593] = 12'hfff;
rom[3594] = 12'hfff;
rom[3595] = 12'hfff;
rom[3596] = 12'hfff;
rom[3597] = 12'hfff;
rom[3598] = 12'hfff;
rom[3599] = 12'hfff;
rom[3600] = 12'hfff;
rom[3601] = 12'hfff;
rom[3602] = 12'hfff;
rom[3603] = 12'hfff;
rom[3604] = 12'hfff;
rom[3605] = 12'hfff;
rom[3606] = 12'hfff;
rom[3607] = 12'hfff;
rom[3608] = 12'hfff;
rom[3609] = 12'hfff;
rom[3610] = 12'hfff;
rom[3611] = 12'hfff;
rom[3612] = 12'hfff;
rom[3613] = 12'hfff;
rom[3614] = 12'hfff;
rom[3615] = 12'hfff;
rom[3616] = 12'hfff;
rom[3617] = 12'hfff;
rom[3618] = 12'heef;
rom[3619] = 12'h77e;
rom[3620] = 12'h11d;
rom[3621] = 12'h  c;
rom[3622] = 12'h  c;
rom[3623] = 12'h  c;
rom[3624] = 12'h  c;
rom[3625] = 12'h  c;
rom[3626] = 12'h  c;
rom[3627] = 12'h  c;
rom[3628] = 12'hddf;
rom[3629] = 12'hfff;
rom[3630] = 12'hfff;
rom[3631] = 12'hfff;
rom[3632] = 12'hfff;
rom[3633] = 12'hfff;
rom[3634] = 12'hfff;
rom[3635] = 12'hfff;
rom[3636] = 12'hfff;
rom[3637] = 12'hfff;
rom[3638] = 12'hfff;
rom[3639] = 12'hfff;
rom[3640] = 12'hfff;
rom[3641] = 12'hfff;
rom[3642] = 12'hfff;
rom[3643] = 12'hfff;
rom[3644] = 12'hfff;
rom[3645] = 12'hfff;
rom[3646] = 12'hfff;
rom[3647] = 12'hfff;
rom[3648] = 12'hfff;
rom[3649] = 12'hfff;
rom[3650] = 12'hfff;
rom[3651] = 12'hfff;
rom[3652] = 12'hfff;
rom[3653] = 12'hfff;
rom[3654] = 12'hfff;
rom[3655] = 12'hfff;
rom[3656] = 12'hfff;
rom[3657] = 12'hfff;
rom[3658] = 12'hfff;
rom[3659] = 12'hfff;
rom[3660] = 12'heef;
rom[3661] = 12'h11d;
rom[3662] = 12'h  c;
rom[3663] = 12'h11d;
rom[3664] = 12'h  c;
rom[3665] = 12'h  c;
rom[3666] = 12'h  c;
rom[3667] = 12'h  c;
rom[3668] = 12'h  c;
rom[3669] = 12'h  c;
rom[3670] = 12'h  c;
rom[3671] = 12'h  c;
rom[3672] = 12'h  c;
rom[3673] = 12'h  c;
rom[3674] = 12'h  c;
rom[3675] = 12'h  c;
rom[3676] = 12'h  c;
rom[3677] = 12'h  c;
rom[3678] = 12'h  c;
rom[3679] = 12'h  c;
rom[3680] = 12'h  c;
rom[3681] = 12'h  c;
rom[3682] = 12'h11d;
rom[3683] = 12'haae;
rom[3684] = 12'hbbf;
rom[3685] = 12'hbbf;
rom[3686] = 12'hbbf;
rom[3687] = 12'hbbf;
rom[3688] = 12'hbbf;
rom[3689] = 12'hbbf;
rom[3690] = 12'hbbf;
rom[3691] = 12'h99e;
rom[3692] = 12'h22d;
rom[3693] = 12'h  c;
rom[3694] = 12'h  c;
rom[3695] = 12'h  c;
rom[3696] = 12'h  c;
rom[3697] = 12'h  c;
rom[3698] = 12'h  c;
rom[3699] = 12'h  c;
rom[3700] = 12'h  c;
rom[3701] = 12'h  c;
rom[3702] = 12'h  c;
rom[3703] = 12'h22d;
rom[3704] = 12'hfff;
rom[3705] = 12'hfff;
rom[3706] = 12'hfff;
rom[3707] = 12'hfff;
rom[3708] = 12'hfff;
rom[3709] = 12'hfff;
rom[3710] = 12'hfff;
rom[3711] = 12'hfff;
rom[3712] = 12'hfff;
rom[3713] = 12'hfff;
rom[3714] = 12'hfff;
rom[3715] = 12'hfff;
rom[3716] = 12'hfff;
rom[3717] = 12'hfff;
rom[3718] = 12'hfff;
rom[3719] = 12'hfff;
rom[3720] = 12'hfff;
rom[3721] = 12'hfff;
rom[3722] = 12'hfff;
rom[3723] = 12'hfff;
rom[3724] = 12'hfff;
rom[3725] = 12'hfff;
rom[3726] = 12'hfff;
rom[3727] = 12'hfff;
rom[3728] = 12'hfff;
rom[3729] = 12'hfff;
rom[3730] = 12'hfff;
rom[3731] = 12'hfff;
rom[3732] = 12'hfff;
rom[3733] = 12'hfff;
rom[3734] = 12'hfff;
rom[3735] = 12'hfff;
rom[3736] = 12'hfff;
rom[3737] = 12'hfff;
rom[3738] = 12'hfff;
rom[3739] = 12'hfff;
rom[3740] = 12'hfff;
rom[3741] = 12'hfff;
rom[3742] = 12'hfff;
rom[3743] = 12'hfff;
rom[3744] = 12'hfff;
rom[3745] = 12'hfff;
rom[3746] = 12'hfff;
rom[3747] = 12'hfff;
rom[3748] = 12'hddf;
rom[3749] = 12'h88e;
rom[3750] = 12'h22d;
rom[3751] = 12'h  c;
rom[3752] = 12'h  c;
rom[3753] = 12'h  c;
rom[3754] = 12'h  c;
rom[3755] = 12'h  c;
rom[3756] = 12'h11d;
rom[3757] = 12'heef;
rom[3758] = 12'hfff;
rom[3759] = 12'hfff;
rom[3760] = 12'hfff;
rom[3761] = 12'hfff;
rom[3762] = 12'hfff;
rom[3763] = 12'hfff;
rom[3764] = 12'hfff;
rom[3765] = 12'hfff;
rom[3766] = 12'hfff;
rom[3767] = 12'hfff;
rom[3768] = 12'hfff;
rom[3769] = 12'hfff;
rom[3770] = 12'hfff;
rom[3771] = 12'hfff;
rom[3772] = 12'hfff;
rom[3773] = 12'hfff;
rom[3774] = 12'hfff;
rom[3775] = 12'hfff;
rom[3776] = 12'hfff;
rom[3777] = 12'hfff;
rom[3778] = 12'hfff;
rom[3779] = 12'hfff;
rom[3780] = 12'hfff;
rom[3781] = 12'hfff;
rom[3782] = 12'hfff;
rom[3783] = 12'hfff;
rom[3784] = 12'hfff;
rom[3785] = 12'hfff;
rom[3786] = 12'hfff;
rom[3787] = 12'hfff;
rom[3788] = 12'h22d;
rom[3789] = 12'h  c;
rom[3790] = 12'h  c;
rom[3791] = 12'h  c;
rom[3792] = 12'h  c;
rom[3793] = 12'h  c;
rom[3794] = 12'h  c;
rom[3795] = 12'h  c;
rom[3796] = 12'h  c;
rom[3797] = 12'h  c;
rom[3798] = 12'h33d;
rom[3799] = 12'h99e;
rom[3800] = 12'hbbf;
rom[3801] = 12'haae;
rom[3802] = 12'haae;
rom[3803] = 12'haae;
rom[3804] = 12'haae;
rom[3805] = 12'h99e;
rom[3806] = 12'h99e;
rom[3807] = 12'h88e;
rom[3808] = 12'h88e;
rom[3809] = 12'h99e;
rom[3810] = 12'heef;
rom[3811] = 12'hfff;
rom[3812] = 12'hfff;
rom[3813] = 12'hfff;
rom[3814] = 12'hfff;
rom[3815] = 12'hfff;
rom[3816] = 12'hfff;
rom[3817] = 12'hfff;
rom[3818] = 12'hfff;
rom[3819] = 12'hfff;
rom[3820] = 12'heef;
rom[3821] = 12'h88e;
rom[3822] = 12'h22d;
rom[3823] = 12'h  c;
rom[3824] = 12'h  c;
rom[3825] = 12'h  c;
rom[3826] = 12'h  c;
rom[3827] = 12'h  c;
rom[3828] = 12'h  c;
rom[3829] = 12'h  c;
rom[3830] = 12'h  c;
rom[3831] = 12'h  c;
rom[3832] = 12'h33d;
rom[3833] = 12'heef;
rom[3834] = 12'hfff;
rom[3835] = 12'hfff;
rom[3836] = 12'hfff;
rom[3837] = 12'hfff;
rom[3838] = 12'hfff;
rom[3839] = 12'hfff;
rom[3840] = 12'hfff;
rom[3841] = 12'hfff;
rom[3842] = 12'hfff;
rom[3843] = 12'hfff;
rom[3844] = 12'hfff;
rom[3845] = 12'hfff;
rom[3846] = 12'hfff;
rom[3847] = 12'hfff;
rom[3848] = 12'hfff;
rom[3849] = 12'hfff;
rom[3850] = 12'hfff;
rom[3851] = 12'hfff;
rom[3852] = 12'hfff;
rom[3853] = 12'hfff;
rom[3854] = 12'hfff;
rom[3855] = 12'hfff;
rom[3856] = 12'hfff;
rom[3857] = 12'hfff;
rom[3858] = 12'hfff;
rom[3859] = 12'hfff;
rom[3860] = 12'hfff;
rom[3861] = 12'hfff;
rom[3862] = 12'hfff;
rom[3863] = 12'hfff;
rom[3864] = 12'hfff;
rom[3865] = 12'hfff;
rom[3866] = 12'hfff;
rom[3867] = 12'hfff;
rom[3868] = 12'hfff;
rom[3869] = 12'hfff;
rom[3870] = 12'hfff;
rom[3871] = 12'hfff;
rom[3872] = 12'hfff;
rom[3873] = 12'hfff;
rom[3874] = 12'hfff;
rom[3875] = 12'hfff;
rom[3876] = 12'hfff;
rom[3877] = 12'heef;
rom[3878] = 12'h77e;
rom[3879] = 12'h11d;
rom[3880] = 12'h  c;
rom[3881] = 12'h  c;
rom[3882] = 12'h  c;
rom[3883] = 12'h  c;
rom[3884] = 12'h  c;
rom[3885] = 12'h22d;
rom[3886] = 12'hbbf;
rom[3887] = 12'heef;
rom[3888] = 12'hfff;
rom[3889] = 12'hfff;
rom[3890] = 12'hfff;
rom[3891] = 12'hfff;
rom[3892] = 12'hfff;
rom[3893] = 12'hfff;
rom[3894] = 12'hfff;
rom[3895] = 12'hfff;
rom[3896] = 12'hfff;
rom[3897] = 12'hfff;
rom[3898] = 12'hfff;
rom[3899] = 12'hfff;
rom[3900] = 12'hfff;
rom[3901] = 12'hfff;
rom[3902] = 12'hfff;
rom[3903] = 12'hfff;
rom[3904] = 12'hfff;
rom[3905] = 12'hfff;
rom[3906] = 12'hfff;
rom[3907] = 12'hfff;
rom[3908] = 12'hfff;
rom[3909] = 12'hfff;
rom[3910] = 12'hfff;
rom[3911] = 12'hfff;
rom[3912] = 12'hfff;
rom[3913] = 12'hfff;
rom[3914] = 12'hfff;
rom[3915] = 12'h77e;
rom[3916] = 12'h  c;
rom[3917] = 12'h  c;
rom[3918] = 12'h  c;
rom[3919] = 12'h  c;
rom[3920] = 12'h  c;
rom[3921] = 12'h  c;
rom[3922] = 12'h  c;
rom[3923] = 12'h33d;
rom[3924] = 12'h99e;
rom[3925] = 12'haae;
rom[3926] = 12'hfff;
rom[3927] = 12'hfff;
rom[3928] = 12'hfff;
rom[3929] = 12'hfff;
rom[3930] = 12'hfff;
rom[3931] = 12'hfff;
rom[3932] = 12'hfff;
rom[3933] = 12'hfff;
rom[3934] = 12'hfff;
rom[3935] = 12'hfff;
rom[3936] = 12'hfff;
rom[3937] = 12'hfff;
rom[3938] = 12'hfff;
rom[3939] = 12'hfff;
rom[3940] = 12'hfff;
rom[3941] = 12'hfff;
rom[3942] = 12'hfff;
rom[3943] = 12'hfff;
rom[3944] = 12'hfff;
rom[3945] = 12'hfff;
rom[3946] = 12'hfff;
rom[3947] = 12'hfff;
rom[3948] = 12'hfff;
rom[3949] = 12'hfff;
rom[3950] = 12'hfff;
rom[3951] = 12'haae;
rom[3952] = 12'haae;
rom[3953] = 12'h88e;
rom[3954] = 12'h33d;
rom[3955] = 12'h  c;
rom[3956] = 12'h  c;
rom[3957] = 12'h  c;
rom[3958] = 12'h  c;
rom[3959] = 12'h  c;
rom[3960] = 12'h  c;
rom[3961] = 12'h11d;
rom[3962] = 12'h77e;
rom[3963] = 12'heef;
rom[3964] = 12'hfff;
rom[3965] = 12'hfff;
rom[3966] = 12'hfff;
rom[3967] = 12'hfff;
rom[3968] = 12'hfff;
rom[3969] = 12'hfff;
rom[3970] = 12'hfff;
rom[3971] = 12'hfff;
rom[3972] = 12'hfff;
rom[3973] = 12'hfff;
rom[3974] = 12'hfff;
rom[3975] = 12'hfff;
rom[3976] = 12'hfff;
rom[3977] = 12'hfff;
rom[3978] = 12'hfff;
rom[3979] = 12'hfff;
rom[3980] = 12'hfff;
rom[3981] = 12'hfff;
rom[3982] = 12'hfff;
rom[3983] = 12'hfff;
rom[3984] = 12'hfff;
rom[3985] = 12'hfff;
rom[3986] = 12'hfff;
rom[3987] = 12'hfff;
rom[3988] = 12'hfff;
rom[3989] = 12'hfff;
rom[3990] = 12'hfff;
rom[3991] = 12'hfff;
rom[3992] = 12'hfff;
rom[3993] = 12'hfff;
rom[3994] = 12'hfff;
rom[3995] = 12'hfff;
rom[3996] = 12'hfff;
rom[3997] = 12'hfff;
rom[3998] = 12'hfff;
rom[3999] = 12'hfff;
rom[4000] = 12'hfff;
rom[4001] = 12'hfff;
rom[4002] = 12'hfff;
rom[4003] = 12'hfff;
rom[4004] = 12'hfff;
rom[4005] = 12'hfff;
rom[4006] = 12'hfff;
rom[4007] = 12'hddf;
rom[4008] = 12'h55d;
rom[4009] = 12'h11d;
rom[4010] = 12'h  c;
rom[4011] = 12'h  c;
rom[4012] = 12'h  c;
rom[4013] = 12'h  c;
rom[4014] = 12'h  c;
rom[4015] = 12'h11d;
rom[4016] = 12'haae;
rom[4017] = 12'hfff;
rom[4018] = 12'hfff;
rom[4019] = 12'hfff;
rom[4020] = 12'hfff;
rom[4021] = 12'hfff;
rom[4022] = 12'hfff;
rom[4023] = 12'hfff;
rom[4024] = 12'hfff;
rom[4025] = 12'hfff;
rom[4026] = 12'hfff;
rom[4027] = 12'hfff;
rom[4028] = 12'hfff;
rom[4029] = 12'hfff;
rom[4030] = 12'hfff;
rom[4031] = 12'hfff;
rom[4032] = 12'hfff;
rom[4033] = 12'hfff;
rom[4034] = 12'hfff;
rom[4035] = 12'hfff;
rom[4036] = 12'hfff;
rom[4037] = 12'hfff;
rom[4038] = 12'hfff;
rom[4039] = 12'hfff;
rom[4040] = 12'hfff;
rom[4041] = 12'hfff;
rom[4042] = 12'hddf;
rom[4043] = 12'h  c;
rom[4044] = 12'h  c;
rom[4045] = 12'h  c;
rom[4046] = 12'h  c;
rom[4047] = 12'h  c;
rom[4048] = 12'h  c;
rom[4049] = 12'h  c;
rom[4050] = 12'h55d;
rom[4051] = 12'hfff;
rom[4052] = 12'hfff;
rom[4053] = 12'hfff;
rom[4054] = 12'hfff;
rom[4055] = 12'hfff;
rom[4056] = 12'hfff;
rom[4057] = 12'hfff;
rom[4058] = 12'hfff;
rom[4059] = 12'hfff;
rom[4060] = 12'hfff;
rom[4061] = 12'hfff;
rom[4062] = 12'hfff;
rom[4063] = 12'hfff;
rom[4064] = 12'hfff;
rom[4065] = 12'hfff;
rom[4066] = 12'hfff;
rom[4067] = 12'hfff;
rom[4068] = 12'hfff;
rom[4069] = 12'hfff;
rom[4070] = 12'hfff;
rom[4071] = 12'hfff;
rom[4072] = 12'hfff;
rom[4073] = 12'hfff;
rom[4074] = 12'hfff;
rom[4075] = 12'hfff;
rom[4076] = 12'hfff;
rom[4077] = 12'hfff;
rom[4078] = 12'hfff;
rom[4079] = 12'hfff;
rom[4080] = 12'hfff;
rom[4081] = 12'hfff;
rom[4082] = 12'hfff;
rom[4083] = 12'h99e;
rom[4084] = 12'h11d;
rom[4085] = 12'h  c;
rom[4086] = 12'h  c;
rom[4087] = 12'h  c;
rom[4088] = 12'h  c;
rom[4089] = 12'h  c;
rom[4090] = 12'h  c;
rom[4091] = 12'h22d;
rom[4092] = 12'hfff;
rom[4093] = 12'hfff;
rom[4094] = 12'hfff;
rom[4095] = 12'hfff;
rom[4096] = 12'hfff;
rom[4097] = 12'hfff;
rom[4098] = 12'hfff;
rom[4099] = 12'hfff;
rom[4100] = 12'hfff;
rom[4101] = 12'hfff;
rom[4102] = 12'hfff;
rom[4103] = 12'hfff;
rom[4104] = 12'hfff;
rom[4105] = 12'hfff;
rom[4106] = 12'hfff;
rom[4107] = 12'hfff;
rom[4108] = 12'hfff;
rom[4109] = 12'hfff;
rom[4110] = 12'hfff;
rom[4111] = 12'hfff;
rom[4112] = 12'hfff;
rom[4113] = 12'hfff;
rom[4114] = 12'hfff;
rom[4115] = 12'hfff;
rom[4116] = 12'hfff;
rom[4117] = 12'hfff;
rom[4118] = 12'hfff;
rom[4119] = 12'hfff;
rom[4120] = 12'hfff;
rom[4121] = 12'hfff;
rom[4122] = 12'hfff;
rom[4123] = 12'hfff;
rom[4124] = 12'hfff;
rom[4125] = 12'hfff;
rom[4126] = 12'hfff;
rom[4127] = 12'hfff;
rom[4128] = 12'hfff;
rom[4129] = 12'hfff;
rom[4130] = 12'hfff;
rom[4131] = 12'hfff;
rom[4132] = 12'hfff;
rom[4133] = 12'hfff;
rom[4134] = 12'hfff;
rom[4135] = 12'hfff;
rom[4136] = 12'heef;
rom[4137] = 12'h11d;
rom[4138] = 12'h  c;
rom[4139] = 12'h  c;
rom[4140] = 12'h  c;
rom[4141] = 12'h  c;
rom[4142] = 12'h  c;
rom[4143] = 12'h  c;
rom[4144] = 12'h  c;
rom[4145] = 12'h88e;
rom[4146] = 12'hfff;
rom[4147] = 12'hfff;
rom[4148] = 12'hfff;
rom[4149] = 12'hfff;
rom[4150] = 12'hfff;
rom[4151] = 12'hfff;
rom[4152] = 12'hfff;
rom[4153] = 12'hfff;
rom[4154] = 12'hfff;
rom[4155] = 12'hfff;
rom[4156] = 12'hfff;
rom[4157] = 12'hfff;
rom[4158] = 12'hfff;
rom[4159] = 12'hfff;
rom[4160] = 12'hfff;
rom[4161] = 12'hfff;
rom[4162] = 12'hfff;
rom[4163] = 12'hfff;
rom[4164] = 12'hfff;
rom[4165] = 12'hfff;
rom[4166] = 12'hfff;
rom[4167] = 12'hfff;
rom[4168] = 12'hfff;
rom[4169] = 12'hfff;
rom[4170] = 12'h66e;
rom[4171] = 12'h  c;
rom[4172] = 12'h  c;
rom[4173] = 12'h  c;
rom[4174] = 12'h11d;
rom[4175] = 12'h33d;
rom[4176] = 12'h88e;
rom[4177] = 12'h99e;
rom[4178] = 12'hfff;
rom[4179] = 12'hfff;
rom[4180] = 12'hfff;
rom[4181] = 12'hfff;
rom[4182] = 12'hfff;
rom[4183] = 12'hfff;
rom[4184] = 12'hfff;
rom[4185] = 12'hfff;
rom[4186] = 12'hfff;
rom[4187] = 12'hfff;
rom[4188] = 12'hfff;
rom[4189] = 12'hfff;
rom[4190] = 12'hfff;
rom[4191] = 12'hfff;
rom[4192] = 12'hfff;
rom[4193] = 12'hfff;
rom[4194] = 12'hfff;
rom[4195] = 12'hfff;
rom[4196] = 12'hfff;
rom[4197] = 12'hfff;
rom[4198] = 12'hfff;
rom[4199] = 12'hfff;
rom[4200] = 12'hfff;
rom[4201] = 12'hfff;
rom[4202] = 12'hfff;
rom[4203] = 12'hfff;
rom[4204] = 12'hfff;
rom[4205] = 12'hfff;
rom[4206] = 12'hfff;
rom[4207] = 12'hfff;
rom[4208] = 12'hfff;
rom[4209] = 12'hfff;
rom[4210] = 12'hfff;
rom[4211] = 12'hfff;
rom[4212] = 12'heef;
rom[4213] = 12'h33d;
rom[4214] = 12'h  c;
rom[4215] = 12'h  c;
rom[4216] = 12'h  c;
rom[4217] = 12'h  c;
rom[4218] = 12'h  c;
rom[4219] = 12'h  c;
rom[4220] = 12'h99e;
rom[4221] = 12'hfff;
rom[4222] = 12'hfff;
rom[4223] = 12'hfff;
rom[4224] = 12'hfff;
rom[4225] = 12'hfff;
rom[4226] = 12'hfff;
rom[4227] = 12'hfff;
rom[4228] = 12'hfff;
rom[4229] = 12'hfff;
rom[4230] = 12'hfff;
rom[4231] = 12'hfff;
rom[4232] = 12'hfff;
rom[4233] = 12'hfff;
rom[4234] = 12'hfff;
rom[4235] = 12'hfff;
rom[4236] = 12'hfff;
rom[4237] = 12'hfff;
rom[4238] = 12'hfff;
rom[4239] = 12'hfff;
rom[4240] = 12'hfff;
rom[4241] = 12'hfff;
rom[4242] = 12'hfff;
rom[4243] = 12'hfff;
rom[4244] = 12'hfff;
rom[4245] = 12'hfff;
rom[4246] = 12'hfff;
rom[4247] = 12'hfff;
rom[4248] = 12'hfff;
rom[4249] = 12'hfff;
rom[4250] = 12'hfff;
rom[4251] = 12'hfff;
rom[4252] = 12'hfff;
rom[4253] = 12'hfff;
rom[4254] = 12'hfff;
rom[4255] = 12'hfff;
rom[4256] = 12'hfff;
rom[4257] = 12'hfff;
rom[4258] = 12'hfff;
rom[4259] = 12'hfff;
rom[4260] = 12'hfff;
rom[4261] = 12'hfff;
rom[4262] = 12'hfff;
rom[4263] = 12'hfff;
rom[4264] = 12'hfff;
rom[4265] = 12'hddf;
rom[4266] = 12'h  c;
rom[4267] = 12'h  c;
rom[4268] = 12'h  c;
rom[4269] = 12'h  c;
rom[4270] = 12'h  c;
rom[4271] = 12'h  c;
rom[4272] = 12'h  c;
rom[4273] = 12'h  c;
rom[4274] = 12'h77e;
rom[4275] = 12'hfff;
rom[4276] = 12'hfff;
rom[4277] = 12'hfff;
rom[4278] = 12'hfff;
rom[4279] = 12'hfff;
rom[4280] = 12'hfff;
rom[4281] = 12'hfff;
rom[4282] = 12'hfff;
rom[4283] = 12'hfff;
rom[4284] = 12'hfff;
rom[4285] = 12'hfff;
rom[4286] = 12'hfff;
rom[4287] = 12'hfff;
rom[4288] = 12'hfff;
rom[4289] = 12'hfff;
rom[4290] = 12'hfff;
rom[4291] = 12'hfff;
rom[4292] = 12'hfff;
rom[4293] = 12'hfff;
rom[4294] = 12'hfff;
rom[4295] = 12'hfff;
rom[4296] = 12'hfff;
rom[4297] = 12'heef;
rom[4298] = 12'h  c;
rom[4299] = 12'h  c;
rom[4300] = 12'h  c;
rom[4301] = 12'h  c;
rom[4302] = 12'h11d;
rom[4303] = 12'h99e;
rom[4304] = 12'hfff;
rom[4305] = 12'hfff;
rom[4306] = 12'hfff;
rom[4307] = 12'hfff;
rom[4308] = 12'hfff;
rom[4309] = 12'hfff;
rom[4310] = 12'hfff;
rom[4311] = 12'hfff;
rom[4312] = 12'hfff;
rom[4313] = 12'hfff;
rom[4314] = 12'hfff;
rom[4315] = 12'hfff;
rom[4316] = 12'hfff;
rom[4317] = 12'hfff;
rom[4318] = 12'hfff;
rom[4319] = 12'hfff;
rom[4320] = 12'hfff;
rom[4321] = 12'hfff;
rom[4322] = 12'hfff;
rom[4323] = 12'hfff;
rom[4324] = 12'hfff;
rom[4325] = 12'hfff;
rom[4326] = 12'hfff;
rom[4327] = 12'hfff;
rom[4328] = 12'hfff;
rom[4329] = 12'hfff;
rom[4330] = 12'hfff;
rom[4331] = 12'hfff;
rom[4332] = 12'hfff;
rom[4333] = 12'hfff;
rom[4334] = 12'hfff;
rom[4335] = 12'hfff;
rom[4336] = 12'hfff;
rom[4337] = 12'hfff;
rom[4338] = 12'hfff;
rom[4339] = 12'hfff;
rom[4340] = 12'hfff;
rom[4341] = 12'hfff;
rom[4342] = 12'h22d;
rom[4343] = 12'h  c;
rom[4344] = 12'h  c;
rom[4345] = 12'h  c;
rom[4346] = 12'h  c;
rom[4347] = 12'h  c;
rom[4348] = 12'h  c;
rom[4349] = 12'h77e;
rom[4350] = 12'hddf;
rom[4351] = 12'hfff;
rom[4352] = 12'hfff;
rom[4353] = 12'hfff;
rom[4354] = 12'hfff;
rom[4355] = 12'hfff;
rom[4356] = 12'hfff;
rom[4357] = 12'hfff;
rom[4358] = 12'hfff;
rom[4359] = 12'hfff;
rom[4360] = 12'hfff;
rom[4361] = 12'hfff;
rom[4362] = 12'hfff;
rom[4363] = 12'hfff;
rom[4364] = 12'hfff;
rom[4365] = 12'hfff;
rom[4366] = 12'hfff;
rom[4367] = 12'hfff;
rom[4368] = 12'hfff;
rom[4369] = 12'hfff;
rom[4370] = 12'hfff;
rom[4371] = 12'hfff;
rom[4372] = 12'hfff;
rom[4373] = 12'hfff;
rom[4374] = 12'hfff;
rom[4375] = 12'hfff;
rom[4376] = 12'hfff;
rom[4377] = 12'hfff;
rom[4378] = 12'hfff;
rom[4379] = 12'hfff;
rom[4380] = 12'hfff;
rom[4381] = 12'hfff;
rom[4382] = 12'hfff;
rom[4383] = 12'hfff;
rom[4384] = 12'hfff;
rom[4385] = 12'hfff;
rom[4386] = 12'hfff;
rom[4387] = 12'hfff;
rom[4388] = 12'hfff;
rom[4389] = 12'hfff;
rom[4390] = 12'hfff;
rom[4391] = 12'hfff;
rom[4392] = 12'hfff;
rom[4393] = 12'hfff;
rom[4394] = 12'hccf;
rom[4395] = 12'h33d;
rom[4396] = 12'h  c;
rom[4397] = 12'h  c;
rom[4398] = 12'h  c;
rom[4399] = 12'h  c;
rom[4400] = 12'h  c;
rom[4401] = 12'h  c;
rom[4402] = 12'h  c;
rom[4403] = 12'h88e;
rom[4404] = 12'hfff;
rom[4405] = 12'hfff;
rom[4406] = 12'hfff;
rom[4407] = 12'hfff;
rom[4408] = 12'hfff;
rom[4409] = 12'hfff;
rom[4410] = 12'hfff;
rom[4411] = 12'hfff;
rom[4412] = 12'hfff;
rom[4413] = 12'hfff;
rom[4414] = 12'hfff;
rom[4415] = 12'hfff;
rom[4416] = 12'hfff;
rom[4417] = 12'hfff;
rom[4418] = 12'hfff;
rom[4419] = 12'hfff;
rom[4420] = 12'hfff;
rom[4421] = 12'hfff;
rom[4422] = 12'hfff;
rom[4423] = 12'hfff;
rom[4424] = 12'hfff;
rom[4425] = 12'h88e;
rom[4426] = 12'h  c;
rom[4427] = 12'h  c;
rom[4428] = 12'h  c;
rom[4429] = 12'h  c;
rom[4430] = 12'h11d;
rom[4431] = 12'hfff;
rom[4432] = 12'hfff;
rom[4433] = 12'hfff;
rom[4434] = 12'hfff;
rom[4435] = 12'hfff;
rom[4436] = 12'hfff;
rom[4437] = 12'hfff;
rom[4438] = 12'hfff;
rom[4439] = 12'hfff;
rom[4440] = 12'hfff;
rom[4441] = 12'hfff;
rom[4442] = 12'hfff;
rom[4443] = 12'hfff;
rom[4444] = 12'hfff;
rom[4445] = 12'hfff;
rom[4446] = 12'hfff;
rom[4447] = 12'hfff;
rom[4448] = 12'hfff;
rom[4449] = 12'hfff;
rom[4450] = 12'hfff;
rom[4451] = 12'hfff;
rom[4452] = 12'hfff;
rom[4453] = 12'hfff;
rom[4454] = 12'hfff;
rom[4455] = 12'hfff;
rom[4456] = 12'hfff;
rom[4457] = 12'hfff;
rom[4458] = 12'hfff;
rom[4459] = 12'hfff;
rom[4460] = 12'hfff;
rom[4461] = 12'hfff;
rom[4462] = 12'hfff;
rom[4463] = 12'hfff;
rom[4464] = 12'hfff;
rom[4465] = 12'hfff;
rom[4466] = 12'hfff;
rom[4467] = 12'hfff;
rom[4468] = 12'hfff;
rom[4469] = 12'hfff;
rom[4470] = 12'hfff;
rom[4471] = 12'hbbf;
rom[4472] = 12'h  c;
rom[4473] = 12'h  c;
rom[4474] = 12'h  c;
rom[4475] = 12'h  c;
rom[4476] = 12'h  c;
rom[4477] = 12'h  c;
rom[4478] = 12'h  c;
rom[4479] = 12'hccf;
rom[4480] = 12'hfff;
rom[4481] = 12'hfff;
rom[4482] = 12'hfff;
rom[4483] = 12'hfff;
rom[4484] = 12'hfff;
rom[4485] = 12'hfff;
rom[4486] = 12'hfff;
rom[4487] = 12'hfff;
rom[4488] = 12'hfff;
rom[4489] = 12'hfff;
rom[4490] = 12'hfff;
rom[4491] = 12'hfff;
rom[4492] = 12'hfff;
rom[4493] = 12'hfff;
rom[4494] = 12'hfff;
rom[4495] = 12'hfff;
rom[4496] = 12'hfff;
rom[4497] = 12'hfff;
rom[4498] = 12'hfff;
rom[4499] = 12'hfff;
rom[4500] = 12'hfff;
rom[4501] = 12'hfff;
rom[4502] = 12'hfff;
rom[4503] = 12'hfff;
rom[4504] = 12'hfff;
rom[4505] = 12'hfff;
rom[4506] = 12'hfff;
rom[4507] = 12'hfff;
rom[4508] = 12'hfff;
rom[4509] = 12'hfff;
rom[4510] = 12'hfff;
rom[4511] = 12'hfff;
rom[4512] = 12'hfff;
rom[4513] = 12'hfff;
rom[4514] = 12'hfff;
rom[4515] = 12'hfff;
rom[4516] = 12'hfff;
rom[4517] = 12'hfff;
rom[4518] = 12'hfff;
rom[4519] = 12'hfff;
rom[4520] = 12'hfff;
rom[4521] = 12'hfff;
rom[4522] = 12'hfff;
rom[4523] = 12'hfff;
rom[4524] = 12'hddf;
rom[4525] = 12'h88e;
rom[4526] = 12'h22d;
rom[4527] = 12'h  c;
rom[4528] = 12'h  c;
rom[4529] = 12'h  c;
rom[4530] = 12'h  c;
rom[4531] = 12'h  c;
rom[4532] = 12'haae;
rom[4533] = 12'hfff;
rom[4534] = 12'hfff;
rom[4535] = 12'hfff;
rom[4536] = 12'hfff;
rom[4537] = 12'hfff;
rom[4538] = 12'hfff;
rom[4539] = 12'hfff;
rom[4540] = 12'hfff;
rom[4541] = 12'hfff;
rom[4542] = 12'hfff;
rom[4543] = 12'hfff;
rom[4544] = 12'hfff;
rom[4545] = 12'hfff;
rom[4546] = 12'hfff;
rom[4547] = 12'hfff;
rom[4548] = 12'hfff;
rom[4549] = 12'hfff;
rom[4550] = 12'hfff;
rom[4551] = 12'hfff;
rom[4552] = 12'hfff;
rom[4553] = 12'h33d;
rom[4554] = 12'h  c;
rom[4555] = 12'h  c;
rom[4556] = 12'h  c;
rom[4557] = 12'h  c;
rom[4558] = 12'h77e;
rom[4559] = 12'hfff;
rom[4560] = 12'hfff;
rom[4561] = 12'hfff;
rom[4562] = 12'hfff;
rom[4563] = 12'hfff;
rom[4564] = 12'hfff;
rom[4565] = 12'hfff;
rom[4566] = 12'hfff;
rom[4567] = 12'hfff;
rom[4568] = 12'hfff;
rom[4569] = 12'hfff;
rom[4570] = 12'hfff;
rom[4571] = 12'hfff;
rom[4572] = 12'hfff;
rom[4573] = 12'hfff;
rom[4574] = 12'hfff;
rom[4575] = 12'hfff;
rom[4576] = 12'hfff;
rom[4577] = 12'hfff;
rom[4578] = 12'hfff;
rom[4579] = 12'hfff;
rom[4580] = 12'hfff;
rom[4581] = 12'hfff;
rom[4582] = 12'hfff;
rom[4583] = 12'hfff;
rom[4584] = 12'hfff;
rom[4585] = 12'hfff;
rom[4586] = 12'hfff;
rom[4587] = 12'hfff;
rom[4588] = 12'hfff;
rom[4589] = 12'hfff;
rom[4590] = 12'hfff;
rom[4591] = 12'hfff;
rom[4592] = 12'hfff;
rom[4593] = 12'hfff;
rom[4594] = 12'hfff;
rom[4595] = 12'hfff;
rom[4596] = 12'hfff;
rom[4597] = 12'hfff;
rom[4598] = 12'hfff;
rom[4599] = 12'hfff;
rom[4600] = 12'h66e;
rom[4601] = 12'h  c;
rom[4602] = 12'h  c;
rom[4603] = 12'h  c;
rom[4604] = 12'h  c;
rom[4605] = 12'h  c;
rom[4606] = 12'h  c;
rom[4607] = 12'h11d;
rom[4608] = 12'hfff;
rom[4609] = 12'hfff;
rom[4610] = 12'hfff;
rom[4611] = 12'hfff;
rom[4612] = 12'hfff;
rom[4613] = 12'hfff;
rom[4614] = 12'hfff;
rom[4615] = 12'hfff;
rom[4616] = 12'hfff;
rom[4617] = 12'hfff;
rom[4618] = 12'hfff;
rom[4619] = 12'hfff;
rom[4620] = 12'hfff;
rom[4621] = 12'hfff;
rom[4622] = 12'hfff;
rom[4623] = 12'hfff;
rom[4624] = 12'hfff;
rom[4625] = 12'hfff;
rom[4626] = 12'hfff;
rom[4627] = 12'hfff;
rom[4628] = 12'hfff;
rom[4629] = 12'hfff;
rom[4630] = 12'hfff;
rom[4631] = 12'hfff;
rom[4632] = 12'hfff;
rom[4633] = 12'hfff;
rom[4634] = 12'hfff;
rom[4635] = 12'hfff;
rom[4636] = 12'hfff;
rom[4637] = 12'hfff;
rom[4638] = 12'hfff;
rom[4639] = 12'hfff;
rom[4640] = 12'hfff;
rom[4641] = 12'hfff;
rom[4642] = 12'hfff;
rom[4643] = 12'hfff;
rom[4644] = 12'hfff;
rom[4645] = 12'hfff;
rom[4646] = 12'hfff;
rom[4647] = 12'hfff;
rom[4648] = 12'hfff;
rom[4649] = 12'hfff;
rom[4650] = 12'hfff;
rom[4651] = 12'hfff;
rom[4652] = 12'hfff;
rom[4653] = 12'hfff;
rom[4654] = 12'h77e;
rom[4655] = 12'h  c;
rom[4656] = 12'h  c;
rom[4657] = 12'h  c;
rom[4658] = 12'h  c;
rom[4659] = 12'h  c;
rom[4660] = 12'h22d;
rom[4661] = 12'hfff;
rom[4662] = 12'hfff;
rom[4663] = 12'hfff;
rom[4664] = 12'hfff;
rom[4665] = 12'hfff;
rom[4666] = 12'hfff;
rom[4667] = 12'hfff;
rom[4668] = 12'hfff;
rom[4669] = 12'hfff;
rom[4670] = 12'hfff;
rom[4671] = 12'hfff;
rom[4672] = 12'hfff;
rom[4673] = 12'hfff;
rom[4674] = 12'hfff;
rom[4675] = 12'hfff;
rom[4676] = 12'hfff;
rom[4677] = 12'hfff;
rom[4678] = 12'hfff;
rom[4679] = 12'hfff;
rom[4680] = 12'hfff;
rom[4681] = 12'h11d;
rom[4682] = 12'h  c;
rom[4683] = 12'h  c;
rom[4684] = 12'h  c;
rom[4685] = 12'h  c;
rom[4686] = 12'hddf;
rom[4687] = 12'hfff;
rom[4688] = 12'hfff;
rom[4689] = 12'hfff;
rom[4690] = 12'hfff;
rom[4691] = 12'hfff;
rom[4692] = 12'hfff;
rom[4693] = 12'hfff;
rom[4694] = 12'hfff;
rom[4695] = 12'hfff;
rom[4696] = 12'hfff;
rom[4697] = 12'hfff;
rom[4698] = 12'hfff;
rom[4699] = 12'hfff;
rom[4700] = 12'hfff;
rom[4701] = 12'hfff;
rom[4702] = 12'hfff;
rom[4703] = 12'hfff;
rom[4704] = 12'hfff;
rom[4705] = 12'hfff;
rom[4706] = 12'hfff;
rom[4707] = 12'hfff;
rom[4708] = 12'hfff;
rom[4709] = 12'hfff;
rom[4710] = 12'hfff;
rom[4711] = 12'hfff;
rom[4712] = 12'hfff;
rom[4713] = 12'hfff;
rom[4714] = 12'hfff;
rom[4715] = 12'hfff;
rom[4716] = 12'hfff;
rom[4717] = 12'hfff;
rom[4718] = 12'hfff;
rom[4719] = 12'hfff;
rom[4720] = 12'hfff;
rom[4721] = 12'hfff;
rom[4722] = 12'hfff;
rom[4723] = 12'hfff;
rom[4724] = 12'hfff;
rom[4725] = 12'hfff;
rom[4726] = 12'hfff;
rom[4727] = 12'hfff;
rom[4728] = 12'heef;
rom[4729] = 12'h22d;
rom[4730] = 12'h  c;
rom[4731] = 12'h22d;
rom[4732] = 12'h  c;
rom[4733] = 12'h  c;
rom[4734] = 12'h  c;
rom[4735] = 12'h  c;
rom[4736] = 12'hfff;
rom[4737] = 12'hfff;
rom[4738] = 12'hfff;
rom[4739] = 12'hfff;
rom[4740] = 12'hfff;
rom[4741] = 12'hfff;
rom[4742] = 12'hfff;
rom[4743] = 12'hfff;
rom[4744] = 12'hfff;
rom[4745] = 12'hfff;
rom[4746] = 12'hfff;
rom[4747] = 12'hfff;
rom[4748] = 12'hfff;
rom[4749] = 12'hfff;
rom[4750] = 12'hfff;
rom[4751] = 12'hfff;
rom[4752] = 12'hfff;
rom[4753] = 12'hfff;
rom[4754] = 12'hfff;
rom[4755] = 12'hfff;
rom[4756] = 12'hfff;
rom[4757] = 12'hfff;
rom[4758] = 12'hfff;
rom[4759] = 12'hfff;
rom[4760] = 12'hfff;
rom[4761] = 12'hfff;
rom[4762] = 12'hfff;
rom[4763] = 12'hfff;
rom[4764] = 12'hfff;
rom[4765] = 12'hfff;
rom[4766] = 12'hfff;
rom[4767] = 12'hfff;
rom[4768] = 12'hfff;
rom[4769] = 12'hfff;
rom[4770] = 12'hfff;
rom[4771] = 12'hfff;
rom[4772] = 12'hfff;
rom[4773] = 12'hfff;
rom[4774] = 12'hfff;
rom[4775] = 12'hfff;
rom[4776] = 12'hfff;
rom[4777] = 12'hfff;
rom[4778] = 12'hfff;
rom[4779] = 12'hfff;
rom[4780] = 12'hfff;
rom[4781] = 12'hfff;
rom[4782] = 12'hfff;
rom[4783] = 12'h77e;
rom[4784] = 12'h  c;
rom[4785] = 12'h  c;
rom[4786] = 12'h  c;
rom[4787] = 12'h  c;
rom[4788] = 12'h  c;
rom[4789] = 12'h99e;
rom[4790] = 12'hfff;
rom[4791] = 12'hfff;
rom[4792] = 12'hfff;
rom[4793] = 12'hfff;
rom[4794] = 12'hfff;
rom[4795] = 12'hfff;
rom[4796] = 12'hfff;
rom[4797] = 12'hfff;
rom[4798] = 12'hfff;
rom[4799] = 12'hfff;
rom[4800] = 12'hfff;
rom[4801] = 12'hfff;
rom[4802] = 12'hfff;
rom[4803] = 12'hfff;
rom[4804] = 12'hfff;
rom[4805] = 12'hfff;
rom[4806] = 12'hfff;
rom[4807] = 12'heef;
rom[4808] = 12'h33d;
rom[4809] = 12'h  c;
rom[4810] = 12'h  c;
rom[4811] = 12'h  c;
rom[4812] = 12'h  c;
rom[4813] = 12'h33d;
rom[4814] = 12'hfff;
rom[4815] = 12'hfff;
rom[4816] = 12'hfff;
rom[4817] = 12'hfff;
rom[4818] = 12'hfff;
rom[4819] = 12'hfff;
rom[4820] = 12'hfff;
rom[4821] = 12'hfff;
rom[4822] = 12'hfff;
rom[4823] = 12'hfff;
rom[4824] = 12'hfff;
rom[4825] = 12'hfff;
rom[4826] = 12'hfff;
rom[4827] = 12'hfff;
rom[4828] = 12'hfff;
rom[4829] = 12'hfff;
rom[4830] = 12'hfff;
rom[4831] = 12'hfff;
rom[4832] = 12'hfff;
rom[4833] = 12'hfff;
rom[4834] = 12'hfff;
rom[4835] = 12'hfff;
rom[4836] = 12'hfff;
rom[4837] = 12'hfff;
rom[4838] = 12'hfff;
rom[4839] = 12'hfff;
rom[4840] = 12'hfff;
rom[4841] = 12'hfff;
rom[4842] = 12'hfff;
rom[4843] = 12'hfff;
rom[4844] = 12'hfff;
rom[4845] = 12'hfff;
rom[4846] = 12'hfff;
rom[4847] = 12'hfff;
rom[4848] = 12'hfff;
rom[4849] = 12'hfff;
rom[4850] = 12'hfff;
rom[4851] = 12'hfff;
rom[4852] = 12'hfff;
rom[4853] = 12'hfff;
rom[4854] = 12'hfff;
rom[4855] = 12'hfff;
rom[4856] = 12'hfff;
rom[4857] = 12'heef;
rom[4858] = 12'haae;
rom[4859] = 12'h66e;
rom[4860] = 12'h  c;
rom[4861] = 12'h  c;
rom[4862] = 12'h  c;
rom[4863] = 12'h  c;
rom[4864] = 12'hfff;
rom[4865] = 12'hfff;
rom[4866] = 12'hfff;
rom[4867] = 12'hfff;
rom[4868] = 12'hfff;
rom[4869] = 12'hfff;
rom[4870] = 12'hfff;
rom[4871] = 12'hfff;
rom[4872] = 12'hfff;
rom[4873] = 12'hfff;
rom[4874] = 12'hfff;
rom[4875] = 12'hfff;
rom[4876] = 12'hfff;
rom[4877] = 12'hfff;
rom[4878] = 12'hfff;
rom[4879] = 12'hfff;
rom[4880] = 12'hfff;
rom[4881] = 12'hfff;
rom[4882] = 12'hfff;
rom[4883] = 12'hfff;
rom[4884] = 12'hfff;
rom[4885] = 12'hfff;
rom[4886] = 12'hfff;
rom[4887] = 12'hfff;
rom[4888] = 12'hfff;
rom[4889] = 12'hfff;
rom[4890] = 12'hfff;
rom[4891] = 12'hfff;
rom[4892] = 12'hfff;
rom[4893] = 12'hfff;
rom[4894] = 12'hfff;
rom[4895] = 12'hfff;
rom[4896] = 12'hfff;
rom[4897] = 12'hfff;
rom[4898] = 12'hfff;
rom[4899] = 12'hfff;
rom[4900] = 12'hfff;
rom[4901] = 12'hfff;
rom[4902] = 12'hfff;
rom[4903] = 12'hfff;
rom[4904] = 12'hfff;
rom[4905] = 12'hfff;
rom[4906] = 12'hfff;
rom[4907] = 12'hfff;
rom[4908] = 12'hfff;
rom[4909] = 12'hfff;
rom[4910] = 12'hfff;
rom[4911] = 12'hfff;
rom[4912] = 12'h55d;
rom[4913] = 12'h  c;
rom[4914] = 12'h  c;
rom[4915] = 12'h  c;
rom[4916] = 12'h  c;
rom[4917] = 12'h88e;
rom[4918] = 12'hfff;
rom[4919] = 12'hfff;
rom[4920] = 12'hfff;
rom[4921] = 12'hfff;
rom[4922] = 12'hfff;
rom[4923] = 12'hfff;
rom[4924] = 12'hfff;
rom[4925] = 12'hfff;
rom[4926] = 12'hfff;
rom[4927] = 12'hfff;
rom[4928] = 12'hfff;
rom[4929] = 12'hfff;
rom[4930] = 12'hfff;
rom[4931] = 12'hfff;
rom[4932] = 12'hfff;
rom[4933] = 12'hfff;
rom[4934] = 12'hfff;
rom[4935] = 12'h99e;
rom[4936] = 12'h  c;
rom[4937] = 12'h  c;
rom[4938] = 12'h  c;
rom[4939] = 12'h  c;
rom[4940] = 12'h  c;
rom[4941] = 12'haae;
rom[4942] = 12'hfff;
rom[4943] = 12'hfff;
rom[4944] = 12'hfff;
rom[4945] = 12'hfff;
rom[4946] = 12'hfff;
rom[4947] = 12'hfff;
rom[4948] = 12'hfff;
rom[4949] = 12'hfff;
rom[4950] = 12'hfff;
rom[4951] = 12'hfff;
rom[4952] = 12'hfff;
rom[4953] = 12'hfff;
rom[4954] = 12'hfff;
rom[4955] = 12'hfff;
rom[4956] = 12'hfff;
rom[4957] = 12'hfff;
rom[4958] = 12'hfff;
rom[4959] = 12'hfff;
rom[4960] = 12'hfff;
rom[4961] = 12'hfff;
rom[4962] = 12'hfff;
rom[4963] = 12'hfff;
rom[4964] = 12'hfff;
rom[4965] = 12'hfff;
rom[4966] = 12'hfff;
rom[4967] = 12'hfff;
rom[4968] = 12'hfff;
rom[4969] = 12'hfff;
rom[4970] = 12'hfff;
rom[4971] = 12'hfff;
rom[4972] = 12'hfff;
rom[4973] = 12'hfff;
rom[4974] = 12'hfff;
rom[4975] = 12'hfff;
rom[4976] = 12'hfff;
rom[4977] = 12'hfff;
rom[4978] = 12'hfff;
rom[4979] = 12'hfff;
rom[4980] = 12'hfff;
rom[4981] = 12'hfff;
rom[4982] = 12'hfff;
rom[4983] = 12'hfff;
rom[4984] = 12'hfff;
rom[4985] = 12'hfff;
rom[4986] = 12'hfff;
rom[4987] = 12'hccf;
rom[4988] = 12'h  c;
rom[4989] = 12'h  c;
rom[4990] = 12'h  c;
rom[4991] = 12'h  c;
rom[4992] = 12'hfff;
rom[4993] = 12'hfff;
rom[4994] = 12'hfff;
rom[4995] = 12'hfff;
rom[4996] = 12'hfff;
rom[4997] = 12'hfff;
rom[4998] = 12'hfff;
rom[4999] = 12'hfff;
rom[5000] = 12'hfff;
rom[5001] = 12'hfff;
rom[5002] = 12'hfff;
rom[5003] = 12'hfff;
rom[5004] = 12'hfff;
rom[5005] = 12'hfff;
rom[5006] = 12'hfff;
rom[5007] = 12'hfff;
rom[5008] = 12'hfff;
rom[5009] = 12'hfff;
rom[5010] = 12'hfff;
rom[5011] = 12'hfff;
rom[5012] = 12'hfff;
rom[5013] = 12'hfff;
rom[5014] = 12'hfff;
rom[5015] = 12'hfff;
rom[5016] = 12'hfff;
rom[5017] = 12'hfff;
rom[5018] = 12'hfff;
rom[5019] = 12'hfff;
rom[5020] = 12'hfff;
rom[5021] = 12'hfff;
rom[5022] = 12'hfff;
rom[5023] = 12'hfff;
rom[5024] = 12'hfff;
rom[5025] = 12'hfff;
rom[5026] = 12'hfff;
rom[5027] = 12'hfff;
rom[5028] = 12'hfff;
rom[5029] = 12'hfff;
rom[5030] = 12'hfff;
rom[5031] = 12'hfff;
rom[5032] = 12'hfff;
rom[5033] = 12'hfff;
rom[5034] = 12'hfff;
rom[5035] = 12'hfff;
rom[5036] = 12'hfff;
rom[5037] = 12'hfff;
rom[5038] = 12'hfff;
rom[5039] = 12'hfff;
rom[5040] = 12'hbbf;
rom[5041] = 12'h11d;
rom[5042] = 12'h  c;
rom[5043] = 12'h  c;
rom[5044] = 12'h  c;
rom[5045] = 12'h44d;
rom[5046] = 12'heef;
rom[5047] = 12'hfff;
rom[5048] = 12'hfff;
rom[5049] = 12'hfff;
rom[5050] = 12'hfff;
rom[5051] = 12'hfff;
rom[5052] = 12'hfff;
rom[5053] = 12'hfff;
rom[5054] = 12'hfff;
rom[5055] = 12'hfff;
rom[5056] = 12'hfff;
rom[5057] = 12'hfff;
rom[5058] = 12'hfff;
rom[5059] = 12'hfff;
rom[5060] = 12'hfff;
rom[5061] = 12'hfff;
rom[5062] = 12'hfff;
rom[5063] = 12'h77e;
rom[5064] = 12'h  c;
rom[5065] = 12'h  c;
rom[5066] = 12'h  c;
rom[5067] = 12'h  c;
rom[5068] = 12'h33d;
rom[5069] = 12'hfff;
rom[5070] = 12'hfff;
rom[5071] = 12'hfff;
rom[5072] = 12'hfff;
rom[5073] = 12'hfff;
rom[5074] = 12'hfff;
rom[5075] = 12'hfff;
rom[5076] = 12'hfff;
rom[5077] = 12'hfff;
rom[5078] = 12'hfff;
rom[5079] = 12'hfff;
rom[5080] = 12'hfff;
rom[5081] = 12'hfff;
rom[5082] = 12'hfff;
rom[5083] = 12'hfff;
rom[5084] = 12'hfff;
rom[5085] = 12'hfff;
rom[5086] = 12'hfff;
rom[5087] = 12'hfff;
rom[5088] = 12'hfff;
rom[5089] = 12'hfff;
rom[5090] = 12'hfff;
rom[5091] = 12'hfff;
rom[5092] = 12'hfff;
rom[5093] = 12'hfff;
rom[5094] = 12'hfff;
rom[5095] = 12'hfff;
rom[5096] = 12'hfff;
rom[5097] = 12'hfff;
rom[5098] = 12'hfff;
rom[5099] = 12'hfff;
rom[5100] = 12'hfff;
rom[5101] = 12'hfff;
rom[5102] = 12'hfff;
rom[5103] = 12'hfff;
rom[5104] = 12'hfff;
rom[5105] = 12'hfff;
rom[5106] = 12'hfff;
rom[5107] = 12'hfff;
rom[5108] = 12'hfff;
rom[5109] = 12'hfff;
rom[5110] = 12'hfff;
rom[5111] = 12'hfff;
rom[5112] = 12'hfff;
rom[5113] = 12'hfff;
rom[5114] = 12'hfff;
rom[5115] = 12'hfff;
rom[5116] = 12'h66e;
rom[5117] = 12'h  c;
rom[5118] = 12'h  c;
rom[5119] = 12'h  c;
rom[5120] = 12'hfff;
rom[5121] = 12'hfff;
rom[5122] = 12'hfff;
rom[5123] = 12'hfff;
rom[5124] = 12'hfff;
rom[5125] = 12'hfff;
rom[5126] = 12'hfff;
rom[5127] = 12'hfff;
rom[5128] = 12'hfff;
rom[5129] = 12'hfff;
rom[5130] = 12'hfff;
rom[5131] = 12'hfff;
rom[5132] = 12'hfff;
rom[5133] = 12'hfff;
rom[5134] = 12'hfff;
rom[5135] = 12'hfff;
rom[5136] = 12'hfff;
rom[5137] = 12'hfff;
rom[5138] = 12'hfff;
rom[5139] = 12'hfff;
rom[5140] = 12'hfff;
rom[5141] = 12'hfff;
rom[5142] = 12'hfff;
rom[5143] = 12'hfff;
rom[5144] = 12'hfff;
rom[5145] = 12'hfff;
rom[5146] = 12'hfff;
rom[5147] = 12'hfff;
rom[5148] = 12'hfff;
rom[5149] = 12'hfff;
rom[5150] = 12'hfff;
rom[5151] = 12'hfff;
rom[5152] = 12'hfff;
rom[5153] = 12'hfff;
rom[5154] = 12'hfff;
rom[5155] = 12'hfff;
rom[5156] = 12'hfff;
rom[5157] = 12'hfff;
rom[5158] = 12'hfff;
rom[5159] = 12'hfff;
rom[5160] = 12'hfff;
rom[5161] = 12'hfff;
rom[5162] = 12'hfff;
rom[5163] = 12'hfff;
rom[5164] = 12'hfff;
rom[5165] = 12'hfff;
rom[5166] = 12'hfff;
rom[5167] = 12'hfff;
rom[5168] = 12'h99e;
rom[5169] = 12'h  c;
rom[5170] = 12'h  c;
rom[5171] = 12'h  c;
rom[5172] = 12'h  c;
rom[5173] = 12'h11d;
rom[5174] = 12'h22d;
rom[5175] = 12'heef;
rom[5176] = 12'hfff;
rom[5177] = 12'hfff;
rom[5178] = 12'hfff;
rom[5179] = 12'hfff;
rom[5180] = 12'hfff;
rom[5181] = 12'hfff;
rom[5182] = 12'hfff;
rom[5183] = 12'hfff;
rom[5184] = 12'hfff;
rom[5185] = 12'hfff;
rom[5186] = 12'hfff;
rom[5187] = 12'hfff;
rom[5188] = 12'hfff;
rom[5189] = 12'hfff;
rom[5190] = 12'hfff;
rom[5191] = 12'h77e;
rom[5192] = 12'h  c;
rom[5193] = 12'h  c;
rom[5194] = 12'h  c;
rom[5195] = 12'h11d;
rom[5196] = 12'h88e;
rom[5197] = 12'hfff;
rom[5198] = 12'hfff;
rom[5199] = 12'hfff;
rom[5200] = 12'hfff;
rom[5201] = 12'hfff;
rom[5202] = 12'hfff;
rom[5203] = 12'hfff;
rom[5204] = 12'hfff;
rom[5205] = 12'hfff;
rom[5206] = 12'hfff;
rom[5207] = 12'hfff;
rom[5208] = 12'hfff;
rom[5209] = 12'hfff;
rom[5210] = 12'hfff;
rom[5211] = 12'hfff;
rom[5212] = 12'hfff;
rom[5213] = 12'hfff;
rom[5214] = 12'hfff;
rom[5215] = 12'hfff;
rom[5216] = 12'hfff;
rom[5217] = 12'hfff;
rom[5218] = 12'hfff;
rom[5219] = 12'hfff;
rom[5220] = 12'hfff;
rom[5221] = 12'hfff;
rom[5222] = 12'hfff;
rom[5223] = 12'hfff;
rom[5224] = 12'hfff;
rom[5225] = 12'hfff;
rom[5226] = 12'hfff;
rom[5227] = 12'hfff;
rom[5228] = 12'hfff;
rom[5229] = 12'hfff;
rom[5230] = 12'hfff;
rom[5231] = 12'hfff;
rom[5232] = 12'hfff;
rom[5233] = 12'hfff;
rom[5234] = 12'hfff;
rom[5235] = 12'hfff;
rom[5236] = 12'hfff;
rom[5237] = 12'hfff;
rom[5238] = 12'hfff;
rom[5239] = 12'hfff;
rom[5240] = 12'hfff;
rom[5241] = 12'hfff;
rom[5242] = 12'hfff;
rom[5243] = 12'hfff;
rom[5244] = 12'heef;
rom[5245] = 12'h11d;
rom[5246] = 12'h  c;
rom[5247] = 12'h  c;
rom[5248] = 12'hfff;
rom[5249] = 12'hfff;
rom[5250] = 12'hfff;
rom[5251] = 12'hfff;
rom[5252] = 12'hfff;
rom[5253] = 12'hfff;
rom[5254] = 12'hfff;
rom[5255] = 12'hfff;
rom[5256] = 12'hfff;
rom[5257] = 12'hfff;
rom[5258] = 12'hfff;
rom[5259] = 12'hfff;
rom[5260] = 12'hfff;
rom[5261] = 12'hfff;
rom[5262] = 12'hfff;
rom[5263] = 12'hfff;
rom[5264] = 12'hfff;
rom[5265] = 12'hfff;
rom[5266] = 12'hfff;
rom[5267] = 12'hfff;
rom[5268] = 12'hfff;
rom[5269] = 12'hfff;
rom[5270] = 12'hfff;
rom[5271] = 12'hfff;
rom[5272] = 12'hfff;
rom[5273] = 12'hfff;
rom[5274] = 12'hfff;
rom[5275] = 12'hfff;
rom[5276] = 12'hfff;
rom[5277] = 12'hfff;
rom[5278] = 12'hfff;
rom[5279] = 12'hfff;
rom[5280] = 12'hfff;
rom[5281] = 12'hfff;
rom[5282] = 12'hfff;
rom[5283] = 12'hfff;
rom[5284] = 12'hfff;
rom[5285] = 12'hfff;
rom[5286] = 12'hfff;
rom[5287] = 12'hfff;
rom[5288] = 12'hfff;
rom[5289] = 12'hfff;
rom[5290] = 12'hfff;
rom[5291] = 12'hfff;
rom[5292] = 12'hfff;
rom[5293] = 12'hfff;
rom[5294] = 12'hfff;
rom[5295] = 12'hfff;
rom[5296] = 12'heef;
rom[5297] = 12'h11d;
rom[5298] = 12'h  c;
rom[5299] = 12'h  c;
rom[5300] = 12'h  c;
rom[5301] = 12'h  c;
rom[5302] = 12'h  c;
rom[5303] = 12'h33d;
rom[5304] = 12'heef;
rom[5305] = 12'hfff;
rom[5306] = 12'hfff;
rom[5307] = 12'hfff;
rom[5308] = 12'hfff;
rom[5309] = 12'hfff;
rom[5310] = 12'hfff;
rom[5311] = 12'hfff;
rom[5312] = 12'hfff;
rom[5313] = 12'hfff;
rom[5314] = 12'hfff;
rom[5315] = 12'hfff;
rom[5316] = 12'hfff;
rom[5317] = 12'hfff;
rom[5318] = 12'hfff;
rom[5319] = 12'h88e;
rom[5320] = 12'h  c;
rom[5321] = 12'h  c;
rom[5322] = 12'h  c;
rom[5323] = 12'h  c;
rom[5324] = 12'h77e;
rom[5325] = 12'hfff;
rom[5326] = 12'hfff;
rom[5327] = 12'hfff;
rom[5328] = 12'hfff;
rom[5329] = 12'hfff;
rom[5330] = 12'hfff;
rom[5331] = 12'hfff;
rom[5332] = 12'hfff;
rom[5333] = 12'hfff;
rom[5334] = 12'hfff;
rom[5335] = 12'hfff;
rom[5336] = 12'hfff;
rom[5337] = 12'hfff;
rom[5338] = 12'hfff;
rom[5339] = 12'hfff;
rom[5340] = 12'hfff;
rom[5341] = 12'hfff;
rom[5342] = 12'hfff;
rom[5343] = 12'hfff;
rom[5344] = 12'hfff;
rom[5345] = 12'hfff;
rom[5346] = 12'hfff;
rom[5347] = 12'hfff;
rom[5348] = 12'hfff;
rom[5349] = 12'hfff;
rom[5350] = 12'hfff;
rom[5351] = 12'hfff;
rom[5352] = 12'hfff;
rom[5353] = 12'hfff;
rom[5354] = 12'hfff;
rom[5355] = 12'hfff;
rom[5356] = 12'hfff;
rom[5357] = 12'hfff;
rom[5358] = 12'hfff;
rom[5359] = 12'hfff;
rom[5360] = 12'hfff;
rom[5361] = 12'hfff;
rom[5362] = 12'hfff;
rom[5363] = 12'hfff;
rom[5364] = 12'hfff;
rom[5365] = 12'hfff;
rom[5366] = 12'hfff;
rom[5367] = 12'hfff;
rom[5368] = 12'hfff;
rom[5369] = 12'hfff;
rom[5370] = 12'hfff;
rom[5371] = 12'hfff;
rom[5372] = 12'hfff;
rom[5373] = 12'heef;
rom[5374] = 12'hccf;
rom[5375] = 12'h44d;
rom[5376] = 12'hfff;
rom[5377] = 12'hfff;
rom[5378] = 12'hfff;
rom[5379] = 12'hfff;
rom[5380] = 12'hfff;
rom[5381] = 12'hfff;
rom[5382] = 12'hfff;
rom[5383] = 12'hfff;
rom[5384] = 12'hfff;
rom[5385] = 12'hfff;
rom[5386] = 12'hfff;
rom[5387] = 12'hfff;
rom[5388] = 12'hfff;
rom[5389] = 12'hfff;
rom[5390] = 12'hfff;
rom[5391] = 12'hfff;
rom[5392] = 12'hfff;
rom[5393] = 12'hfff;
rom[5394] = 12'hfff;
rom[5395] = 12'hfff;
rom[5396] = 12'hfff;
rom[5397] = 12'hfff;
rom[5398] = 12'hfff;
rom[5399] = 12'hfff;
rom[5400] = 12'hfff;
rom[5401] = 12'hfff;
rom[5402] = 12'hfff;
rom[5403] = 12'hfff;
rom[5404] = 12'hfff;
rom[5405] = 12'hfff;
rom[5406] = 12'hfff;
rom[5407] = 12'hfff;
rom[5408] = 12'hfff;
rom[5409] = 12'hfff;
rom[5410] = 12'hfff;
rom[5411] = 12'hfff;
rom[5412] = 12'hfff;
rom[5413] = 12'hfff;
rom[5414] = 12'hfff;
rom[5415] = 12'hfff;
rom[5416] = 12'hfff;
rom[5417] = 12'hfff;
rom[5418] = 12'hfff;
rom[5419] = 12'hfff;
rom[5420] = 12'hfff;
rom[5421] = 12'hfff;
rom[5422] = 12'hfff;
rom[5423] = 12'hfff;
rom[5424] = 12'hfff;
rom[5425] = 12'hccf;
rom[5426] = 12'h  c;
rom[5427] = 12'h  c;
rom[5428] = 12'h  c;
rom[5429] = 12'h  c;
rom[5430] = 12'h  c;
rom[5431] = 12'h  c;
rom[5432] = 12'h22d;
rom[5433] = 12'hfff;
rom[5434] = 12'hfff;
rom[5435] = 12'hfff;
rom[5436] = 12'hfff;
rom[5437] = 12'hfff;
rom[5438] = 12'hfff;
rom[5439] = 12'hfff;
rom[5440] = 12'hfff;
rom[5441] = 12'hfff;
rom[5442] = 12'hfff;
rom[5443] = 12'hfff;
rom[5444] = 12'hfff;
rom[5445] = 12'hfff;
rom[5446] = 12'hfff;
rom[5447] = 12'h33d;
rom[5448] = 12'h  c;
rom[5449] = 12'h  c;
rom[5450] = 12'h  c;
rom[5451] = 12'h  c;
rom[5452] = 12'h77e;
rom[5453] = 12'hfff;
rom[5454] = 12'hfff;
rom[5455] = 12'hfff;
rom[5456] = 12'hfff;
rom[5457] = 12'hfff;
rom[5458] = 12'hfff;
rom[5459] = 12'hfff;
rom[5460] = 12'hfff;
rom[5461] = 12'hfff;
rom[5462] = 12'hfff;
rom[5463] = 12'hfff;
rom[5464] = 12'hfff;
rom[5465] = 12'hfff;
rom[5466] = 12'hfff;
rom[5467] = 12'hfff;
rom[5468] = 12'hfff;
rom[5469] = 12'hfff;
rom[5470] = 12'hfff;
rom[5471] = 12'hfff;
rom[5472] = 12'hfff;
rom[5473] = 12'hfff;
rom[5474] = 12'hfff;
rom[5475] = 12'hfff;
rom[5476] = 12'hfff;
rom[5477] = 12'hfff;
rom[5478] = 12'hfff;
rom[5479] = 12'hfff;
rom[5480] = 12'hfff;
rom[5481] = 12'hfff;
rom[5482] = 12'hfff;
rom[5483] = 12'hfff;
rom[5484] = 12'hfff;
rom[5485] = 12'hfff;
rom[5486] = 12'hfff;
rom[5487] = 12'hfff;
rom[5488] = 12'hfff;
rom[5489] = 12'hfff;
rom[5490] = 12'hfff;
rom[5491] = 12'hfff;
rom[5492] = 12'hfff;
rom[5493] = 12'hfff;
rom[5494] = 12'hfff;
rom[5495] = 12'hfff;
rom[5496] = 12'hfff;
rom[5497] = 12'hfff;
rom[5498] = 12'hfff;
rom[5499] = 12'hfff;
rom[5500] = 12'hfff;
rom[5501] = 12'hfff;
rom[5502] = 12'hfff;
rom[5503] = 12'hfff;
rom[5504] = 12'hfff;
rom[5505] = 12'hfff;
rom[5506] = 12'hfff;
rom[5507] = 12'hfff;
rom[5508] = 12'hfff;
rom[5509] = 12'hfff;
rom[5510] = 12'hfff;
rom[5511] = 12'hfff;
rom[5512] = 12'hfff;
rom[5513] = 12'hfff;
rom[5514] = 12'hfff;
rom[5515] = 12'hfff;
rom[5516] = 12'hfff;
rom[5517] = 12'hfff;
rom[5518] = 12'hfff;
rom[5519] = 12'hfff;
rom[5520] = 12'hfff;
rom[5521] = 12'hfff;
rom[5522] = 12'hfff;
rom[5523] = 12'hfff;
rom[5524] = 12'hfff;
rom[5525] = 12'hfff;
rom[5526] = 12'hfff;
rom[5527] = 12'hfff;
rom[5528] = 12'hfff;
rom[5529] = 12'hfff;
rom[5530] = 12'hfff;
rom[5531] = 12'hfff;
rom[5532] = 12'hfff;
rom[5533] = 12'hfff;
rom[5534] = 12'hfff;
rom[5535] = 12'hfff;
rom[5536] = 12'hfff;
rom[5537] = 12'hfff;
rom[5538] = 12'hfff;
rom[5539] = 12'hfff;
rom[5540] = 12'hfff;
rom[5541] = 12'hfff;
rom[5542] = 12'hfff;
rom[5543] = 12'hfff;
rom[5544] = 12'hfff;
rom[5545] = 12'hfff;
rom[5546] = 12'hfff;
rom[5547] = 12'hfff;
rom[5548] = 12'hfff;
rom[5549] = 12'hfff;
rom[5550] = 12'hfff;
rom[5551] = 12'hfff;
rom[5552] = 12'hfff;
rom[5553] = 12'hfff;
rom[5554] = 12'hccf;
rom[5555] = 12'h11c;
rom[5556] = 12'h  c;
rom[5557] = 12'h  c;
rom[5558] = 12'h  c;
rom[5559] = 12'h  c;
rom[5560] = 12'h  c;
rom[5561] = 12'h77e;
rom[5562] = 12'heef;
rom[5563] = 12'hfff;
rom[5564] = 12'hfff;
rom[5565] = 12'hfff;
rom[5566] = 12'hfff;
rom[5567] = 12'hfff;
rom[5568] = 12'hfff;
rom[5569] = 12'hfff;
rom[5570] = 12'hfff;
rom[5571] = 12'hfff;
rom[5572] = 12'hfff;
rom[5573] = 12'hfff;
rom[5574] = 12'h77e;
rom[5575] = 12'h  c;
rom[5576] = 12'h  c;
rom[5577] = 12'h  c;
rom[5578] = 12'h  c;
rom[5579] = 12'h  c;
rom[5580] = 12'hbbf;
rom[5581] = 12'hfff;
rom[5582] = 12'hfff;
rom[5583] = 12'hfff;
rom[5584] = 12'hfff;
rom[5585] = 12'hfff;
rom[5586] = 12'hfff;
rom[5587] = 12'hfff;
rom[5588] = 12'hfff;
rom[5589] = 12'hfff;
rom[5590] = 12'hfff;
rom[5591] = 12'hfff;
rom[5592] = 12'hfff;
rom[5593] = 12'hfff;
rom[5594] = 12'hfff;
rom[5595] = 12'hfff;
rom[5596] = 12'hfff;
rom[5597] = 12'hfff;
rom[5598] = 12'hfff;
rom[5599] = 12'hfff;
rom[5600] = 12'hfff;
rom[5601] = 12'hfff;
rom[5602] = 12'hfff;
rom[5603] = 12'hfff;
rom[5604] = 12'hfff;
rom[5605] = 12'hfff;
rom[5606] = 12'hfff;
rom[5607] = 12'hfff;
rom[5608] = 12'hfff;
rom[5609] = 12'hfff;
rom[5610] = 12'hfff;
rom[5611] = 12'hfff;
rom[5612] = 12'hfff;
rom[5613] = 12'hfff;
rom[5614] = 12'hfff;
rom[5615] = 12'hfff;
rom[5616] = 12'hfff;
rom[5617] = 12'hfff;
rom[5618] = 12'hfff;
rom[5619] = 12'hfff;
rom[5620] = 12'hfff;
rom[5621] = 12'hfff;
rom[5622] = 12'hfff;
rom[5623] = 12'hfff;
rom[5624] = 12'hfff;
rom[5625] = 12'hfff;
rom[5626] = 12'hfff;
rom[5627] = 12'hfff;
rom[5628] = 12'hfff;
rom[5629] = 12'hfff;
rom[5630] = 12'hfff;
rom[5631] = 12'hfff;
rom[5632] = 12'hfff;
rom[5633] = 12'hfff;
rom[5634] = 12'hfff;
rom[5635] = 12'hfff;
rom[5636] = 12'hfff;
rom[5637] = 12'hfff;
rom[5638] = 12'hfff;
rom[5639] = 12'hfff;
rom[5640] = 12'hfff;
rom[5641] = 12'hfff;
rom[5642] = 12'hfff;
rom[5643] = 12'hfff;
rom[5644] = 12'hfff;
rom[5645] = 12'hfff;
rom[5646] = 12'hfff;
rom[5647] = 12'hfff;
rom[5648] = 12'hfff;
rom[5649] = 12'hfff;
rom[5650] = 12'hfff;
rom[5651] = 12'hfff;
rom[5652] = 12'hfff;
rom[5653] = 12'hfff;
rom[5654] = 12'hfff;
rom[5655] = 12'hfff;
rom[5656] = 12'hfff;
rom[5657] = 12'hfff;
rom[5658] = 12'hfff;
rom[5659] = 12'hfff;
rom[5660] = 12'hfff;
rom[5661] = 12'hfff;
rom[5662] = 12'hfff;
rom[5663] = 12'hfff;
rom[5664] = 12'hfff;
rom[5665] = 12'hfff;
rom[5666] = 12'hfff;
rom[5667] = 12'hfff;
rom[5668] = 12'hfff;
rom[5669] = 12'hfff;
rom[5670] = 12'hfff;
rom[5671] = 12'hfff;
rom[5672] = 12'hfff;
rom[5673] = 12'hfff;
rom[5674] = 12'hfff;
rom[5675] = 12'hfff;
rom[5676] = 12'hfff;
rom[5677] = 12'hfff;
rom[5678] = 12'hfff;
rom[5679] = 12'hfff;
rom[5680] = 12'hfff;
rom[5681] = 12'hfff;
rom[5682] = 12'hfff;
rom[5683] = 12'hddf;
rom[5684] = 12'h22d;
rom[5685] = 12'h  c;
rom[5686] = 12'h  c;
rom[5687] = 12'h  c;
rom[5688] = 12'h  c;
rom[5689] = 12'h  c;
rom[5690] = 12'h22d;
rom[5691] = 12'heef;
rom[5692] = 12'hfff;
rom[5693] = 12'hfff;
rom[5694] = 12'hfff;
rom[5695] = 12'hfff;
rom[5696] = 12'hfff;
rom[5697] = 12'hfff;
rom[5698] = 12'hfff;
rom[5699] = 12'hfff;
rom[5700] = 12'hfff;
rom[5701] = 12'hfff;
rom[5702] = 12'h11d;
rom[5703] = 12'h  c;
rom[5704] = 12'h  c;
rom[5705] = 12'h  c;
rom[5706] = 12'h  c;
rom[5707] = 12'h44d;
rom[5708] = 12'hfff;
rom[5709] = 12'hfff;
rom[5710] = 12'hfff;
rom[5711] = 12'hfff;
rom[5712] = 12'hfff;
rom[5713] = 12'hfff;
rom[5714] = 12'hfff;
rom[5715] = 12'hfff;
rom[5716] = 12'hfff;
rom[5717] = 12'hfff;
rom[5718] = 12'hfff;
rom[5719] = 12'hfff;
rom[5720] = 12'hfff;
rom[5721] = 12'hfff;
rom[5722] = 12'hfff;
rom[5723] = 12'hfff;
rom[5724] = 12'hfff;
rom[5725] = 12'hfff;
rom[5726] = 12'hfff;
rom[5727] = 12'hfff;
rom[5728] = 12'hfff;
rom[5729] = 12'hfff;
rom[5730] = 12'hfff;
rom[5731] = 12'hfff;
rom[5732] = 12'hfff;
rom[5733] = 12'hfff;
rom[5734] = 12'hfff;
rom[5735] = 12'hfff;
rom[5736] = 12'hfff;
rom[5737] = 12'hfff;
rom[5738] = 12'hfff;
rom[5739] = 12'hfff;
rom[5740] = 12'hfff;
rom[5741] = 12'hfff;
rom[5742] = 12'hfff;
rom[5743] = 12'hfff;
rom[5744] = 12'hfff;
rom[5745] = 12'hfff;
rom[5746] = 12'hfff;
rom[5747] = 12'hfff;
rom[5748] = 12'hfff;
rom[5749] = 12'hfff;
rom[5750] = 12'hfff;
rom[5751] = 12'hfff;
rom[5752] = 12'hfff;
rom[5753] = 12'hfff;
rom[5754] = 12'hfff;
rom[5755] = 12'hfff;
rom[5756] = 12'hfff;
rom[5757] = 12'hfff;
rom[5758] = 12'hfff;
rom[5759] = 12'hfff;
rom[5760] = 12'hfff;
rom[5761] = 12'hfff;
rom[5762] = 12'hfff;
rom[5763] = 12'hfff;
rom[5764] = 12'hfff;
rom[5765] = 12'hfff;
rom[5766] = 12'hfff;
rom[5767] = 12'hfff;
rom[5768] = 12'hfff;
rom[5769] = 12'hfff;
rom[5770] = 12'hfff;
rom[5771] = 12'hfff;
rom[5772] = 12'hfff;
rom[5773] = 12'hfff;
rom[5774] = 12'hfff;
rom[5775] = 12'hfff;
rom[5776] = 12'hfff;
rom[5777] = 12'hfff;
rom[5778] = 12'hfff;
rom[5779] = 12'hfff;
rom[5780] = 12'hfff;
rom[5781] = 12'hfff;
rom[5782] = 12'hfff;
rom[5783] = 12'hfff;
rom[5784] = 12'hfff;
rom[5785] = 12'hfff;
rom[5786] = 12'hfff;
rom[5787] = 12'hfff;
rom[5788] = 12'hfff;
rom[5789] = 12'hfff;
rom[5790] = 12'hfff;
rom[5791] = 12'hfff;
rom[5792] = 12'hfff;
rom[5793] = 12'hfff;
rom[5794] = 12'hfff;
rom[5795] = 12'hfff;
rom[5796] = 12'hfff;
rom[5797] = 12'hfff;
rom[5798] = 12'hfff;
rom[5799] = 12'hfff;
rom[5800] = 12'hfff;
rom[5801] = 12'hfff;
rom[5802] = 12'hfff;
rom[5803] = 12'hfff;
rom[5804] = 12'hfff;
rom[5805] = 12'hfff;
rom[5806] = 12'hfff;
rom[5807] = 12'hfff;
rom[5808] = 12'hfff;
rom[5809] = 12'hfff;
rom[5810] = 12'hfff;
rom[5811] = 12'hfff;
rom[5812] = 12'heef;
rom[5813] = 12'h11d;
rom[5814] = 12'h  c;
rom[5815] = 12'h  c;
rom[5816] = 12'h  c;
rom[5817] = 12'h  c;
rom[5818] = 12'h  c;
rom[5819] = 12'h66e;
rom[5820] = 12'hfff;
rom[5821] = 12'hfff;
rom[5822] = 12'hfff;
rom[5823] = 12'hfff;
rom[5824] = 12'hfff;
rom[5825] = 12'hfff;
rom[5826] = 12'hfff;
rom[5827] = 12'hfff;
rom[5828] = 12'hfff;
rom[5829] = 12'heef;
rom[5830] = 12'h  c;
rom[5831] = 12'h  c;
rom[5832] = 12'h  c;
rom[5833] = 12'h  c;
rom[5834] = 12'h  c;
rom[5835] = 12'heef;
rom[5836] = 12'hfff;
rom[5837] = 12'hfff;
rom[5838] = 12'hfff;
rom[5839] = 12'hfff;
rom[5840] = 12'hfff;
rom[5841] = 12'hfff;
rom[5842] = 12'hfff;
rom[5843] = 12'hfff;
rom[5844] = 12'hfff;
rom[5845] = 12'hfff;
rom[5846] = 12'hfff;
rom[5847] = 12'hfff;
rom[5848] = 12'hfff;
rom[5849] = 12'hfff;
rom[5850] = 12'hfff;
rom[5851] = 12'hfff;
rom[5852] = 12'hfff;
rom[5853] = 12'hfff;
rom[5854] = 12'hfff;
rom[5855] = 12'hfff;
rom[5856] = 12'hfff;
rom[5857] = 12'hfff;
rom[5858] = 12'hfff;
rom[5859] = 12'hfff;
rom[5860] = 12'hfff;
rom[5861] = 12'hfff;
rom[5862] = 12'hfff;
rom[5863] = 12'hfff;
rom[5864] = 12'hfff;
rom[5865] = 12'hfff;
rom[5866] = 12'hfff;
rom[5867] = 12'hfff;
rom[5868] = 12'hfff;
rom[5869] = 12'hfff;
rom[5870] = 12'hfff;
rom[5871] = 12'hfff;
rom[5872] = 12'hfff;
rom[5873] = 12'hfff;
rom[5874] = 12'hfff;
rom[5875] = 12'hfff;
rom[5876] = 12'hfff;
rom[5877] = 12'hfff;
rom[5878] = 12'hfff;
rom[5879] = 12'hfff;
rom[5880] = 12'hfff;
rom[5881] = 12'hfff;
rom[5882] = 12'hfff;
rom[5883] = 12'hfff;
rom[5884] = 12'hfff;
rom[5885] = 12'hfff;
rom[5886] = 12'hfff;
rom[5887] = 12'hfff;
rom[5888] = 12'hfff;
rom[5889] = 12'hfff;
rom[5890] = 12'hfff;
rom[5891] = 12'hfff;
rom[5892] = 12'hfff;
rom[5893] = 12'hfff;
rom[5894] = 12'hfff;
rom[5895] = 12'hfff;
rom[5896] = 12'hfff;
rom[5897] = 12'hfff;
rom[5898] = 12'hfff;
rom[5899] = 12'hfff;
rom[5900] = 12'hfff;
rom[5901] = 12'hfff;
rom[5902] = 12'hfff;
rom[5903] = 12'hfff;
rom[5904] = 12'hfff;
rom[5905] = 12'hfff;
rom[5906] = 12'hfff;
rom[5907] = 12'hfff;
rom[5908] = 12'hfff;
rom[5909] = 12'hfff;
rom[5910] = 12'hfff;
rom[5911] = 12'hfff;
rom[5912] = 12'hfff;
rom[5913] = 12'hfff;
rom[5914] = 12'hfff;
rom[5915] = 12'hfff;
rom[5916] = 12'hfff;
rom[5917] = 12'hfff;
rom[5918] = 12'hfff;
rom[5919] = 12'hfff;
rom[5920] = 12'hfff;
rom[5921] = 12'hfff;
rom[5922] = 12'hfff;
rom[5923] = 12'hfff;
rom[5924] = 12'hfff;
rom[5925] = 12'hfff;
rom[5926] = 12'hfff;
rom[5927] = 12'hfff;
rom[5928] = 12'hfff;
rom[5929] = 12'hfff;
rom[5930] = 12'hfff;
rom[5931] = 12'hfff;
rom[5932] = 12'hfff;
rom[5933] = 12'hfff;
rom[5934] = 12'hfff;
rom[5935] = 12'hfff;
rom[5936] = 12'hfff;
rom[5937] = 12'hfff;
rom[5938] = 12'hfff;
rom[5939] = 12'hfff;
rom[5940] = 12'hfff;
rom[5941] = 12'h77e;
rom[5942] = 12'h  c;
rom[5943] = 12'h  c;
rom[5944] = 12'h  c;
rom[5945] = 12'h  c;
rom[5946] = 12'h  c;
rom[5947] = 12'h  c;
rom[5948] = 12'hccf;
rom[5949] = 12'hfff;
rom[5950] = 12'hfff;
rom[5951] = 12'hfff;
rom[5952] = 12'hfff;
rom[5953] = 12'hfff;
rom[5954] = 12'hfff;
rom[5955] = 12'hfff;
rom[5956] = 12'hfff;
rom[5957] = 12'hccf;
rom[5958] = 12'h  c;
rom[5959] = 12'h  c;
rom[5960] = 12'h  c;
rom[5961] = 12'h  c;
rom[5962] = 12'h33d;
rom[5963] = 12'hfff;
rom[5964] = 12'hfff;
rom[5965] = 12'hfff;
rom[5966] = 12'hfff;
rom[5967] = 12'hfff;
rom[5968] = 12'hfff;
rom[5969] = 12'hfff;
rom[5970] = 12'hfff;
rom[5971] = 12'hfff;
rom[5972] = 12'hfff;
rom[5973] = 12'hfff;
rom[5974] = 12'hfff;
rom[5975] = 12'hfff;
rom[5976] = 12'hfff;
rom[5977] = 12'hfff;
rom[5978] = 12'hfff;
rom[5979] = 12'hfff;
rom[5980] = 12'hfff;
rom[5981] = 12'hfff;
rom[5982] = 12'hfff;
rom[5983] = 12'hfff;
rom[5984] = 12'hfff;
rom[5985] = 12'hfff;
rom[5986] = 12'hfff;
rom[5987] = 12'hfff;
rom[5988] = 12'hfff;
rom[5989] = 12'hfff;
rom[5990] = 12'hfff;
rom[5991] = 12'hfff;
rom[5992] = 12'hfff;
rom[5993] = 12'hfff;
rom[5994] = 12'hfff;
rom[5995] = 12'hfff;
rom[5996] = 12'hfff;
rom[5997] = 12'hfff;
rom[5998] = 12'hfff;
rom[5999] = 12'hfff;
rom[6000] = 12'hfff;
rom[6001] = 12'hfff;
rom[6002] = 12'hfff;
rom[6003] = 12'hfff;
rom[6004] = 12'hfff;
rom[6005] = 12'hfff;
rom[6006] = 12'hfff;
rom[6007] = 12'hfff;
rom[6008] = 12'hfff;
rom[6009] = 12'hfff;
rom[6010] = 12'hfff;
rom[6011] = 12'hfff;
rom[6012] = 12'hfff;
rom[6013] = 12'hfff;
rom[6014] = 12'hfff;
rom[6015] = 12'hfff;
rom[6016] = 12'hfff;
rom[6017] = 12'hfff;
rom[6018] = 12'hfff;
rom[6019] = 12'hfff;
rom[6020] = 12'hfff;
rom[6021] = 12'hfff;
rom[6022] = 12'hfff;
rom[6023] = 12'hfff;
rom[6024] = 12'hfff;
rom[6025] = 12'hfff;
rom[6026] = 12'hfff;
rom[6027] = 12'hfff;
rom[6028] = 12'hfff;
rom[6029] = 12'hfff;
rom[6030] = 12'hfff;
rom[6031] = 12'hfff;
rom[6032] = 12'hfff;
rom[6033] = 12'hfff;
rom[6034] = 12'hfff;
rom[6035] = 12'hfff;
rom[6036] = 12'hfff;
rom[6037] = 12'hfff;
rom[6038] = 12'hfff;
rom[6039] = 12'hfff;
rom[6040] = 12'hfff;
rom[6041] = 12'hfff;
rom[6042] = 12'hfff;
rom[6043] = 12'hfff;
rom[6044] = 12'hfff;
rom[6045] = 12'hfff;
rom[6046] = 12'hfff;
rom[6047] = 12'hfff;
rom[6048] = 12'hfff;
rom[6049] = 12'hfff;
rom[6050] = 12'hfff;
rom[6051] = 12'hfff;
rom[6052] = 12'hfff;
rom[6053] = 12'hfff;
rom[6054] = 12'hfff;
rom[6055] = 12'hfff;
rom[6056] = 12'hfff;
rom[6057] = 12'hfff;
rom[6058] = 12'hfff;
rom[6059] = 12'hfff;
rom[6060] = 12'hfff;
rom[6061] = 12'hfff;
rom[6062] = 12'hfff;
rom[6063] = 12'hfff;
rom[6064] = 12'hfff;
rom[6065] = 12'hfff;
rom[6066] = 12'hfff;
rom[6067] = 12'hfff;
rom[6068] = 12'hfff;
rom[6069] = 12'hfff;
rom[6070] = 12'h99e;
rom[6071] = 12'h11d;
rom[6072] = 12'h  c;
rom[6073] = 12'h  c;
rom[6074] = 12'h  c;
rom[6075] = 12'h  c;
rom[6076] = 12'h44d;
rom[6077] = 12'hfff;
rom[6078] = 12'hfff;
rom[6079] = 12'hfff;
rom[6080] = 12'hfff;
rom[6081] = 12'hfff;
rom[6082] = 12'hfff;
rom[6083] = 12'hfff;
rom[6084] = 12'hfff;
rom[6085] = 12'h99e;
rom[6086] = 12'h  c;
rom[6087] = 12'h  c;
rom[6088] = 12'h  c;
rom[6089] = 12'h  c;
rom[6090] = 12'h55d;
rom[6091] = 12'hfff;
rom[6092] = 12'hfff;
rom[6093] = 12'hfff;
rom[6094] = 12'hfff;
rom[6095] = 12'hfff;
rom[6096] = 12'hfff;
rom[6097] = 12'hfff;
rom[6098] = 12'hfff;
rom[6099] = 12'hfff;
rom[6100] = 12'hfff;
rom[6101] = 12'hfff;
rom[6102] = 12'hfff;
rom[6103] = 12'hfff;
rom[6104] = 12'hfff;
rom[6105] = 12'hfff;
rom[6106] = 12'hfff;
rom[6107] = 12'hfff;
rom[6108] = 12'hfff;
rom[6109] = 12'hfff;
rom[6110] = 12'hfff;
rom[6111] = 12'hfff;
rom[6112] = 12'hfff;
rom[6113] = 12'hfff;
rom[6114] = 12'hfff;
rom[6115] = 12'hfff;
rom[6116] = 12'hfff;
rom[6117] = 12'hfff;
rom[6118] = 12'hfff;
rom[6119] = 12'hfff;
rom[6120] = 12'hfff;
rom[6121] = 12'hfff;
rom[6122] = 12'hfff;
rom[6123] = 12'hfff;
rom[6124] = 12'hfff;
rom[6125] = 12'hfff;
rom[6126] = 12'hfff;
rom[6127] = 12'hfff;
rom[6128] = 12'hfff;
rom[6129] = 12'hfff;
rom[6130] = 12'hfff;
rom[6131] = 12'hfff;
rom[6132] = 12'hfff;
rom[6133] = 12'hfff;
rom[6134] = 12'hfff;
rom[6135] = 12'hfff;
rom[6136] = 12'hfff;
rom[6137] = 12'hfff;
rom[6138] = 12'hfff;
rom[6139] = 12'hfff;
rom[6140] = 12'hfff;
rom[6141] = 12'hfff;
rom[6142] = 12'hfff;
rom[6143] = 12'hfff;
rom[6144] = 12'hfff;
rom[6145] = 12'hfff;
rom[6146] = 12'hfff;
rom[6147] = 12'hfff;
rom[6148] = 12'hfff;
rom[6149] = 12'hfff;
rom[6150] = 12'hfff;
rom[6151] = 12'hfff;
rom[6152] = 12'hfff;
rom[6153] = 12'hfff;
rom[6154] = 12'hfff;
rom[6155] = 12'hfff;
rom[6156] = 12'hfff;
rom[6157] = 12'hfff;
rom[6158] = 12'hfff;
rom[6159] = 12'hfff;
rom[6160] = 12'hfff;
rom[6161] = 12'hfff;
rom[6162] = 12'hfff;
rom[6163] = 12'hfff;
rom[6164] = 12'hfff;
rom[6165] = 12'hfff;
rom[6166] = 12'hfff;
rom[6167] = 12'hfff;
rom[6168] = 12'hfff;
rom[6169] = 12'hfff;
rom[6170] = 12'hfff;
rom[6171] = 12'hfff;
rom[6172] = 12'hfff;
rom[6173] = 12'hfff;
rom[6174] = 12'hfff;
rom[6175] = 12'hfff;
rom[6176] = 12'hfff;
rom[6177] = 12'hfff;
rom[6178] = 12'hfff;
rom[6179] = 12'hfff;
rom[6180] = 12'hfff;
rom[6181] = 12'hfff;
rom[6182] = 12'hfff;
rom[6183] = 12'hfff;
rom[6184] = 12'hfff;
rom[6185] = 12'hfff;
rom[6186] = 12'hfff;
rom[6187] = 12'hfff;
rom[6188] = 12'hfff;
rom[6189] = 12'hfff;
rom[6190] = 12'hfff;
rom[6191] = 12'hfff;
rom[6192] = 12'hfff;
rom[6193] = 12'hfff;
rom[6194] = 12'hfff;
rom[6195] = 12'hfff;
rom[6196] = 12'hfff;
rom[6197] = 12'hfff;
rom[6198] = 12'hfff;
rom[6199] = 12'h99e;
rom[6200] = 12'h  c;
rom[6201] = 12'h  c;
rom[6202] = 12'h  c;
rom[6203] = 12'h  c;
rom[6204] = 12'h  c;
rom[6205] = 12'h33d;
rom[6206] = 12'heef;
rom[6207] = 12'hfff;
rom[6208] = 12'hfff;
rom[6209] = 12'hfff;
rom[6210] = 12'hfff;
rom[6211] = 12'hfff;
rom[6212] = 12'hfff;
rom[6213] = 12'h88e;
rom[6214] = 12'h  c;
rom[6215] = 12'h  c;
rom[6216] = 12'h  c;
rom[6217] = 12'h  c;
rom[6218] = 12'h77e;
rom[6219] = 12'hfff;
rom[6220] = 12'hfff;
rom[6221] = 12'hfff;
rom[6222] = 12'hfff;
rom[6223] = 12'hfff;
rom[6224] = 12'hfff;
rom[6225] = 12'hfff;
rom[6226] = 12'hfff;
rom[6227] = 12'hfff;
rom[6228] = 12'hfff;
rom[6229] = 12'hfff;
rom[6230] = 12'hfff;
rom[6231] = 12'hfff;
rom[6232] = 12'hfff;
rom[6233] = 12'hfff;
rom[6234] = 12'hfff;
rom[6235] = 12'hfff;
rom[6236] = 12'hfff;
rom[6237] = 12'hfff;
rom[6238] = 12'hfff;
rom[6239] = 12'hfff;
rom[6240] = 12'hfff;
rom[6241] = 12'hfff;
rom[6242] = 12'hfff;
rom[6243] = 12'hfff;
rom[6244] = 12'hfff;
rom[6245] = 12'hfff;
rom[6246] = 12'hfff;
rom[6247] = 12'hfff;
rom[6248] = 12'hfff;
rom[6249] = 12'hfff;
rom[6250] = 12'hfff;
rom[6251] = 12'hfff;
rom[6252] = 12'hfff;
rom[6253] = 12'hfff;
rom[6254] = 12'hfff;
rom[6255] = 12'hfff;
rom[6256] = 12'hfff;
rom[6257] = 12'hfff;
rom[6258] = 12'hfff;
rom[6259] = 12'hfff;
rom[6260] = 12'hfff;
rom[6261] = 12'hfff;
rom[6262] = 12'hfff;
rom[6263] = 12'hfff;
rom[6264] = 12'hfff;
rom[6265] = 12'hfff;
rom[6266] = 12'hfff;
rom[6267] = 12'hfff;
rom[6268] = 12'hfff;
rom[6269] = 12'hfff;
rom[6270] = 12'hfff;
rom[6271] = 12'hfff;
rom[6272] = 12'hfff;
rom[6273] = 12'hfff;
rom[6274] = 12'hfff;
rom[6275] = 12'hfff;
rom[6276] = 12'hfff;
rom[6277] = 12'hfff;
rom[6278] = 12'hfff;
rom[6279] = 12'hfff;
rom[6280] = 12'hfff;
rom[6281] = 12'hfff;
rom[6282] = 12'hfff;
rom[6283] = 12'hfff;
rom[6284] = 12'hfff;
rom[6285] = 12'hfff;
rom[6286] = 12'hfff;
rom[6287] = 12'hfff;
rom[6288] = 12'hfff;
rom[6289] = 12'hfff;
rom[6290] = 12'hfff;
rom[6291] = 12'hfff;
rom[6292] = 12'hfff;
rom[6293] = 12'hfff;
rom[6294] = 12'hfff;
rom[6295] = 12'hfff;
rom[6296] = 12'hfff;
rom[6297] = 12'hfff;
rom[6298] = 12'hfff;
rom[6299] = 12'hfff;
rom[6300] = 12'hfff;
rom[6301] = 12'hfff;
rom[6302] = 12'hfff;
rom[6303] = 12'hfff;
rom[6304] = 12'hfff;
rom[6305] = 12'hfff;
rom[6306] = 12'hfff;
rom[6307] = 12'hfff;
rom[6308] = 12'hfff;
rom[6309] = 12'hfff;
rom[6310] = 12'hfff;
rom[6311] = 12'hfff;
rom[6312] = 12'hfff;
rom[6313] = 12'hfff;
rom[6314] = 12'hfff;
rom[6315] = 12'hfff;
rom[6316] = 12'hfff;
rom[6317] = 12'hfff;
rom[6318] = 12'hfff;
rom[6319] = 12'hfff;
rom[6320] = 12'hfff;
rom[6321] = 12'hfff;
rom[6322] = 12'hfff;
rom[6323] = 12'hfff;
rom[6324] = 12'hfff;
rom[6325] = 12'hfff;
rom[6326] = 12'hfff;
rom[6327] = 12'heef;
rom[6328] = 12'h11d;
rom[6329] = 12'h  c;
rom[6330] = 12'h  c;
rom[6331] = 12'h  c;
rom[6332] = 12'h  c;
rom[6333] = 12'h  c;
rom[6334] = 12'h22d;
rom[6335] = 12'hddf;
rom[6336] = 12'hfff;
rom[6337] = 12'hfff;
rom[6338] = 12'hfff;
rom[6339] = 12'hfff;
rom[6340] = 12'hfff;
rom[6341] = 12'h77e;
rom[6342] = 12'h  c;
rom[6343] = 12'h  c;
rom[6344] = 12'h  c;
rom[6345] = 12'h  c;
rom[6346] = 12'h88e;
rom[6347] = 12'hfff;
rom[6348] = 12'hfff;
rom[6349] = 12'hfff;
rom[6350] = 12'hfff;
rom[6351] = 12'hfff;
rom[6352] = 12'hfff;
rom[6353] = 12'hfff;
rom[6354] = 12'hfff;
rom[6355] = 12'hfff;
rom[6356] = 12'hfff;
rom[6357] = 12'hfff;
rom[6358] = 12'hfff;
rom[6359] = 12'hfff;
rom[6360] = 12'hfff;
rom[6361] = 12'hfff;
rom[6362] = 12'hfff;
rom[6363] = 12'hfff;
rom[6364] = 12'hfff;
rom[6365] = 12'hfff;
rom[6366] = 12'hfff;
rom[6367] = 12'hfff;
rom[6368] = 12'hfff;
rom[6369] = 12'hfff;
rom[6370] = 12'hfff;
rom[6371] = 12'hfff;
rom[6372] = 12'hfff;
rom[6373] = 12'hfff;
rom[6374] = 12'hfff;
rom[6375] = 12'hfff;
rom[6376] = 12'hfff;
rom[6377] = 12'hfff;
rom[6378] = 12'hfff;
rom[6379] = 12'hfff;
rom[6380] = 12'hfff;
rom[6381] = 12'hfff;
rom[6382] = 12'hfff;
rom[6383] = 12'hfff;
rom[6384] = 12'hfff;
rom[6385] = 12'hfff;
rom[6386] = 12'hfff;
rom[6387] = 12'hfff;
rom[6388] = 12'hfff;
rom[6389] = 12'hfff;
rom[6390] = 12'hfff;
rom[6391] = 12'hfff;
rom[6392] = 12'hfff;
rom[6393] = 12'hfff;
rom[6394] = 12'hfff;
rom[6395] = 12'hfff;
rom[6396] = 12'hfff;
rom[6397] = 12'hfff;
rom[6398] = 12'hfff;
rom[6399] = 12'hfff;
rom[6400] = 12'hfff;
rom[6401] = 12'hfff;
rom[6402] = 12'hfff;
rom[6403] = 12'hfff;
rom[6404] = 12'hfff;
rom[6405] = 12'hfff;
rom[6406] = 12'hfff;
rom[6407] = 12'hfff;
rom[6408] = 12'hfff;
rom[6409] = 12'hfff;
rom[6410] = 12'hfff;
rom[6411] = 12'hfff;
rom[6412] = 12'hfff;
rom[6413] = 12'hfff;
rom[6414] = 12'hfff;
rom[6415] = 12'hfff;
rom[6416] = 12'hfff;
rom[6417] = 12'hfff;
rom[6418] = 12'hfff;
rom[6419] = 12'hfff;
rom[6420] = 12'hfff;
rom[6421] = 12'hfff;
rom[6422] = 12'hfff;
rom[6423] = 12'hfff;
rom[6424] = 12'hfff;
rom[6425] = 12'hfff;
rom[6426] = 12'hfff;
rom[6427] = 12'hfff;
rom[6428] = 12'hfff;
rom[6429] = 12'hfff;
rom[6430] = 12'hfff;
rom[6431] = 12'hfff;
rom[6432] = 12'hfff;
rom[6433] = 12'hfff;
rom[6434] = 12'hfff;
rom[6435] = 12'hfff;
rom[6436] = 12'hfff;
rom[6437] = 12'hfff;
rom[6438] = 12'hfff;
rom[6439] = 12'hfff;
rom[6440] = 12'hfff;
rom[6441] = 12'hfff;
rom[6442] = 12'hfff;
rom[6443] = 12'hfff;
rom[6444] = 12'hfff;
rom[6445] = 12'hfff;
rom[6446] = 12'hfff;
rom[6447] = 12'hfff;
rom[6448] = 12'hfff;
rom[6449] = 12'hfff;
rom[6450] = 12'hfff;
rom[6451] = 12'hfff;
rom[6452] = 12'hfff;
rom[6453] = 12'hfff;
rom[6454] = 12'hfff;
rom[6455] = 12'hfff;
rom[6456] = 12'hbbf;
rom[6457] = 12'h  c;
rom[6458] = 12'h  c;
rom[6459] = 12'h  c;
rom[6460] = 12'h  c;
rom[6461] = 12'h  c;
rom[6462] = 12'h  c;
rom[6463] = 12'h11d;
rom[6464] = 12'hccf;
rom[6465] = 12'hfff;
rom[6466] = 12'hfff;
rom[6467] = 12'hfff;
rom[6468] = 12'hfff;
rom[6469] = 12'h66e;
rom[6470] = 12'h  c;
rom[6471] = 12'h  c;
rom[6472] = 12'h  c;
rom[6473] = 12'h  c;
rom[6474] = 12'h99e;
rom[6475] = 12'hfff;
rom[6476] = 12'hfff;
rom[6477] = 12'hfff;
rom[6478] = 12'hfff;
rom[6479] = 12'hfff;
rom[6480] = 12'hfff;
rom[6481] = 12'hfff;
rom[6482] = 12'hfff;
rom[6483] = 12'hfff;
rom[6484] = 12'hfff;
rom[6485] = 12'hfff;
rom[6486] = 12'hfff;
rom[6487] = 12'hfff;
rom[6488] = 12'hfff;
rom[6489] = 12'hfff;
rom[6490] = 12'hfff;
rom[6491] = 12'hfff;
rom[6492] = 12'hfff;
rom[6493] = 12'hfff;
rom[6494] = 12'hfff;
rom[6495] = 12'hfff;
rom[6496] = 12'hfff;
rom[6497] = 12'hfff;
rom[6498] = 12'hfff;
rom[6499] = 12'hfff;
rom[6500] = 12'hfff;
rom[6501] = 12'hfff;
rom[6502] = 12'hfff;
rom[6503] = 12'hfff;
rom[6504] = 12'hfff;
rom[6505] = 12'hfff;
rom[6506] = 12'hfff;
rom[6507] = 12'hfff;
rom[6508] = 12'hfff;
rom[6509] = 12'hfff;
rom[6510] = 12'hfff;
rom[6511] = 12'hfff;
rom[6512] = 12'hfff;
rom[6513] = 12'hfff;
rom[6514] = 12'hfff;
rom[6515] = 12'hfff;
rom[6516] = 12'hfff;
rom[6517] = 12'hfff;
rom[6518] = 12'hfff;
rom[6519] = 12'hfff;
rom[6520] = 12'hfff;
rom[6521] = 12'hfff;
rom[6522] = 12'hfff;
rom[6523] = 12'hfff;
rom[6524] = 12'hfff;
rom[6525] = 12'hfff;
rom[6526] = 12'hfff;
rom[6527] = 12'hfff;
rom[6528] = 12'hfff;
rom[6529] = 12'hfff;
rom[6530] = 12'hfff;
rom[6531] = 12'hfff;
rom[6532] = 12'hfff;
rom[6533] = 12'hfff;
rom[6534] = 12'hfff;
rom[6535] = 12'hfff;
rom[6536] = 12'hfff;
rom[6537] = 12'hfff;
rom[6538] = 12'hfff;
rom[6539] = 12'hfff;
rom[6540] = 12'hfff;
rom[6541] = 12'hfff;
rom[6542] = 12'hfff;
rom[6543] = 12'hfff;
rom[6544] = 12'hfff;
rom[6545] = 12'hfff;
rom[6546] = 12'hfff;
rom[6547] = 12'hfff;
rom[6548] = 12'hfff;
rom[6549] = 12'hfff;
rom[6550] = 12'hfff;
rom[6551] = 12'hfff;
rom[6552] = 12'hfff;
rom[6553] = 12'hfff;
rom[6554] = 12'hfff;
rom[6555] = 12'hfff;
rom[6556] = 12'hfff;
rom[6557] = 12'hfff;
rom[6558] = 12'hfff;
rom[6559] = 12'hfff;
rom[6560] = 12'hfff;
rom[6561] = 12'hfff;
rom[6562] = 12'hfff;
rom[6563] = 12'hfff;
rom[6564] = 12'hfff;
rom[6565] = 12'hfff;
rom[6566] = 12'hfff;
rom[6567] = 12'hfff;
rom[6568] = 12'hfff;
rom[6569] = 12'hfff;
rom[6570] = 12'hfff;
rom[6571] = 12'hfff;
rom[6572] = 12'hfff;
rom[6573] = 12'hfff;
rom[6574] = 12'hfff;
rom[6575] = 12'hfff;
rom[6576] = 12'hfff;
rom[6577] = 12'hfff;
rom[6578] = 12'hfff;
rom[6579] = 12'hfff;
rom[6580] = 12'hfff;
rom[6581] = 12'hfff;
rom[6582] = 12'hfff;
rom[6583] = 12'hfff;
rom[6584] = 12'hfff;
rom[6585] = 12'hbbf;
rom[6586] = 12'h  c;
rom[6587] = 12'h  c;
rom[6588] = 12'h  c;
rom[6589] = 12'h  c;
rom[6590] = 12'h  c;
rom[6591] = 12'h  c;
rom[6592] = 12'h  c;
rom[6593] = 12'hbbe;
rom[6594] = 12'hfff;
rom[6595] = 12'hfff;
rom[6596] = 12'hfff;
rom[6597] = 12'h55d;
rom[6598] = 12'h  c;
rom[6599] = 12'h  c;
rom[6600] = 12'h  c;
rom[6601] = 12'h  c;
rom[6602] = 12'haae;
rom[6603] = 12'hfff;
rom[6604] = 12'hfff;
rom[6605] = 12'hfff;
rom[6606] = 12'hfff;
rom[6607] = 12'hfff;
rom[6608] = 12'hfff;
rom[6609] = 12'hfff;
rom[6610] = 12'hfff;
rom[6611] = 12'hfff;
rom[6612] = 12'hfff;
rom[6613] = 12'hfff;
rom[6614] = 12'hfff;
rom[6615] = 12'hfff;
rom[6616] = 12'hfff;
rom[6617] = 12'hfff;
rom[6618] = 12'hfff;
rom[6619] = 12'hfff;
rom[6620] = 12'hfff;
rom[6621] = 12'hfff;
rom[6622] = 12'hfff;
rom[6623] = 12'hfff;
rom[6624] = 12'hfff;
rom[6625] = 12'hfff;
rom[6626] = 12'hfff;
rom[6627] = 12'hfff;
rom[6628] = 12'hfff;
rom[6629] = 12'hfff;
rom[6630] = 12'hfff;
rom[6631] = 12'hfff;
rom[6632] = 12'hfff;
rom[6633] = 12'hfff;
rom[6634] = 12'hfff;
rom[6635] = 12'hfff;
rom[6636] = 12'hfff;
rom[6637] = 12'hfff;
rom[6638] = 12'hfff;
rom[6639] = 12'hfff;
rom[6640] = 12'hfff;
rom[6641] = 12'hfff;
rom[6642] = 12'hfff;
rom[6643] = 12'hfff;
rom[6644] = 12'hfff;
rom[6645] = 12'hfff;
rom[6646] = 12'hfff;
rom[6647] = 12'hfff;
rom[6648] = 12'hfff;
rom[6649] = 12'hfff;
rom[6650] = 12'hfff;
rom[6651] = 12'hfff;
rom[6652] = 12'hfff;
rom[6653] = 12'hfff;
rom[6654] = 12'hfff;
rom[6655] = 12'hfff;
rom[6656] = 12'hfff;
rom[6657] = 12'hfff;
rom[6658] = 12'hfff;
rom[6659] = 12'hfff;
rom[6660] = 12'hfff;
rom[6661] = 12'hfff;
rom[6662] = 12'hfff;
rom[6663] = 12'hfff;
rom[6664] = 12'hfff;
rom[6665] = 12'hfff;
rom[6666] = 12'hfff;
rom[6667] = 12'hfff;
rom[6668] = 12'hfff;
rom[6669] = 12'hfff;
rom[6670] = 12'hfff;
rom[6671] = 12'hfff;
rom[6672] = 12'hfff;
rom[6673] = 12'hfff;
rom[6674] = 12'hfff;
rom[6675] = 12'hfff;
rom[6676] = 12'hfff;
rom[6677] = 12'hfff;
rom[6678] = 12'hfff;
rom[6679] = 12'hfff;
rom[6680] = 12'hfff;
rom[6681] = 12'hfff;
rom[6682] = 12'hfff;
rom[6683] = 12'hfff;
rom[6684] = 12'hfff;
rom[6685] = 12'hfff;
rom[6686] = 12'hfff;
rom[6687] = 12'hfff;
rom[6688] = 12'hfff;
rom[6689] = 12'hfff;
rom[6690] = 12'hfff;
rom[6691] = 12'hfff;
rom[6692] = 12'hfff;
rom[6693] = 12'hfff;
rom[6694] = 12'hfff;
rom[6695] = 12'hfff;
rom[6696] = 12'hfff;
rom[6697] = 12'hfff;
rom[6698] = 12'hfff;
rom[6699] = 12'hfff;
rom[6700] = 12'hfff;
rom[6701] = 12'hfff;
rom[6702] = 12'hfff;
rom[6703] = 12'hfff;
rom[6704] = 12'hfff;
rom[6705] = 12'hfff;
rom[6706] = 12'hfff;
rom[6707] = 12'hfff;
rom[6708] = 12'hfff;
rom[6709] = 12'hfff;
rom[6710] = 12'hfff;
rom[6711] = 12'hfff;
rom[6712] = 12'hfff;
rom[6713] = 12'hfff;
rom[6714] = 12'hccf;
rom[6715] = 12'h11d;
rom[6716] = 12'h  c;
rom[6717] = 12'h  c;
rom[6718] = 12'h  c;
rom[6719] = 12'h  c;
rom[6720] = 12'h  c;
rom[6721] = 12'h  c;
rom[6722] = 12'hbbf;
rom[6723] = 12'hfff;
rom[6724] = 12'hfff;
rom[6725] = 12'h44d;
rom[6726] = 12'h  c;
rom[6727] = 12'h  c;
rom[6728] = 12'h  c;
rom[6729] = 12'h  c;
rom[6730] = 12'hbbf;
rom[6731] = 12'hfff;
rom[6732] = 12'hfff;
rom[6733] = 12'hfff;
rom[6734] = 12'hfff;
rom[6735] = 12'hfff;
rom[6736] = 12'hfff;
rom[6737] = 12'hfff;
rom[6738] = 12'hfff;
rom[6739] = 12'hfff;
rom[6740] = 12'hfff;
rom[6741] = 12'hfff;
rom[6742] = 12'hfff;
rom[6743] = 12'hfff;
rom[6744] = 12'hfff;
rom[6745] = 12'hfff;
rom[6746] = 12'hfff;
rom[6747] = 12'hfff;
rom[6748] = 12'hfff;
rom[6749] = 12'hfff;
rom[6750] = 12'hfff;
rom[6751] = 12'hfff;
rom[6752] = 12'hfff;
rom[6753] = 12'hfff;
rom[6754] = 12'hfff;
rom[6755] = 12'hfff;
rom[6756] = 12'hfff;
rom[6757] = 12'hfff;
rom[6758] = 12'hfff;
rom[6759] = 12'hfff;
rom[6760] = 12'hfff;
rom[6761] = 12'hfff;
rom[6762] = 12'hfff;
rom[6763] = 12'hfff;
rom[6764] = 12'hfff;
rom[6765] = 12'hfff;
rom[6766] = 12'hfff;
rom[6767] = 12'hfff;
rom[6768] = 12'hfff;
rom[6769] = 12'hfff;
rom[6770] = 12'hfff;
rom[6771] = 12'hfff;
rom[6772] = 12'hfff;
rom[6773] = 12'hfff;
rom[6774] = 12'hfff;
rom[6775] = 12'hfff;
rom[6776] = 12'hfff;
rom[6777] = 12'hfff;
rom[6778] = 12'hfff;
rom[6779] = 12'hfff;
rom[6780] = 12'hfff;
rom[6781] = 12'hfff;
rom[6782] = 12'hfff;
rom[6783] = 12'hfff;
rom[6784] = 12'hfff;
rom[6785] = 12'hfff;
rom[6786] = 12'hfff;
rom[6787] = 12'hfff;
rom[6788] = 12'hfff;
rom[6789] = 12'hfff;
rom[6790] = 12'hfff;
rom[6791] = 12'hfff;
rom[6792] = 12'hfff;
rom[6793] = 12'hfff;
rom[6794] = 12'hfff;
rom[6795] = 12'hfff;
rom[6796] = 12'hfff;
rom[6797] = 12'hfff;
rom[6798] = 12'hfff;
rom[6799] = 12'hfff;
rom[6800] = 12'hfff;
rom[6801] = 12'hfff;
rom[6802] = 12'hfff;
rom[6803] = 12'hfff;
rom[6804] = 12'hfff;
rom[6805] = 12'hfff;
rom[6806] = 12'hfff;
rom[6807] = 12'hfff;
rom[6808] = 12'hfff;
rom[6809] = 12'hfff;
rom[6810] = 12'hfff;
rom[6811] = 12'hfff;
rom[6812] = 12'hfff;
rom[6813] = 12'hfff;
rom[6814] = 12'hfff;
rom[6815] = 12'hfff;
rom[6816] = 12'hfff;
rom[6817] = 12'hfff;
rom[6818] = 12'hfff;
rom[6819] = 12'hfff;
rom[6820] = 12'hfff;
rom[6821] = 12'hfff;
rom[6822] = 12'hfff;
rom[6823] = 12'hfff;
rom[6824] = 12'hfff;
rom[6825] = 12'hfff;
rom[6826] = 12'hfff;
rom[6827] = 12'hfff;
rom[6828] = 12'hfff;
rom[6829] = 12'hfff;
rom[6830] = 12'hfff;
rom[6831] = 12'hfff;
rom[6832] = 12'hfff;
rom[6833] = 12'hfff;
rom[6834] = 12'hfff;
rom[6835] = 12'hfff;
rom[6836] = 12'hfff;
rom[6837] = 12'hfff;
rom[6838] = 12'hfff;
rom[6839] = 12'hfff;
rom[6840] = 12'hfff;
rom[6841] = 12'hfff;
rom[6842] = 12'hfff;
rom[6843] = 12'hddf;
rom[6844] = 12'h22d;
rom[6845] = 12'h  c;
rom[6846] = 12'h  c;
rom[6847] = 12'h  c;
rom[6848] = 12'h  c;
rom[6849] = 12'h  c;
rom[6850] = 12'h11d;
rom[6851] = 12'hfff;
rom[6852] = 12'hfff;
rom[6853] = 12'h44d;
rom[6854] = 12'h  c;
rom[6855] = 12'h  c;
rom[6856] = 12'h  c;
rom[6857] = 12'h  c;
rom[6858] = 12'hbbf;
rom[6859] = 12'hfff;
rom[6860] = 12'hfff;
rom[6861] = 12'hfff;
rom[6862] = 12'hfff;
rom[6863] = 12'hfff;
rom[6864] = 12'hfff;
rom[6865] = 12'hfff;
rom[6866] = 12'hfff;
rom[6867] = 12'hfff;
rom[6868] = 12'hfff;
rom[6869] = 12'hfff;
rom[6870] = 12'hfff;
rom[6871] = 12'hfff;
rom[6872] = 12'hfff;
rom[6873] = 12'hfff;
rom[6874] = 12'hfff;
rom[6875] = 12'hfff;
rom[6876] = 12'hfff;
rom[6877] = 12'hfff;
rom[6878] = 12'hfff;
rom[6879] = 12'hfff;
rom[6880] = 12'hfff;
rom[6881] = 12'hfff;
rom[6882] = 12'hfff;
rom[6883] = 12'hfff;
rom[6884] = 12'hfff;
rom[6885] = 12'hfff;
rom[6886] = 12'hfff;
rom[6887] = 12'hfff;
rom[6888] = 12'hfff;
rom[6889] = 12'hfff;
rom[6890] = 12'hfff;
rom[6891] = 12'hfff;
rom[6892] = 12'hfff;
rom[6893] = 12'hfff;
rom[6894] = 12'hfff;
rom[6895] = 12'hfff;
rom[6896] = 12'hfff;
rom[6897] = 12'hfff;
rom[6898] = 12'hfff;
rom[6899] = 12'hfff;
rom[6900] = 12'hfff;
rom[6901] = 12'hfff;
rom[6902] = 12'hfff;
rom[6903] = 12'hfff;
rom[6904] = 12'hfff;
rom[6905] = 12'hfff;
rom[6906] = 12'hfff;
rom[6907] = 12'hfff;
rom[6908] = 12'hfff;
rom[6909] = 12'hfff;
rom[6910] = 12'hfff;
rom[6911] = 12'hfff;
rom[6912] = 12'hfff;
rom[6913] = 12'hfff;
rom[6914] = 12'hfff;
rom[6915] = 12'hfff;
rom[6916] = 12'hfff;
rom[6917] = 12'hfff;
rom[6918] = 12'hfff;
rom[6919] = 12'hfff;
rom[6920] = 12'hfff;
rom[6921] = 12'hfff;
rom[6922] = 12'hfff;
rom[6923] = 12'hfff;
rom[6924] = 12'hfff;
rom[6925] = 12'hfff;
rom[6926] = 12'hfff;
rom[6927] = 12'hfff;
rom[6928] = 12'hfff;
rom[6929] = 12'hfff;
rom[6930] = 12'hfff;
rom[6931] = 12'hfff;
rom[6932] = 12'hfff;
rom[6933] = 12'hfff;
rom[6934] = 12'hfff;
rom[6935] = 12'hfff;
rom[6936] = 12'hfff;
rom[6937] = 12'hfff;
rom[6938] = 12'hfff;
rom[6939] = 12'hfff;
rom[6940] = 12'hfff;
rom[6941] = 12'hfff;
rom[6942] = 12'hfff;
rom[6943] = 12'hfff;
rom[6944] = 12'hfff;
rom[6945] = 12'hfff;
rom[6946] = 12'hfff;
rom[6947] = 12'hfff;
rom[6948] = 12'hfff;
rom[6949] = 12'hfff;
rom[6950] = 12'hfff;
rom[6951] = 12'hfff;
rom[6952] = 12'hfff;
rom[6953] = 12'hfff;
rom[6954] = 12'hfff;
rom[6955] = 12'hfff;
rom[6956] = 12'hfff;
rom[6957] = 12'hfff;
rom[6958] = 12'hfff;
rom[6959] = 12'hfff;
rom[6960] = 12'hfff;
rom[6961] = 12'hfff;
rom[6962] = 12'hfff;
rom[6963] = 12'hfff;
rom[6964] = 12'hfff;
rom[6965] = 12'hfff;
rom[6966] = 12'hfff;
rom[6967] = 12'hfff;
rom[6968] = 12'hfff;
rom[6969] = 12'hfff;
rom[6970] = 12'hfff;
rom[6971] = 12'hfff;
rom[6972] = 12'heef;
rom[6973] = 12'h33d;
rom[6974] = 12'h  c;
rom[6975] = 12'h  c;
rom[6976] = 12'h  c;
rom[6977] = 12'h  c;
rom[6978] = 12'h  c;
rom[6979] = 12'haae;
rom[6980] = 12'hfff;
rom[6981] = 12'h44d;
rom[6982] = 12'h  c;
rom[6983] = 12'h  c;
rom[6984] = 12'h  c;
rom[6985] = 12'h  c;
rom[6986] = 12'hbbf;
rom[6987] = 12'hfff;
rom[6988] = 12'hfff;
rom[6989] = 12'hfff;
rom[6990] = 12'hfff;
rom[6991] = 12'hfff;
rom[6992] = 12'hfff;
rom[6993] = 12'hfff;
rom[6994] = 12'hfff;
rom[6995] = 12'hfff;
rom[6996] = 12'hfff;
rom[6997] = 12'hfff;
rom[6998] = 12'hfff;
rom[6999] = 12'hfff;
rom[7000] = 12'hfff;
rom[7001] = 12'hfff;
rom[7002] = 12'hfff;
rom[7003] = 12'hfff;
rom[7004] = 12'hfff;
rom[7005] = 12'hfff;
rom[7006] = 12'hfff;
rom[7007] = 12'hfff;
rom[7008] = 12'hfff;
rom[7009] = 12'hfff;
rom[7010] = 12'hfff;
rom[7011] = 12'hfff;
rom[7012] = 12'hfff;
rom[7013] = 12'hfff;
rom[7014] = 12'hfff;
rom[7015] = 12'hfff;
rom[7016] = 12'hfff;
rom[7017] = 12'hfff;
rom[7018] = 12'hfff;
rom[7019] = 12'hfff;
rom[7020] = 12'hfff;
rom[7021] = 12'hfff;
rom[7022] = 12'hfff;
rom[7023] = 12'hfff;
rom[7024] = 12'hfff;
rom[7025] = 12'hfff;
rom[7026] = 12'hfff;
rom[7027] = 12'hfff;
rom[7028] = 12'hfff;
rom[7029] = 12'hfff;
rom[7030] = 12'hfff;
rom[7031] = 12'hfff;
rom[7032] = 12'hfff;
rom[7033] = 12'hfff;
rom[7034] = 12'hfff;
rom[7035] = 12'hfff;
rom[7036] = 12'hfff;
rom[7037] = 12'hfff;
rom[7038] = 12'hfff;
rom[7039] = 12'hfff;
rom[7040] = 12'hfff;
rom[7041] = 12'hfff;
rom[7042] = 12'hfff;
rom[7043] = 12'hfff;
rom[7044] = 12'hfff;
rom[7045] = 12'hfff;
rom[7046] = 12'hfff;
rom[7047] = 12'hfff;
rom[7048] = 12'hfff;
rom[7049] = 12'hfff;
rom[7050] = 12'hfff;
rom[7051] = 12'hfff;
rom[7052] = 12'hfff;
rom[7053] = 12'hfff;
rom[7054] = 12'hfff;
rom[7055] = 12'hfff;
rom[7056] = 12'hfff;
rom[7057] = 12'hfff;
rom[7058] = 12'hfff;
rom[7059] = 12'hfff;
rom[7060] = 12'hfff;
rom[7061] = 12'hfff;
rom[7062] = 12'hfff;
rom[7063] = 12'hfff;
rom[7064] = 12'hfff;
rom[7065] = 12'hfff;
rom[7066] = 12'hfff;
rom[7067] = 12'hfff;
rom[7068] = 12'hfff;
rom[7069] = 12'hfff;
rom[7070] = 12'hfff;
rom[7071] = 12'hfff;
rom[7072] = 12'hfff;
rom[7073] = 12'hfff;
rom[7074] = 12'hfff;
rom[7075] = 12'hfff;
rom[7076] = 12'hfff;
rom[7077] = 12'hfff;
rom[7078] = 12'hfff;
rom[7079] = 12'hfff;
rom[7080] = 12'hfff;
rom[7081] = 12'hfff;
rom[7082] = 12'hfff;
rom[7083] = 12'hfff;
rom[7084] = 12'hfff;
rom[7085] = 12'hfff;
rom[7086] = 12'hfff;
rom[7087] = 12'hfff;
rom[7088] = 12'hfff;
rom[7089] = 12'hfff;
rom[7090] = 12'hfff;
rom[7091] = 12'hfff;
rom[7092] = 12'hfff;
rom[7093] = 12'hfff;
rom[7094] = 12'hfff;
rom[7095] = 12'hfff;
rom[7096] = 12'hfff;
rom[7097] = 12'hfff;
rom[7098] = 12'hfff;
rom[7099] = 12'hfff;
rom[7100] = 12'hfff;
rom[7101] = 12'hfff;
rom[7102] = 12'h44d;
rom[7103] = 12'h  c;
rom[7104] = 12'h  c;
rom[7105] = 12'h  c;
rom[7106] = 12'h  c;
rom[7107] = 12'h44d;
rom[7108] = 12'hfff;
rom[7109] = 12'h33d;
rom[7110] = 12'h  c;
rom[7111] = 12'h  c;
rom[7112] = 12'h  c;
rom[7113] = 12'h  c;
rom[7114] = 12'hccf;
rom[7115] = 12'hfff;
rom[7116] = 12'hfff;
rom[7117] = 12'hfff;
rom[7118] = 12'hfff;
rom[7119] = 12'hfff;
rom[7120] = 12'hfff;
rom[7121] = 12'hfff;
rom[7122] = 12'hfff;
rom[7123] = 12'hfff;
rom[7124] = 12'hfff;
rom[7125] = 12'hfff;
rom[7126] = 12'hfff;
rom[7127] = 12'hfff;
rom[7128] = 12'hfff;
rom[7129] = 12'hfff;
rom[7130] = 12'hfff;
rom[7131] = 12'hfff;
rom[7132] = 12'hfff;
rom[7133] = 12'hfff;
rom[7134] = 12'hfff;
rom[7135] = 12'hfff;
rom[7136] = 12'hfff;
rom[7137] = 12'hfff;
rom[7138] = 12'hfff;
rom[7139] = 12'hfff;
rom[7140] = 12'hfff;
rom[7141] = 12'hfff;
rom[7142] = 12'hfff;
rom[7143] = 12'hfff;
rom[7144] = 12'hfff;
rom[7145] = 12'hfff;
rom[7146] = 12'hfff;
rom[7147] = 12'hfff;
rom[7148] = 12'hfff;
rom[7149] = 12'hfff;
rom[7150] = 12'hfff;
rom[7151] = 12'hfff;
rom[7152] = 12'hfff;
rom[7153] = 12'hfff;
rom[7154] = 12'hfff;
rom[7155] = 12'hfff;
rom[7156] = 12'hfff;
rom[7157] = 12'hfff;
rom[7158] = 12'hfff;
rom[7159] = 12'hfff;
rom[7160] = 12'hfff;
rom[7161] = 12'hfff;
rom[7162] = 12'hfff;
rom[7163] = 12'hfff;
rom[7164] = 12'hfff;
rom[7165] = 12'hfff;
rom[7166] = 12'hfff;
rom[7167] = 12'hfff;
rom[7168] = 12'hfff;
rom[7169] = 12'hfff;
rom[7170] = 12'hfff;
rom[7171] = 12'hfff;
rom[7172] = 12'hfff;
rom[7173] = 12'hfff;
rom[7174] = 12'hfff;
rom[7175] = 12'hfff;
rom[7176] = 12'hfff;
rom[7177] = 12'hfff;
rom[7178] = 12'hfff;
rom[7179] = 12'hfff;
rom[7180] = 12'hfff;
rom[7181] = 12'hfff;
rom[7182] = 12'hfff;
rom[7183] = 12'hfff;
rom[7184] = 12'hfff;
rom[7185] = 12'hfff;
rom[7186] = 12'hfff;
rom[7187] = 12'hfff;
rom[7188] = 12'hfff;
rom[7189] = 12'hfff;
rom[7190] = 12'hfff;
rom[7191] = 12'hfff;
rom[7192] = 12'hfff;
rom[7193] = 12'hfff;
rom[7194] = 12'hfff;
rom[7195] = 12'hfff;
rom[7196] = 12'hfff;
rom[7197] = 12'hfff;
rom[7198] = 12'hfff;
rom[7199] = 12'hfff;
rom[7200] = 12'hfff;
rom[7201] = 12'hfff;
rom[7202] = 12'hfff;
rom[7203] = 12'hfff;
rom[7204] = 12'hfff;
rom[7205] = 12'hfff;
rom[7206] = 12'hfff;
rom[7207] = 12'hfff;
rom[7208] = 12'hfff;
rom[7209] = 12'hfff;
rom[7210] = 12'hfff;
rom[7211] = 12'hfff;
rom[7212] = 12'hfff;
rom[7213] = 12'hfff;
rom[7214] = 12'hfff;
rom[7215] = 12'hfff;
rom[7216] = 12'hfff;
rom[7217] = 12'hfff;
rom[7218] = 12'hfff;
rom[7219] = 12'hfff;
rom[7220] = 12'hfff;
rom[7221] = 12'hfff;
rom[7222] = 12'hfff;
rom[7223] = 12'hfff;
rom[7224] = 12'hfff;
rom[7225] = 12'hfff;
rom[7226] = 12'hfff;
rom[7227] = 12'hfff;
rom[7228] = 12'hfff;
rom[7229] = 12'hfff;
rom[7230] = 12'h99e;
rom[7231] = 12'h  c;
rom[7232] = 12'h  c;
rom[7233] = 12'h  c;
rom[7234] = 12'h  c;
rom[7235] = 12'h  c;
rom[7236] = 12'h33d;
rom[7237] = 12'h33d;
rom[7238] = 12'h  c;
rom[7239] = 12'h  c;
rom[7240] = 12'h  c;
rom[7241] = 12'h  c;
rom[7242] = 12'hccf;
rom[7243] = 12'hfff;
rom[7244] = 12'hfff;
rom[7245] = 12'hfff;
rom[7246] = 12'hfff;
rom[7247] = 12'hfff;
rom[7248] = 12'hfff;
rom[7249] = 12'hfff;
rom[7250] = 12'hfff;
rom[7251] = 12'hfff;
rom[7252] = 12'hfff;
rom[7253] = 12'hfff;
rom[7254] = 12'hfff;
rom[7255] = 12'hfff;
rom[7256] = 12'hfff;
rom[7257] = 12'hfff;
rom[7258] = 12'hfff;
rom[7259] = 12'hfff;
rom[7260] = 12'hfff;
rom[7261] = 12'hfff;
rom[7262] = 12'hfff;
rom[7263] = 12'hfff;
rom[7264] = 12'hfff;
rom[7265] = 12'hfff;
rom[7266] = 12'hfff;
rom[7267] = 12'hfff;
rom[7268] = 12'hfff;
rom[7269] = 12'hfff;
rom[7270] = 12'hfff;
rom[7271] = 12'hfff;
rom[7272] = 12'hfff;
rom[7273] = 12'hfff;
rom[7274] = 12'hfff;
rom[7275] = 12'hfff;
rom[7276] = 12'hfff;
rom[7277] = 12'hfff;
rom[7278] = 12'hfff;
rom[7279] = 12'hfff;
rom[7280] = 12'hfff;
rom[7281] = 12'hfff;
rom[7282] = 12'hfff;
rom[7283] = 12'hfff;
rom[7284] = 12'hfff;
rom[7285] = 12'hfff;
rom[7286] = 12'hfff;
rom[7287] = 12'hfff;
rom[7288] = 12'hfff;
rom[7289] = 12'hfff;
rom[7290] = 12'hfff;
rom[7291] = 12'hfff;
rom[7292] = 12'hfff;
rom[7293] = 12'hfff;
rom[7294] = 12'hfff;
rom[7295] = 12'hfff;
rom[7296] = 12'hfff;
rom[7297] = 12'hfff;
rom[7298] = 12'hfff;
rom[7299] = 12'hfff;
rom[7300] = 12'hfff;
rom[7301] = 12'hfff;
rom[7302] = 12'hfff;
rom[7303] = 12'hfff;
rom[7304] = 12'hfff;
rom[7305] = 12'hfff;
rom[7306] = 12'hfff;
rom[7307] = 12'hfff;
rom[7308] = 12'hfff;
rom[7309] = 12'hfff;
rom[7310] = 12'hfff;
rom[7311] = 12'hfff;
rom[7312] = 12'hfff;
rom[7313] = 12'hfff;
rom[7314] = 12'hfff;
rom[7315] = 12'hfff;
rom[7316] = 12'hfff;
rom[7317] = 12'hfff;
rom[7318] = 12'hfff;
rom[7319] = 12'hfff;
rom[7320] = 12'hfff;
rom[7321] = 12'hfff;
rom[7322] = 12'hfff;
rom[7323] = 12'hfff;
rom[7324] = 12'hfff;
rom[7325] = 12'hfff;
rom[7326] = 12'hfff;
rom[7327] = 12'hfff;
rom[7328] = 12'hfff;
rom[7329] = 12'hfff;
rom[7330] = 12'hfff;
rom[7331] = 12'hfff;
rom[7332] = 12'hfff;
rom[7333] = 12'hfff;
rom[7334] = 12'hfff;
rom[7335] = 12'hfff;
rom[7336] = 12'hfff;
rom[7337] = 12'hfff;
rom[7338] = 12'hfff;
rom[7339] = 12'hfff;
rom[7340] = 12'hfff;
rom[7341] = 12'hfff;
rom[7342] = 12'hfff;
rom[7343] = 12'hfff;
rom[7344] = 12'hfff;
rom[7345] = 12'hfff;
rom[7346] = 12'hfff;
rom[7347] = 12'hfff;
rom[7348] = 12'hfff;
rom[7349] = 12'hfff;
rom[7350] = 12'hfff;
rom[7351] = 12'hfff;
rom[7352] = 12'hfff;
rom[7353] = 12'hfff;
rom[7354] = 12'hfff;
rom[7355] = 12'hfff;
rom[7356] = 12'hfff;
rom[7357] = 12'hfff;
rom[7358] = 12'heef;
rom[7359] = 12'h11d;
rom[7360] = 12'h  c;
rom[7361] = 12'h  c;
rom[7362] = 12'h  c;
rom[7363] = 12'h  c;
rom[7364] = 12'h  c;
rom[7365] = 12'h  c;
rom[7366] = 12'h  c;
rom[7367] = 12'h  c;
rom[7368] = 12'h  c;
rom[7369] = 12'h  c;
rom[7370] = 12'hbbf;
rom[7371] = 12'hfff;
rom[7372] = 12'hfff;
rom[7373] = 12'hfff;
rom[7374] = 12'hfff;
rom[7375] = 12'hfff;
rom[7376] = 12'hfff;
rom[7377] = 12'hfff;
rom[7378] = 12'hfff;
rom[7379] = 12'hfff;
rom[7380] = 12'hfff;
rom[7381] = 12'hfff;
rom[7382] = 12'hfff;
rom[7383] = 12'hfff;
rom[7384] = 12'hfff;
rom[7385] = 12'hfff;
rom[7386] = 12'hfff;
rom[7387] = 12'hfff;
rom[7388] = 12'hfff;
rom[7389] = 12'hfff;
rom[7390] = 12'hfff;
rom[7391] = 12'hfff;
rom[7392] = 12'hfff;
rom[7393] = 12'hfff;
rom[7394] = 12'hfff;
rom[7395] = 12'hfff;
rom[7396] = 12'hfff;
rom[7397] = 12'hfff;
rom[7398] = 12'hfff;
rom[7399] = 12'hfff;
rom[7400] = 12'hfff;
rom[7401] = 12'hfff;
rom[7402] = 12'hfff;
rom[7403] = 12'hfff;
rom[7404] = 12'hfff;
rom[7405] = 12'hfff;
rom[7406] = 12'hfff;
rom[7407] = 12'hfff;
rom[7408] = 12'hfff;
rom[7409] = 12'hfff;
rom[7410] = 12'hfff;
rom[7411] = 12'hfff;
rom[7412] = 12'hfff;
rom[7413] = 12'hfff;
rom[7414] = 12'hfff;
rom[7415] = 12'hfff;
rom[7416] = 12'hfff;
rom[7417] = 12'hfff;
rom[7418] = 12'hfff;
rom[7419] = 12'hfff;
rom[7420] = 12'hfff;
rom[7421] = 12'hfff;
rom[7422] = 12'hfff;
rom[7423] = 12'hfff;
rom[7424] = 12'hfff;
rom[7425] = 12'hfff;
rom[7426] = 12'hfff;
rom[7427] = 12'hfff;
rom[7428] = 12'hfff;
rom[7429] = 12'hfff;
rom[7430] = 12'hfff;
rom[7431] = 12'hfff;
rom[7432] = 12'hfff;
rom[7433] = 12'hfff;
rom[7434] = 12'hfff;
rom[7435] = 12'hfff;
rom[7436] = 12'hfff;
rom[7437] = 12'hfff;
rom[7438] = 12'hfff;
rom[7439] = 12'hfff;
rom[7440] = 12'hfff;
rom[7441] = 12'hfff;
rom[7442] = 12'hfff;
rom[7443] = 12'hfff;
rom[7444] = 12'hfff;
rom[7445] = 12'hfff;
rom[7446] = 12'hfff;
rom[7447] = 12'hfff;
rom[7448] = 12'hfff;
rom[7449] = 12'hfff;
rom[7450] = 12'hfff;
rom[7451] = 12'hfff;
rom[7452] = 12'hfff;
rom[7453] = 12'hfff;
rom[7454] = 12'hfff;
rom[7455] = 12'hfff;
rom[7456] = 12'hfff;
rom[7457] = 12'hfff;
rom[7458] = 12'hfff;
rom[7459] = 12'hfff;
rom[7460] = 12'hfff;
rom[7461] = 12'hfff;
rom[7462] = 12'hfff;
rom[7463] = 12'hfff;
rom[7464] = 12'hfff;
rom[7465] = 12'hfff;
rom[7466] = 12'hfff;
rom[7467] = 12'hfff;
rom[7468] = 12'hfff;
rom[7469] = 12'hfff;
rom[7470] = 12'hfff;
rom[7471] = 12'hfff;
rom[7472] = 12'hfff;
rom[7473] = 12'hfff;
rom[7474] = 12'hfff;
rom[7475] = 12'hfff;
rom[7476] = 12'hfff;
rom[7477] = 12'hfff;
rom[7478] = 12'hfff;
rom[7479] = 12'hfff;
rom[7480] = 12'hfff;
rom[7481] = 12'hfff;
rom[7482] = 12'hfff;
rom[7483] = 12'hfff;
rom[7484] = 12'hfff;
rom[7485] = 12'hfff;
rom[7486] = 12'hfff;
rom[7487] = 12'hbbf;
rom[7488] = 12'h  c;
rom[7489] = 12'h  c;
rom[7490] = 12'h  c;
rom[7491] = 12'h  c;
rom[7492] = 12'h  c;
rom[7493] = 12'h  c;
rom[7494] = 12'h  c;
rom[7495] = 12'h  c;
rom[7496] = 12'h  c;
rom[7497] = 12'h  c;
rom[7498] = 12'hbbf;
rom[7499] = 12'hfff;
rom[7500] = 12'hfff;
rom[7501] = 12'hfff;
rom[7502] = 12'hfff;
rom[7503] = 12'hfff;
rom[7504] = 12'hfff;
rom[7505] = 12'hfff;
rom[7506] = 12'hfff;
rom[7507] = 12'hfff;
rom[7508] = 12'hfff;
rom[7509] = 12'hfff;
rom[7510] = 12'hfff;
rom[7511] = 12'hfff;
rom[7512] = 12'hfff;
rom[7513] = 12'hfff;
rom[7514] = 12'hfff;
rom[7515] = 12'hfff;
rom[7516] = 12'hfff;
rom[7517] = 12'hfff;
rom[7518] = 12'hfff;
rom[7519] = 12'hfff;
rom[7520] = 12'hfff;
rom[7521] = 12'hfff;
rom[7522] = 12'hfff;
rom[7523] = 12'hfff;
rom[7524] = 12'hfff;
rom[7525] = 12'hfff;
rom[7526] = 12'hfff;
rom[7527] = 12'hfff;
rom[7528] = 12'hfff;
rom[7529] = 12'hfff;
rom[7530] = 12'hfff;
rom[7531] = 12'hfff;
rom[7532] = 12'hfff;
rom[7533] = 12'hfff;
rom[7534] = 12'hfff;
rom[7535] = 12'hfff;
rom[7536] = 12'hfff;
rom[7537] = 12'hfff;
rom[7538] = 12'hfff;
rom[7539] = 12'hfff;
rom[7540] = 12'hfff;
rom[7541] = 12'hfff;
rom[7542] = 12'hfff;
rom[7543] = 12'hfff;
rom[7544] = 12'hfff;
rom[7545] = 12'hfff;
rom[7546] = 12'hfff;
rom[7547] = 12'hfff;
rom[7548] = 12'hfff;
rom[7549] = 12'hfff;
rom[7550] = 12'hfff;
rom[7551] = 12'hfff;
rom[7552] = 12'hfff;
rom[7553] = 12'hfff;
rom[7554] = 12'hfff;
rom[7555] = 12'hfff;
rom[7556] = 12'hfff;
rom[7557] = 12'hfff;
rom[7558] = 12'hfff;
rom[7559] = 12'hfff;
rom[7560] = 12'hfff;
rom[7561] = 12'hfff;
rom[7562] = 12'hfff;
rom[7563] = 12'hfff;
rom[7564] = 12'hfff;
rom[7565] = 12'hfff;
rom[7566] = 12'hfff;
rom[7567] = 12'hfff;
rom[7568] = 12'hfff;
rom[7569] = 12'hfff;
rom[7570] = 12'hfff;
rom[7571] = 12'hfff;
rom[7572] = 12'hfff;
rom[7573] = 12'hfff;
rom[7574] = 12'hfff;
rom[7575] = 12'hfff;
rom[7576] = 12'hfff;
rom[7577] = 12'hfff;
rom[7578] = 12'hfff;
rom[7579] = 12'hfff;
rom[7580] = 12'hfff;
rom[7581] = 12'hfff;
rom[7582] = 12'hfff;
rom[7583] = 12'hfff;
rom[7584] = 12'hfff;
rom[7585] = 12'hfff;
rom[7586] = 12'hfff;
rom[7587] = 12'hfff;
rom[7588] = 12'hfff;
rom[7589] = 12'hfff;
rom[7590] = 12'hfff;
rom[7591] = 12'hfff;
rom[7592] = 12'hfff;
rom[7593] = 12'hfff;
rom[7594] = 12'hfff;
rom[7595] = 12'hfff;
rom[7596] = 12'hfff;
rom[7597] = 12'hfff;
rom[7598] = 12'hfff;
rom[7599] = 12'hfff;
rom[7600] = 12'hfff;
rom[7601] = 12'hfff;
rom[7602] = 12'hfff;
rom[7603] = 12'hfff;
rom[7604] = 12'hfff;
rom[7605] = 12'hfff;
rom[7606] = 12'hfff;
rom[7607] = 12'hfff;
rom[7608] = 12'hfff;
rom[7609] = 12'hfff;
rom[7610] = 12'hfff;
rom[7611] = 12'hfff;
rom[7612] = 12'hfff;
rom[7613] = 12'hfff;
rom[7614] = 12'hfff;
rom[7615] = 12'hfff;
rom[7616] = 12'hbbf;
rom[7617] = 12'h  c;
rom[7618] = 12'h  c;
rom[7619] = 12'h  c;
rom[7620] = 12'h  c;
rom[7621] = 12'h  c;
rom[7622] = 12'h  c;
rom[7623] = 12'h  c;
rom[7624] = 12'h  c;
rom[7625] = 12'h  c;
rom[7626] = 12'hbbf;
rom[7627] = 12'hfff;
rom[7628] = 12'hfff;
rom[7629] = 12'hfff;
rom[7630] = 12'hfff;
rom[7631] = 12'hfff;
rom[7632] = 12'hfff;
rom[7633] = 12'hfff;
rom[7634] = 12'hfff;
rom[7635] = 12'hfff;
rom[7636] = 12'hfff;
rom[7637] = 12'hfff;
rom[7638] = 12'hfff;
rom[7639] = 12'hfff;
rom[7640] = 12'hfff;
rom[7641] = 12'hfff;
rom[7642] = 12'hfff;
rom[7643] = 12'hfff;
rom[7644] = 12'hfff;
rom[7645] = 12'hfff;
rom[7646] = 12'hfff;
rom[7647] = 12'hfff;
rom[7648] = 12'hfff;
rom[7649] = 12'hfff;
rom[7650] = 12'hfff;
rom[7651] = 12'hfff;
rom[7652] = 12'hfff;
rom[7653] = 12'hfff;
rom[7654] = 12'hfff;
rom[7655] = 12'hfff;
rom[7656] = 12'hfff;
rom[7657] = 12'hfff;
rom[7658] = 12'hfff;
rom[7659] = 12'hfff;
rom[7660] = 12'hfff;
rom[7661] = 12'hfff;
rom[7662] = 12'hfff;
rom[7663] = 12'hfff;
rom[7664] = 12'hfff;
rom[7665] = 12'hfff;
rom[7666] = 12'hfff;
rom[7667] = 12'hfff;
rom[7668] = 12'hfff;
rom[7669] = 12'hfff;
rom[7670] = 12'hfff;
rom[7671] = 12'hfff;
rom[7672] = 12'hfff;
rom[7673] = 12'hfff;
rom[7674] = 12'hfff;
rom[7675] = 12'hfff;
rom[7676] = 12'hfff;
rom[7677] = 12'hfff;
rom[7678] = 12'hfff;
rom[7679] = 12'hfff;
rom[7680] = 12'hfff;
rom[7681] = 12'hfff;
rom[7682] = 12'hfff;
rom[7683] = 12'hfff;
rom[7684] = 12'hfff;
rom[7685] = 12'hfff;
rom[7686] = 12'hfff;
rom[7687] = 12'hfff;
rom[7688] = 12'hfff;
rom[7689] = 12'hfff;
rom[7690] = 12'hfff;
rom[7691] = 12'hfff;
rom[7692] = 12'hfff;
rom[7693] = 12'hfff;
rom[7694] = 12'hfff;
rom[7695] = 12'hfff;
rom[7696] = 12'hfff;
rom[7697] = 12'hfff;
rom[7698] = 12'hfff;
rom[7699] = 12'hfff;
rom[7700] = 12'hfff;
rom[7701] = 12'hfff;
rom[7702] = 12'hfff;
rom[7703] = 12'hfff;
rom[7704] = 12'hfff;
rom[7705] = 12'hfff;
rom[7706] = 12'hfff;
rom[7707] = 12'hfff;
rom[7708] = 12'hfff;
rom[7709] = 12'hfff;
rom[7710] = 12'hfff;
rom[7711] = 12'hfff;
rom[7712] = 12'hfff;
rom[7713] = 12'hfff;
rom[7714] = 12'hfff;
rom[7715] = 12'hfff;
rom[7716] = 12'hfff;
rom[7717] = 12'hfff;
rom[7718] = 12'hfff;
rom[7719] = 12'hfff;
rom[7720] = 12'hfff;
rom[7721] = 12'hfff;
rom[7722] = 12'hfff;
rom[7723] = 12'hfff;
rom[7724] = 12'hfff;
rom[7725] = 12'hfff;
rom[7726] = 12'hfff;
rom[7727] = 12'hfff;
rom[7728] = 12'hfff;
rom[7729] = 12'hfff;
rom[7730] = 12'hfff;
rom[7731] = 12'hfff;
rom[7732] = 12'hfff;
rom[7733] = 12'hfff;
rom[7734] = 12'hfff;
rom[7735] = 12'hfff;
rom[7736] = 12'hfff;
rom[7737] = 12'hfff;
rom[7738] = 12'hfff;
rom[7739] = 12'hfff;
rom[7740] = 12'hfff;
rom[7741] = 12'hfff;
rom[7742] = 12'hfff;
rom[7743] = 12'hfff;
rom[7744] = 12'hfff;
rom[7745] = 12'hddf;
rom[7746] = 12'h22d;
rom[7747] = 12'h  c;
rom[7748] = 12'h  c;
rom[7749] = 12'h  c;
rom[7750] = 12'h  c;
rom[7751] = 12'h  c;
rom[7752] = 12'h  c;
rom[7753] = 12'h  c;
rom[7754] = 12'haae;
rom[7755] = 12'hfff;
rom[7756] = 12'hfff;
rom[7757] = 12'hfff;
rom[7758] = 12'hfff;
rom[7759] = 12'hfff;
rom[7760] = 12'hfff;
rom[7761] = 12'hfff;
rom[7762] = 12'hfff;
rom[7763] = 12'hfff;
rom[7764] = 12'hfff;
rom[7765] = 12'hfff;
rom[7766] = 12'hfff;
rom[7767] = 12'hfff;
rom[7768] = 12'hfff;
rom[7769] = 12'hfff;
rom[7770] = 12'hfff;
rom[7771] = 12'hfff;
rom[7772] = 12'hfff;
rom[7773] = 12'hfff;
rom[7774] = 12'hfff;
rom[7775] = 12'hfff;
rom[7776] = 12'hfff;
rom[7777] = 12'hfff;
rom[7778] = 12'hfff;
rom[7779] = 12'hfff;
rom[7780] = 12'hfff;
rom[7781] = 12'hfff;
rom[7782] = 12'hfff;
rom[7783] = 12'hfff;
rom[7784] = 12'hfff;
rom[7785] = 12'hfff;
rom[7786] = 12'hfff;
rom[7787] = 12'hfff;
rom[7788] = 12'hfff;
rom[7789] = 12'hfff;
rom[7790] = 12'hfff;
rom[7791] = 12'hfff;
rom[7792] = 12'hfff;
rom[7793] = 12'hfff;
rom[7794] = 12'hfff;
rom[7795] = 12'hfff;
rom[7796] = 12'hfff;
rom[7797] = 12'hfff;
rom[7798] = 12'hfff;
rom[7799] = 12'hfff;
rom[7800] = 12'hfff;
rom[7801] = 12'hfff;
rom[7802] = 12'hfff;
rom[7803] = 12'hfff;
rom[7804] = 12'hfff;
rom[7805] = 12'hfff;
rom[7806] = 12'hfff;
rom[7807] = 12'hfff;
rom[7808] = 12'hfff;
rom[7809] = 12'hfff;
rom[7810] = 12'hfff;
rom[7811] = 12'hfff;
rom[7812] = 12'hfff;
rom[7813] = 12'hfff;
rom[7814] = 12'hfff;
rom[7815] = 12'hfff;
rom[7816] = 12'hfff;
rom[7817] = 12'hfff;
rom[7818] = 12'hfff;
rom[7819] = 12'hfff;
rom[7820] = 12'hfff;
rom[7821] = 12'hfff;
rom[7822] = 12'hfff;
rom[7823] = 12'hfff;
rom[7824] = 12'hfff;
rom[7825] = 12'hfff;
rom[7826] = 12'hfff;
rom[7827] = 12'hfff;
rom[7828] = 12'hfff;
rom[7829] = 12'hfff;
rom[7830] = 12'hfff;
rom[7831] = 12'hfff;
rom[7832] = 12'hfff;
rom[7833] = 12'hfff;
rom[7834] = 12'hfff;
rom[7835] = 12'hfff;
rom[7836] = 12'hfff;
rom[7837] = 12'hfff;
rom[7838] = 12'hfff;
rom[7839] = 12'hfff;
rom[7840] = 12'hfff;
rom[7841] = 12'hfff;
rom[7842] = 12'hfff;
rom[7843] = 12'hfff;
rom[7844] = 12'hfff;
rom[7845] = 12'hfff;
rom[7846] = 12'hfff;
rom[7847] = 12'hfff;
rom[7848] = 12'hfff;
rom[7849] = 12'hfff;
rom[7850] = 12'hfff;
rom[7851] = 12'hfff;
rom[7852] = 12'hfff;
rom[7853] = 12'hfff;
rom[7854] = 12'hfff;
rom[7855] = 12'hfff;
rom[7856] = 12'hfff;
rom[7857] = 12'hfff;
rom[7858] = 12'hfff;
rom[7859] = 12'hfff;
rom[7860] = 12'hfff;
rom[7861] = 12'hfff;
rom[7862] = 12'hfff;
rom[7863] = 12'hfff;
rom[7864] = 12'hfff;
rom[7865] = 12'hfff;
rom[7866] = 12'hfff;
rom[7867] = 12'hfff;
rom[7868] = 12'hfff;
rom[7869] = 12'hfff;
rom[7870] = 12'hfff;
rom[7871] = 12'hfff;
rom[7872] = 12'hfff;
rom[7873] = 12'hfff;
rom[7874] = 12'hfff;
rom[7875] = 12'h99e;
rom[7876] = 12'h11d;
rom[7877] = 12'h  c;
rom[7878] = 12'h  c;
rom[7879] = 12'h  c;
rom[7880] = 12'h  c;
rom[7881] = 12'h  c;
rom[7882] = 12'h77e;
rom[7883] = 12'hfff;
rom[7884] = 12'hfff;
rom[7885] = 12'hfff;
rom[7886] = 12'hfff;
rom[7887] = 12'hfff;
rom[7888] = 12'hfff;
rom[7889] = 12'hfff;
rom[7890] = 12'hfff;
rom[7891] = 12'hfff;
rom[7892] = 12'hfff;
rom[7893] = 12'hfff;
rom[7894] = 12'hfff;
rom[7895] = 12'hfff;
rom[7896] = 12'hfff;
rom[7897] = 12'hfff;
rom[7898] = 12'hfff;
rom[7899] = 12'hfff;
rom[7900] = 12'hfff;
rom[7901] = 12'hfff;
rom[7902] = 12'hfff;
rom[7903] = 12'hfff;
rom[7904] = 12'hfff;
rom[7905] = 12'hfff;
rom[7906] = 12'hfff;
rom[7907] = 12'hfff;
rom[7908] = 12'hfff;
rom[7909] = 12'hfff;
rom[7910] = 12'hfff;
rom[7911] = 12'hfff;
rom[7912] = 12'hfff;
rom[7913] = 12'hfff;
rom[7914] = 12'hfff;
rom[7915] = 12'hfff;
rom[7916] = 12'hfff;
rom[7917] = 12'hfff;
rom[7918] = 12'hfff;
rom[7919] = 12'hfff;
rom[7920] = 12'hfff;
rom[7921] = 12'hfff;
rom[7922] = 12'hfff;
rom[7923] = 12'hfff;
rom[7924] = 12'hfff;
rom[7925] = 12'hfff;
rom[7926] = 12'hfff;
rom[7927] = 12'hfff;
rom[7928] = 12'hfff;
rom[7929] = 12'hfff;
rom[7930] = 12'hfff;
rom[7931] = 12'hfff;
rom[7932] = 12'hfff;
rom[7933] = 12'hfff;
rom[7934] = 12'hfff;
rom[7935] = 12'hfff;
rom[7936] = 12'hfff;
rom[7937] = 12'hfff;
rom[7938] = 12'hfff;
rom[7939] = 12'hfff;
rom[7940] = 12'hfff;
rom[7941] = 12'hfff;
rom[7942] = 12'hfff;
rom[7943] = 12'hfff;
rom[7944] = 12'hfff;
rom[7945] = 12'hfff;
rom[7946] = 12'hfff;
rom[7947] = 12'hfff;
rom[7948] = 12'hfff;
rom[7949] = 12'hfff;
rom[7950] = 12'hfff;
rom[7951] = 12'hfff;
rom[7952] = 12'hfff;
rom[7953] = 12'hfff;
rom[7954] = 12'hfff;
rom[7955] = 12'hfff;
rom[7956] = 12'hfff;
rom[7957] = 12'hfff;
rom[7958] = 12'hfff;
rom[7959] = 12'hfff;
rom[7960] = 12'hfff;
rom[7961] = 12'hfff;
rom[7962] = 12'hfff;
rom[7963] = 12'hfff;
rom[7964] = 12'hfff;
rom[7965] = 12'hfff;
rom[7966] = 12'hfff;
rom[7967] = 12'hfff;
rom[7968] = 12'hfff;
rom[7969] = 12'hfff;
rom[7970] = 12'hfff;
rom[7971] = 12'hfff;
rom[7972] = 12'hfff;
rom[7973] = 12'hfff;
rom[7974] = 12'hfff;
rom[7975] = 12'hfff;
rom[7976] = 12'hfff;
rom[7977] = 12'hfff;
rom[7978] = 12'hfff;
rom[7979] = 12'hfff;
rom[7980] = 12'hfff;
rom[7981] = 12'hfff;
rom[7982] = 12'hfff;
rom[7983] = 12'hfff;
rom[7984] = 12'hfff;
rom[7985] = 12'hfff;
rom[7986] = 12'hfff;
rom[7987] = 12'hfff;
rom[7988] = 12'hfff;
rom[7989] = 12'hfff;
rom[7990] = 12'hfff;
rom[7991] = 12'hfff;
rom[7992] = 12'hfff;
rom[7993] = 12'hfff;
rom[7994] = 12'hfff;
rom[7995] = 12'hfff;
rom[7996] = 12'hfff;
rom[7997] = 12'hfff;
rom[7998] = 12'hfff;
rom[7999] = 12'hfff;
rom[8000] = 12'hfff;
rom[8001] = 12'hfff;
rom[8002] = 12'hfff;
rom[8003] = 12'hfff;
rom[8004] = 12'heef;
rom[8005] = 12'h11d;
rom[8006] = 12'h  c;
rom[8007] = 12'h  c;
rom[8008] = 12'h  c;
rom[8009] = 12'h  c;
rom[8010] = 12'h33d;
rom[8011] = 12'hfff;
rom[8012] = 12'hfff;
rom[8013] = 12'hfff;
rom[8014] = 12'hfff;
rom[8015] = 12'hfff;
rom[8016] = 12'hfff;
rom[8017] = 12'hfff;
rom[8018] = 12'hfff;
rom[8019] = 12'hfff;
rom[8020] = 12'hfff;
rom[8021] = 12'hfff;
rom[8022] = 12'hfff;
rom[8023] = 12'hfff;
rom[8024] = 12'hfff;
rom[8025] = 12'hfff;
rom[8026] = 12'hfff;
rom[8027] = 12'hfff;
rom[8028] = 12'hfff;
rom[8029] = 12'hfff;
rom[8030] = 12'hfff;
rom[8031] = 12'hfff;
rom[8032] = 12'hfff;
rom[8033] = 12'hfff;
rom[8034] = 12'hfff;
rom[8035] = 12'hfff;
rom[8036] = 12'hfff;
rom[8037] = 12'hfff;
rom[8038] = 12'hfff;
rom[8039] = 12'hfff;
rom[8040] = 12'hfff;
rom[8041] = 12'hfff;
rom[8042] = 12'hfff;
rom[8043] = 12'hfff;
rom[8044] = 12'hfff;
rom[8045] = 12'hfff;
rom[8046] = 12'hfff;
rom[8047] = 12'hfff;
rom[8048] = 12'hfff;
rom[8049] = 12'hfff;
rom[8050] = 12'hfff;
rom[8051] = 12'hfff;
rom[8052] = 12'hfff;
rom[8053] = 12'hfff;
rom[8054] = 12'hfff;
rom[8055] = 12'hfff;
rom[8056] = 12'hfff;
rom[8057] = 12'hfff;
rom[8058] = 12'hfff;
rom[8059] = 12'hfff;
rom[8060] = 12'hfff;
rom[8061] = 12'hfff;
rom[8062] = 12'hfff;
rom[8063] = 12'hfff;
rom[8064] = 12'hfff;
rom[8065] = 12'hfff;
rom[8066] = 12'hfff;
rom[8067] = 12'hfff;
rom[8068] = 12'hfff;
rom[8069] = 12'hfff;
rom[8070] = 12'hfff;
rom[8071] = 12'hfff;
rom[8072] = 12'hfff;
rom[8073] = 12'hfff;
rom[8074] = 12'hfff;
rom[8075] = 12'hfff;
rom[8076] = 12'hfff;
rom[8077] = 12'hfff;
rom[8078] = 12'hfff;
rom[8079] = 12'hfff;
rom[8080] = 12'hfff;
rom[8081] = 12'hfff;
rom[8082] = 12'hfff;
rom[8083] = 12'hfff;
rom[8084] = 12'hfff;
rom[8085] = 12'hfff;
rom[8086] = 12'hfff;
rom[8087] = 12'hfff;
rom[8088] = 12'hfff;
rom[8089] = 12'hfff;
rom[8090] = 12'hfff;
rom[8091] = 12'hfff;
rom[8092] = 12'hfff;
rom[8093] = 12'hfff;
rom[8094] = 12'hfff;
rom[8095] = 12'hfff;
rom[8096] = 12'hfff;
rom[8097] = 12'hfff;
rom[8098] = 12'hfff;
rom[8099] = 12'hfff;
rom[8100] = 12'hfff;
rom[8101] = 12'hfff;
rom[8102] = 12'hfff;
rom[8103] = 12'hfff;
rom[8104] = 12'hfff;
rom[8105] = 12'hfff;
rom[8106] = 12'hfff;
rom[8107] = 12'hfff;
rom[8108] = 12'hfff;
rom[8109] = 12'hfff;
rom[8110] = 12'hfff;
rom[8111] = 12'hfff;
rom[8112] = 12'hfff;
rom[8113] = 12'hfff;
rom[8114] = 12'hfff;
rom[8115] = 12'hfff;
rom[8116] = 12'hfff;
rom[8117] = 12'hfff;
rom[8118] = 12'hfff;
rom[8119] = 12'hfff;
rom[8120] = 12'hfff;
rom[8121] = 12'hfff;
rom[8122] = 12'hfff;
rom[8123] = 12'hfff;
rom[8124] = 12'hfff;
rom[8125] = 12'hfff;
rom[8126] = 12'hfff;
rom[8127] = 12'hfff;
rom[8128] = 12'hfff;
rom[8129] = 12'hfff;
rom[8130] = 12'hfff;
rom[8131] = 12'hfff;
rom[8132] = 12'hfff;
rom[8133] = 12'h44d;
rom[8134] = 12'h  c;
rom[8135] = 12'h  c;
rom[8136] = 12'h  c;
rom[8137] = 12'h  c;
rom[8138] = 12'h  c;
rom[8139] = 12'h44d;
rom[8140] = 12'haae;
rom[8141] = 12'heef;
rom[8142] = 12'hfff;
rom[8143] = 12'hfff;
rom[8144] = 12'hfff;
rom[8145] = 12'hfff;
rom[8146] = 12'hfff;
rom[8147] = 12'hfff;
rom[8148] = 12'hfff;
rom[8149] = 12'hfff;
rom[8150] = 12'hfff;
rom[8151] = 12'hfff;
rom[8152] = 12'hfff;
rom[8153] = 12'hfff;
rom[8154] = 12'hfff;
rom[8155] = 12'hfff;
rom[8156] = 12'hfff;
rom[8157] = 12'hfff;
rom[8158] = 12'hfff;
rom[8159] = 12'hfff;
rom[8160] = 12'hfff;
rom[8161] = 12'hfff;
rom[8162] = 12'hfff;
rom[8163] = 12'hfff;
rom[8164] = 12'hfff;
rom[8165] = 12'hfff;
rom[8166] = 12'hfff;
rom[8167] = 12'hfff;
rom[8168] = 12'hfff;
rom[8169] = 12'hfff;
rom[8170] = 12'hfff;
rom[8171] = 12'hfff;
rom[8172] = 12'hfff;
rom[8173] = 12'hfff;
rom[8174] = 12'hfff;
rom[8175] = 12'hfff;
rom[8176] = 12'hfff;
rom[8177] = 12'hfff;
rom[8178] = 12'hfff;
rom[8179] = 12'hfff;
rom[8180] = 12'hfff;
rom[8181] = 12'hfff;
rom[8182] = 12'hfff;
rom[8183] = 12'hfff;
rom[8184] = 12'hfff;
rom[8185] = 12'hfff;
rom[8186] = 12'hfff;
rom[8187] = 12'hfff;
rom[8188] = 12'hfff;
rom[8189] = 12'hfff;
rom[8190] = 12'hfff;
rom[8191] = 12'h99e;
rom[8192] = 12'hfff;
rom[8193] = 12'hfff;
rom[8194] = 12'hfff;
rom[8195] = 12'hfff;
rom[8196] = 12'hfff;
rom[8197] = 12'hfff;
rom[8198] = 12'hfff;
rom[8199] = 12'hfff;
rom[8200] = 12'hfff;
rom[8201] = 12'hfff;
rom[8202] = 12'hfff;
rom[8203] = 12'hfff;
rom[8204] = 12'hfff;
rom[8205] = 12'hfff;
rom[8206] = 12'hfff;
rom[8207] = 12'hfff;
rom[8208] = 12'hfff;
rom[8209] = 12'hfff;
rom[8210] = 12'hfff;
rom[8211] = 12'hfff;
rom[8212] = 12'hfff;
rom[8213] = 12'hfff;
rom[8214] = 12'hfff;
rom[8215] = 12'hfff;
rom[8216] = 12'hfff;
rom[8217] = 12'hfff;
rom[8218] = 12'hfff;
rom[8219] = 12'hfff;
rom[8220] = 12'hfff;
rom[8221] = 12'hfff;
rom[8222] = 12'hfff;
rom[8223] = 12'hfff;
rom[8224] = 12'hfff;
rom[8225] = 12'hfff;
rom[8226] = 12'hfff;
rom[8227] = 12'hfff;
rom[8228] = 12'hfff;
rom[8229] = 12'hfff;
rom[8230] = 12'hfff;
rom[8231] = 12'hfff;
rom[8232] = 12'hfff;
rom[8233] = 12'hfff;
rom[8234] = 12'hfff;
rom[8235] = 12'hfff;
rom[8236] = 12'hfff;
rom[8237] = 12'hfff;
rom[8238] = 12'hfff;
rom[8239] = 12'hfff;
rom[8240] = 12'hfff;
rom[8241] = 12'hfff;
rom[8242] = 12'hfff;
rom[8243] = 12'hfff;
rom[8244] = 12'hfff;
rom[8245] = 12'hfff;
rom[8246] = 12'hfff;
rom[8247] = 12'hfff;
rom[8248] = 12'hfff;
rom[8249] = 12'hfff;
rom[8250] = 12'hfff;
rom[8251] = 12'hfff;
rom[8252] = 12'hfff;
rom[8253] = 12'hfff;
rom[8254] = 12'hfff;
rom[8255] = 12'hfff;
rom[8256] = 12'hfff;
rom[8257] = 12'hfff;
rom[8258] = 12'hfff;
rom[8259] = 12'hfff;
rom[8260] = 12'hfff;
rom[8261] = 12'h99e;
rom[8262] = 12'h  c;
rom[8263] = 12'h  c;
rom[8264] = 12'h  c;
rom[8265] = 12'h  c;
rom[8266] = 12'h  c;
rom[8267] = 12'h  c;
rom[8268] = 12'h  c;
rom[8269] = 12'h11d;
rom[8270] = 12'hddf;
rom[8271] = 12'hfff;
rom[8272] = 12'hfff;
rom[8273] = 12'hfff;
rom[8274] = 12'hfff;
rom[8275] = 12'hfff;
rom[8276] = 12'hfff;
rom[8277] = 12'hfff;
rom[8278] = 12'hfff;
rom[8279] = 12'hfff;
rom[8280] = 12'hfff;
rom[8281] = 12'hfff;
rom[8282] = 12'hfff;
rom[8283] = 12'hfff;
rom[8284] = 12'hfff;
rom[8285] = 12'hfff;
rom[8286] = 12'hfff;
rom[8287] = 12'hfff;
rom[8288] = 12'hfff;
rom[8289] = 12'hfff;
rom[8290] = 12'hfff;
rom[8291] = 12'hfff;
rom[8292] = 12'hfff;
rom[8293] = 12'hfff;
rom[8294] = 12'hfff;
rom[8295] = 12'hfff;
rom[8296] = 12'hfff;
rom[8297] = 12'hfff;
rom[8298] = 12'hfff;
rom[8299] = 12'hfff;
rom[8300] = 12'hfff;
rom[8301] = 12'hfff;
rom[8302] = 12'hfff;
rom[8303] = 12'hfff;
rom[8304] = 12'hfff;
rom[8305] = 12'hfff;
rom[8306] = 12'hfff;
rom[8307] = 12'hfff;
rom[8308] = 12'hfff;
rom[8309] = 12'hfff;
rom[8310] = 12'hfff;
rom[8311] = 12'hfff;
rom[8312] = 12'hfff;
rom[8313] = 12'hfff;
rom[8314] = 12'hfff;
rom[8315] = 12'hfff;
rom[8316] = 12'hfff;
rom[8317] = 12'hfff;
rom[8318] = 12'heef;
rom[8319] = 12'h11d;
rom[8320] = 12'hfff;
rom[8321] = 12'hfff;
rom[8322] = 12'hfff;
rom[8323] = 12'hfff;
rom[8324] = 12'hfff;
rom[8325] = 12'hfff;
rom[8326] = 12'hfff;
rom[8327] = 12'hfff;
rom[8328] = 12'hfff;
rom[8329] = 12'hfff;
rom[8330] = 12'hfff;
rom[8331] = 12'hfff;
rom[8332] = 12'hfff;
rom[8333] = 12'hfff;
rom[8334] = 12'hfff;
rom[8335] = 12'hfff;
rom[8336] = 12'hfff;
rom[8337] = 12'hfff;
rom[8338] = 12'hfff;
rom[8339] = 12'hfff;
rom[8340] = 12'hfff;
rom[8341] = 12'hfff;
rom[8342] = 12'hfff;
rom[8343] = 12'hfff;
rom[8344] = 12'hfff;
rom[8345] = 12'hfff;
rom[8346] = 12'hfff;
rom[8347] = 12'hfff;
rom[8348] = 12'hfff;
rom[8349] = 12'hfff;
rom[8350] = 12'hfff;
rom[8351] = 12'hfff;
rom[8352] = 12'hfff;
rom[8353] = 12'hfff;
rom[8354] = 12'hfff;
rom[8355] = 12'hfff;
rom[8356] = 12'hfff;
rom[8357] = 12'hfff;
rom[8358] = 12'hfff;
rom[8359] = 12'hfff;
rom[8360] = 12'hfff;
rom[8361] = 12'hfff;
rom[8362] = 12'hfff;
rom[8363] = 12'hfff;
rom[8364] = 12'hfff;
rom[8365] = 12'hfff;
rom[8366] = 12'hfff;
rom[8367] = 12'hfff;
rom[8368] = 12'hfff;
rom[8369] = 12'hfff;
rom[8370] = 12'hfff;
rom[8371] = 12'hfff;
rom[8372] = 12'hfff;
rom[8373] = 12'hfff;
rom[8374] = 12'hfff;
rom[8375] = 12'hfff;
rom[8376] = 12'hfff;
rom[8377] = 12'hfff;
rom[8378] = 12'hfff;
rom[8379] = 12'hfff;
rom[8380] = 12'hfff;
rom[8381] = 12'hfff;
rom[8382] = 12'hfff;
rom[8383] = 12'hfff;
rom[8384] = 12'hfff;
rom[8385] = 12'hfff;
rom[8386] = 12'hfff;
rom[8387] = 12'hfff;
rom[8388] = 12'hfff;
rom[8389] = 12'hccf;
rom[8390] = 12'h  c;
rom[8391] = 12'h  c;
rom[8392] = 12'h  c;
rom[8393] = 12'h  c;
rom[8394] = 12'h  c;
rom[8395] = 12'h  c;
rom[8396] = 12'h  c;
rom[8397] = 12'h  c;
rom[8398] = 12'h  c;
rom[8399] = 12'h55d;
rom[8400] = 12'hccf;
rom[8401] = 12'heef;
rom[8402] = 12'hfff;
rom[8403] = 12'hfff;
rom[8404] = 12'hfff;
rom[8405] = 12'hfff;
rom[8406] = 12'hfff;
rom[8407] = 12'hfff;
rom[8408] = 12'hfff;
rom[8409] = 12'hfff;
rom[8410] = 12'hfff;
rom[8411] = 12'hfff;
rom[8412] = 12'hfff;
rom[8413] = 12'hfff;
rom[8414] = 12'hfff;
rom[8415] = 12'hfff;
rom[8416] = 12'hfff;
rom[8417] = 12'hfff;
rom[8418] = 12'hfff;
rom[8419] = 12'hfff;
rom[8420] = 12'hfff;
rom[8421] = 12'hfff;
rom[8422] = 12'hfff;
rom[8423] = 12'hfff;
rom[8424] = 12'hfff;
rom[8425] = 12'hfff;
rom[8426] = 12'hfff;
rom[8427] = 12'hfff;
rom[8428] = 12'hfff;
rom[8429] = 12'hfff;
rom[8430] = 12'hfff;
rom[8431] = 12'hfff;
rom[8432] = 12'hfff;
rom[8433] = 12'hfff;
rom[8434] = 12'hfff;
rom[8435] = 12'hfff;
rom[8436] = 12'hfff;
rom[8437] = 12'hfff;
rom[8438] = 12'hfff;
rom[8439] = 12'hfff;
rom[8440] = 12'hfff;
rom[8441] = 12'hfff;
rom[8442] = 12'hfff;
rom[8443] = 12'hfff;
rom[8444] = 12'hfff;
rom[8445] = 12'hfff;
rom[8446] = 12'h88e;
rom[8447] = 12'h  c;
rom[8448] = 12'hfff;
rom[8449] = 12'hfff;
rom[8450] = 12'hfff;
rom[8451] = 12'hfff;
rom[8452] = 12'hfff;
rom[8453] = 12'hfff;
rom[8454] = 12'hfff;
rom[8455] = 12'hfff;
rom[8456] = 12'hfff;
rom[8457] = 12'hfff;
rom[8458] = 12'hfff;
rom[8459] = 12'hfff;
rom[8460] = 12'hfff;
rom[8461] = 12'hfff;
rom[8462] = 12'hfff;
rom[8463] = 12'hfff;
rom[8464] = 12'hfff;
rom[8465] = 12'hfff;
rom[8466] = 12'hfff;
rom[8467] = 12'hfff;
rom[8468] = 12'hfff;
rom[8469] = 12'hfff;
rom[8470] = 12'hfff;
rom[8471] = 12'hfff;
rom[8472] = 12'hfff;
rom[8473] = 12'hfff;
rom[8474] = 12'hfff;
rom[8475] = 12'hfff;
rom[8476] = 12'hfff;
rom[8477] = 12'hfff;
rom[8478] = 12'hfff;
rom[8479] = 12'hfff;
rom[8480] = 12'hfff;
rom[8481] = 12'hfff;
rom[8482] = 12'hfff;
rom[8483] = 12'hfff;
rom[8484] = 12'hfff;
rom[8485] = 12'hfff;
rom[8486] = 12'hfff;
rom[8487] = 12'hfff;
rom[8488] = 12'hfff;
rom[8489] = 12'hfff;
rom[8490] = 12'hfff;
rom[8491] = 12'hfff;
rom[8492] = 12'hfff;
rom[8493] = 12'hfff;
rom[8494] = 12'hfff;
rom[8495] = 12'hfff;
rom[8496] = 12'hfff;
rom[8497] = 12'hfff;
rom[8498] = 12'hfff;
rom[8499] = 12'hfff;
rom[8500] = 12'hfff;
rom[8501] = 12'hfff;
rom[8502] = 12'hfff;
rom[8503] = 12'hfff;
rom[8504] = 12'hfff;
rom[8505] = 12'hfff;
rom[8506] = 12'hfff;
rom[8507] = 12'hfff;
rom[8508] = 12'hfff;
rom[8509] = 12'hfff;
rom[8510] = 12'hfff;
rom[8511] = 12'hfff;
rom[8512] = 12'hfff;
rom[8513] = 12'hfff;
rom[8514] = 12'hfff;
rom[8515] = 12'hfff;
rom[8516] = 12'hfff;
rom[8517] = 12'heef;
rom[8518] = 12'h  c;
rom[8519] = 12'h  c;
rom[8520] = 12'h  c;
rom[8521] = 12'h  c;
rom[8522] = 12'h  c;
rom[8523] = 12'h  c;
rom[8524] = 12'h  c;
rom[8525] = 12'h  c;
rom[8526] = 12'h44d;
rom[8527] = 12'h11d;
rom[8528] = 12'h  c;
rom[8529] = 12'h22d;
rom[8530] = 12'hfff;
rom[8531] = 12'hfff;
rom[8532] = 12'hfff;
rom[8533] = 12'hfff;
rom[8534] = 12'hfff;
rom[8535] = 12'hfff;
rom[8536] = 12'hfff;
rom[8537] = 12'hfff;
rom[8538] = 12'hfff;
rom[8539] = 12'hfff;
rom[8540] = 12'hfff;
rom[8541] = 12'hfff;
rom[8542] = 12'hfff;
rom[8543] = 12'hfff;
rom[8544] = 12'hfff;
rom[8545] = 12'hfff;
rom[8546] = 12'hfff;
rom[8547] = 12'hfff;
rom[8548] = 12'hfff;
rom[8549] = 12'hfff;
rom[8550] = 12'hfff;
rom[8551] = 12'hfff;
rom[8552] = 12'hfff;
rom[8553] = 12'hfff;
rom[8554] = 12'hfff;
rom[8555] = 12'hfff;
rom[8556] = 12'hfff;
rom[8557] = 12'hfff;
rom[8558] = 12'hfff;
rom[8559] = 12'hfff;
rom[8560] = 12'hfff;
rom[8561] = 12'hfff;
rom[8562] = 12'hfff;
rom[8563] = 12'hfff;
rom[8564] = 12'hfff;
rom[8565] = 12'hfff;
rom[8566] = 12'hfff;
rom[8567] = 12'hfff;
rom[8568] = 12'hfff;
rom[8569] = 12'hfff;
rom[8570] = 12'hfff;
rom[8571] = 12'hfff;
rom[8572] = 12'hfff;
rom[8573] = 12'heef;
rom[8574] = 12'h11d;
rom[8575] = 12'h  c;
rom[8576] = 12'hfff;
rom[8577] = 12'hfff;
rom[8578] = 12'hfff;
rom[8579] = 12'hfff;
rom[8580] = 12'hfff;
rom[8581] = 12'hfff;
rom[8582] = 12'hfff;
rom[8583] = 12'hfff;
rom[8584] = 12'hfff;
rom[8585] = 12'hfff;
rom[8586] = 12'hfff;
rom[8587] = 12'hfff;
rom[8588] = 12'hfff;
rom[8589] = 12'hfff;
rom[8590] = 12'hfff;
rom[8591] = 12'hfff;
rom[8592] = 12'hfff;
rom[8593] = 12'hfff;
rom[8594] = 12'hfff;
rom[8595] = 12'hfff;
rom[8596] = 12'hfff;
rom[8597] = 12'hfff;
rom[8598] = 12'hfff;
rom[8599] = 12'hfff;
rom[8600] = 12'hfff;
rom[8601] = 12'hfff;
rom[8602] = 12'hfff;
rom[8603] = 12'hfff;
rom[8604] = 12'hfff;
rom[8605] = 12'hfff;
rom[8606] = 12'hfff;
rom[8607] = 12'hfff;
rom[8608] = 12'hfff;
rom[8609] = 12'hfff;
rom[8610] = 12'hfff;
rom[8611] = 12'hfff;
rom[8612] = 12'hfff;
rom[8613] = 12'hfff;
rom[8614] = 12'hfff;
rom[8615] = 12'hfff;
rom[8616] = 12'hfff;
rom[8617] = 12'hfff;
rom[8618] = 12'hfff;
rom[8619] = 12'hfff;
rom[8620] = 12'hfff;
rom[8621] = 12'hfff;
rom[8622] = 12'hfff;
rom[8623] = 12'hfff;
rom[8624] = 12'hfff;
rom[8625] = 12'hfff;
rom[8626] = 12'hfff;
rom[8627] = 12'hfff;
rom[8628] = 12'hfff;
rom[8629] = 12'hfff;
rom[8630] = 12'hfff;
rom[8631] = 12'hfff;
rom[8632] = 12'hfff;
rom[8633] = 12'hfff;
rom[8634] = 12'hfff;
rom[8635] = 12'hfff;
rom[8636] = 12'hfff;
rom[8637] = 12'hfff;
rom[8638] = 12'hfff;
rom[8639] = 12'hfff;
rom[8640] = 12'hfff;
rom[8641] = 12'hfff;
rom[8642] = 12'hfff;
rom[8643] = 12'hfff;
rom[8644] = 12'hfff;
rom[8645] = 12'hfff;
rom[8646] = 12'h11d;
rom[8647] = 12'h  c;
rom[8648] = 12'h  c;
rom[8649] = 12'h  c;
rom[8650] = 12'h  c;
rom[8651] = 12'h  c;
rom[8652] = 12'h  c;
rom[8653] = 12'h  c;
rom[8654] = 12'h  c;
rom[8655] = 12'h  c;
rom[8656] = 12'h  c;
rom[8657] = 12'h  c;
rom[8658] = 12'h77e;
rom[8659] = 12'hfff;
rom[8660] = 12'hfff;
rom[8661] = 12'hfff;
rom[8662] = 12'hfff;
rom[8663] = 12'hfff;
rom[8664] = 12'hfff;
rom[8665] = 12'hfff;
rom[8666] = 12'hfff;
rom[8667] = 12'hfff;
rom[8668] = 12'hfff;
rom[8669] = 12'hfff;
rom[8670] = 12'hfff;
rom[8671] = 12'hfff;
rom[8672] = 12'hfff;
rom[8673] = 12'hfff;
rom[8674] = 12'hfff;
rom[8675] = 12'hfff;
rom[8676] = 12'hfff;
rom[8677] = 12'hfff;
rom[8678] = 12'hfff;
rom[8679] = 12'hfff;
rom[8680] = 12'hfff;
rom[8681] = 12'hfff;
rom[8682] = 12'hfff;
rom[8683] = 12'hfff;
rom[8684] = 12'hfff;
rom[8685] = 12'hfff;
rom[8686] = 12'hfff;
rom[8687] = 12'hfff;
rom[8688] = 12'hfff;
rom[8689] = 12'hfff;
rom[8690] = 12'hfff;
rom[8691] = 12'hfff;
rom[8692] = 12'hfff;
rom[8693] = 12'hfff;
rom[8694] = 12'hfff;
rom[8695] = 12'hfff;
rom[8696] = 12'hfff;
rom[8697] = 12'hfff;
rom[8698] = 12'hfff;
rom[8699] = 12'hfff;
rom[8700] = 12'heef;
rom[8701] = 12'h33d;
rom[8702] = 12'h  c;
rom[8703] = 12'h  c;
rom[8704] = 12'hfff;
rom[8705] = 12'hfff;
rom[8706] = 12'hfff;
rom[8707] = 12'hfff;
rom[8708] = 12'hfff;
rom[8709] = 12'hfff;
rom[8710] = 12'hfff;
rom[8711] = 12'hfff;
rom[8712] = 12'hfff;
rom[8713] = 12'hfff;
rom[8714] = 12'hfff;
rom[8715] = 12'hfff;
rom[8716] = 12'hfff;
rom[8717] = 12'hfff;
rom[8718] = 12'hfff;
rom[8719] = 12'hfff;
rom[8720] = 12'hfff;
rom[8721] = 12'hfff;
rom[8722] = 12'hfff;
rom[8723] = 12'hfff;
rom[8724] = 12'hfff;
rom[8725] = 12'hfff;
rom[8726] = 12'hfff;
rom[8727] = 12'hfff;
rom[8728] = 12'hfff;
rom[8729] = 12'hfff;
rom[8730] = 12'hfff;
rom[8731] = 12'hfff;
rom[8732] = 12'hfff;
rom[8733] = 12'hfff;
rom[8734] = 12'hfff;
rom[8735] = 12'hfff;
rom[8736] = 12'hfff;
rom[8737] = 12'hfff;
rom[8738] = 12'hfff;
rom[8739] = 12'hfff;
rom[8740] = 12'hfff;
rom[8741] = 12'hfff;
rom[8742] = 12'hfff;
rom[8743] = 12'hfff;
rom[8744] = 12'hfff;
rom[8745] = 12'hfff;
rom[8746] = 12'hfff;
rom[8747] = 12'hfff;
rom[8748] = 12'hfff;
rom[8749] = 12'hfff;
rom[8750] = 12'hfff;
rom[8751] = 12'hfff;
rom[8752] = 12'hfff;
rom[8753] = 12'hfff;
rom[8754] = 12'hfff;
rom[8755] = 12'hfff;
rom[8756] = 12'hfff;
rom[8757] = 12'hfff;
rom[8758] = 12'hfff;
rom[8759] = 12'hfff;
rom[8760] = 12'hfff;
rom[8761] = 12'hfff;
rom[8762] = 12'hfff;
rom[8763] = 12'hfff;
rom[8764] = 12'hfff;
rom[8765] = 12'hfff;
rom[8766] = 12'hfff;
rom[8767] = 12'hfff;
rom[8768] = 12'hfff;
rom[8769] = 12'hfff;
rom[8770] = 12'hfff;
rom[8771] = 12'hfff;
rom[8772] = 12'hfff;
rom[8773] = 12'hfff;
rom[8774] = 12'h77e;
rom[8775] = 12'h  c;
rom[8776] = 12'h  c;
rom[8777] = 12'h  c;
rom[8778] = 12'h  c;
rom[8779] = 12'h  c;
rom[8780] = 12'h  c;
rom[8781] = 12'h  c;
rom[8782] = 12'h  c;
rom[8783] = 12'h  c;
rom[8784] = 12'h  c;
rom[8785] = 12'h  c;
rom[8786] = 12'h11d;
rom[8787] = 12'hddf;
rom[8788] = 12'hfff;
rom[8789] = 12'hfff;
rom[8790] = 12'hfff;
rom[8791] = 12'hfff;
rom[8792] = 12'hfff;
rom[8793] = 12'hfff;
rom[8794] = 12'hfff;
rom[8795] = 12'hfff;
rom[8796] = 12'hfff;
rom[8797] = 12'hfff;
rom[8798] = 12'hfff;
rom[8799] = 12'hfff;
rom[8800] = 12'hfff;
rom[8801] = 12'hfff;
rom[8802] = 12'hfff;
rom[8803] = 12'hfff;
rom[8804] = 12'hfff;
rom[8805] = 12'hfff;
rom[8806] = 12'hfff;
rom[8807] = 12'hfff;
rom[8808] = 12'hfff;
rom[8809] = 12'hfff;
rom[8810] = 12'hfff;
rom[8811] = 12'hfff;
rom[8812] = 12'hfff;
rom[8813] = 12'hfff;
rom[8814] = 12'hfff;
rom[8815] = 12'hfff;
rom[8816] = 12'hfff;
rom[8817] = 12'hfff;
rom[8818] = 12'hfff;
rom[8819] = 12'hfff;
rom[8820] = 12'hfff;
rom[8821] = 12'hfff;
rom[8822] = 12'hfff;
rom[8823] = 12'hfff;
rom[8824] = 12'hfff;
rom[8825] = 12'hfff;
rom[8826] = 12'hfff;
rom[8827] = 12'heef;
rom[8828] = 12'h33d;
rom[8829] = 12'h  c;
rom[8830] = 12'h  c;
rom[8831] = 12'h  c;
rom[8832] = 12'hfff;
rom[8833] = 12'hfff;
rom[8834] = 12'hfff;
rom[8835] = 12'hfff;
rom[8836] = 12'hfff;
rom[8837] = 12'hfff;
rom[8838] = 12'hfff;
rom[8839] = 12'hfff;
rom[8840] = 12'hfff;
rom[8841] = 12'hfff;
rom[8842] = 12'hfff;
rom[8843] = 12'hfff;
rom[8844] = 12'hfff;
rom[8845] = 12'hfff;
rom[8846] = 12'hfff;
rom[8847] = 12'hfff;
rom[8848] = 12'hfff;
rom[8849] = 12'hfff;
rom[8850] = 12'hfff;
rom[8851] = 12'hfff;
rom[8852] = 12'hfff;
rom[8853] = 12'hfff;
rom[8854] = 12'hfff;
rom[8855] = 12'hfff;
rom[8856] = 12'hfff;
rom[8857] = 12'hfff;
rom[8858] = 12'hfff;
rom[8859] = 12'hfff;
rom[8860] = 12'hfff;
rom[8861] = 12'hfff;
rom[8862] = 12'hfff;
rom[8863] = 12'hfff;
rom[8864] = 12'hfff;
rom[8865] = 12'hfff;
rom[8866] = 12'hfff;
rom[8867] = 12'hfff;
rom[8868] = 12'hfff;
rom[8869] = 12'hfff;
rom[8870] = 12'hfff;
rom[8871] = 12'hfff;
rom[8872] = 12'hfff;
rom[8873] = 12'hfff;
rom[8874] = 12'hfff;
rom[8875] = 12'hfff;
rom[8876] = 12'hfff;
rom[8877] = 12'hfff;
rom[8878] = 12'hfff;
rom[8879] = 12'hfff;
rom[8880] = 12'hfff;
rom[8881] = 12'hfff;
rom[8882] = 12'hfff;
rom[8883] = 12'hfff;
rom[8884] = 12'hfff;
rom[8885] = 12'hfff;
rom[8886] = 12'hfff;
rom[8887] = 12'hfff;
rom[8888] = 12'hfff;
rom[8889] = 12'hfff;
rom[8890] = 12'hfff;
rom[8891] = 12'hfff;
rom[8892] = 12'hfff;
rom[8893] = 12'hfff;
rom[8894] = 12'hfff;
rom[8895] = 12'hfff;
rom[8896] = 12'hfff;
rom[8897] = 12'hfff;
rom[8898] = 12'hfff;
rom[8899] = 12'hfff;
rom[8900] = 12'hfff;
rom[8901] = 12'hfff;
rom[8902] = 12'heef;
rom[8903] = 12'h11d;
rom[8904] = 12'h  c;
rom[8905] = 12'h  c;
rom[8906] = 12'h  c;
rom[8907] = 12'h  c;
rom[8908] = 12'h  c;
rom[8909] = 12'h  c;
rom[8910] = 12'h  c;
rom[8911] = 12'h  c;
rom[8912] = 12'h  c;
rom[8913] = 12'h  c;
rom[8914] = 12'h  c;
rom[8915] = 12'h11d;
rom[8916] = 12'h55d;
rom[8917] = 12'haae;
rom[8918] = 12'heef;
rom[8919] = 12'hfff;
rom[8920] = 12'hfff;
rom[8921] = 12'hfff;
rom[8922] = 12'hfff;
rom[8923] = 12'hfff;
rom[8924] = 12'hfff;
rom[8925] = 12'hfff;
rom[8926] = 12'hfff;
rom[8927] = 12'hfff;
rom[8928] = 12'hfff;
rom[8929] = 12'hfff;
rom[8930] = 12'hfff;
rom[8931] = 12'hfff;
rom[8932] = 12'hfff;
rom[8933] = 12'hfff;
rom[8934] = 12'hfff;
rom[8935] = 12'hfff;
rom[8936] = 12'hfff;
rom[8937] = 12'hfff;
rom[8938] = 12'hfff;
rom[8939] = 12'hfff;
rom[8940] = 12'hfff;
rom[8941] = 12'hfff;
rom[8942] = 12'hfff;
rom[8943] = 12'hfff;
rom[8944] = 12'hfff;
rom[8945] = 12'hfff;
rom[8946] = 12'hfff;
rom[8947] = 12'hfff;
rom[8948] = 12'hfff;
rom[8949] = 12'hfff;
rom[8950] = 12'hfff;
rom[8951] = 12'hfff;
rom[8952] = 12'hfff;
rom[8953] = 12'hfff;
rom[8954] = 12'heef;
rom[8955] = 12'h33d;
rom[8956] = 12'h  c;
rom[8957] = 12'h  c;
rom[8958] = 12'h  c;
rom[8959] = 12'h  c;
rom[8960] = 12'hfff;
rom[8961] = 12'hfff;
rom[8962] = 12'hfff;
rom[8963] = 12'hfff;
rom[8964] = 12'hfff;
rom[8965] = 12'hfff;
rom[8966] = 12'hfff;
rom[8967] = 12'hfff;
rom[8968] = 12'hfff;
rom[8969] = 12'hfff;
rom[8970] = 12'hfff;
rom[8971] = 12'hfff;
rom[8972] = 12'hfff;
rom[8973] = 12'hfff;
rom[8974] = 12'hfff;
rom[8975] = 12'hfff;
rom[8976] = 12'hfff;
rom[8977] = 12'hfff;
rom[8978] = 12'hfff;
rom[8979] = 12'hfff;
rom[8980] = 12'hfff;
rom[8981] = 12'hfff;
rom[8982] = 12'hfff;
rom[8983] = 12'hfff;
rom[8984] = 12'hfff;
rom[8985] = 12'hfff;
rom[8986] = 12'hfff;
rom[8987] = 12'hfff;
rom[8988] = 12'hfff;
rom[8989] = 12'hfff;
rom[8990] = 12'hfff;
rom[8991] = 12'hfff;
rom[8992] = 12'hfff;
rom[8993] = 12'hfff;
rom[8994] = 12'hfff;
rom[8995] = 12'hfff;
rom[8996] = 12'hfff;
rom[8997] = 12'hfff;
rom[8998] = 12'hfff;
rom[8999] = 12'hfff;
rom[9000] = 12'hfff;
rom[9001] = 12'hfff;
rom[9002] = 12'hfff;
rom[9003] = 12'hfff;
rom[9004] = 12'hfff;
rom[9005] = 12'hfff;
rom[9006] = 12'hfff;
rom[9007] = 12'hfff;
rom[9008] = 12'hfff;
rom[9009] = 12'hfff;
rom[9010] = 12'hfff;
rom[9011] = 12'hfff;
rom[9012] = 12'hfff;
rom[9013] = 12'hfff;
rom[9014] = 12'hfff;
rom[9015] = 12'hfff;
rom[9016] = 12'hfff;
rom[9017] = 12'hfff;
rom[9018] = 12'hfff;
rom[9019] = 12'hfff;
rom[9020] = 12'hfff;
rom[9021] = 12'hfff;
rom[9022] = 12'hfff;
rom[9023] = 12'hfff;
rom[9024] = 12'hfff;
rom[9025] = 12'hfff;
rom[9026] = 12'hfff;
rom[9027] = 12'hfff;
rom[9028] = 12'hfff;
rom[9029] = 12'hfff;
rom[9030] = 12'hfff;
rom[9031] = 12'hbbf;
rom[9032] = 12'h  c;
rom[9033] = 12'h  c;
rom[9034] = 12'h  c;
rom[9035] = 12'h  c;
rom[9036] = 12'h  c;
rom[9037] = 12'h  c;
rom[9038] = 12'h  c;
rom[9039] = 12'h  c;
rom[9040] = 12'h  c;
rom[9041] = 12'h  c;
rom[9042] = 12'h  c;
rom[9043] = 12'h  c;
rom[9044] = 12'h  c;
rom[9045] = 12'h  c;
rom[9046] = 12'h11d;
rom[9047] = 12'heef;
rom[9048] = 12'hfff;
rom[9049] = 12'hfff;
rom[9050] = 12'hfff;
rom[9051] = 12'hfff;
rom[9052] = 12'hfff;
rom[9053] = 12'hfff;
rom[9054] = 12'hfff;
rom[9055] = 12'hfff;
rom[9056] = 12'hfff;
rom[9057] = 12'hfff;
rom[9058] = 12'hfff;
rom[9059] = 12'hfff;
rom[9060] = 12'hfff;
rom[9061] = 12'hfff;
rom[9062] = 12'hfff;
rom[9063] = 12'hfff;
rom[9064] = 12'hfff;
rom[9065] = 12'hfff;
rom[9066] = 12'hfff;
rom[9067] = 12'hfff;
rom[9068] = 12'hfff;
rom[9069] = 12'hfff;
rom[9070] = 12'hfff;
rom[9071] = 12'hfff;
rom[9072] = 12'hfff;
rom[9073] = 12'hfff;
rom[9074] = 12'hfff;
rom[9075] = 12'hfff;
rom[9076] = 12'hfff;
rom[9077] = 12'hfff;
rom[9078] = 12'hfff;
rom[9079] = 12'hfff;
rom[9080] = 12'hfff;
rom[9081] = 12'h99e;
rom[9082] = 12'h11d;
rom[9083] = 12'h  c;
rom[9084] = 12'h  c;
rom[9085] = 12'h  c;
rom[9086] = 12'h  c;
rom[9087] = 12'h  c;
rom[9088] = 12'hfff;
rom[9089] = 12'hfff;
rom[9090] = 12'hfff;
rom[9091] = 12'hfff;
rom[9092] = 12'hfff;
rom[9093] = 12'hfff;
rom[9094] = 12'hfff;
rom[9095] = 12'hfff;
rom[9096] = 12'hfff;
rom[9097] = 12'hfff;
rom[9098] = 12'hfff;
rom[9099] = 12'hfff;
rom[9100] = 12'hfff;
rom[9101] = 12'hfff;
rom[9102] = 12'hfff;
rom[9103] = 12'hfff;
rom[9104] = 12'hfff;
rom[9105] = 12'hfff;
rom[9106] = 12'hfff;
rom[9107] = 12'hfff;
rom[9108] = 12'hfff;
rom[9109] = 12'hfff;
rom[9110] = 12'hfff;
rom[9111] = 12'hfff;
rom[9112] = 12'hfff;
rom[9113] = 12'hfff;
rom[9114] = 12'hfff;
rom[9115] = 12'hfff;
rom[9116] = 12'hfff;
rom[9117] = 12'hfff;
rom[9118] = 12'hfff;
rom[9119] = 12'hfff;
rom[9120] = 12'hfff;
rom[9121] = 12'hfff;
rom[9122] = 12'hfff;
rom[9123] = 12'hfff;
rom[9124] = 12'hfff;
rom[9125] = 12'hfff;
rom[9126] = 12'hfff;
rom[9127] = 12'hfff;
rom[9128] = 12'hfff;
rom[9129] = 12'hfff;
rom[9130] = 12'hfff;
rom[9131] = 12'hfff;
rom[9132] = 12'heef;
rom[9133] = 12'h99e;
rom[9134] = 12'h77e;
rom[9135] = 12'h66e;
rom[9136] = 12'h55d;
rom[9137] = 12'h44d;
rom[9138] = 12'h33d;
rom[9139] = 12'h33d;
rom[9140] = 12'h33d;
rom[9141] = 12'h33d;
rom[9142] = 12'h33d;
rom[9143] = 12'h33d;
rom[9144] = 12'h44d;
rom[9145] = 12'h88e;
rom[9146] = 12'heef;
rom[9147] = 12'hfff;
rom[9148] = 12'hfff;
rom[9149] = 12'hfff;
rom[9150] = 12'hfff;
rom[9151] = 12'hfff;
rom[9152] = 12'hfff;
rom[9153] = 12'hfff;
rom[9154] = 12'hfff;
rom[9155] = 12'hfff;
rom[9156] = 12'hfff;
rom[9157] = 12'hfff;
rom[9158] = 12'hfff;
rom[9159] = 12'hfff;
rom[9160] = 12'haae;
rom[9161] = 12'h  c;
rom[9162] = 12'h  c;
rom[9163] = 12'h  c;
rom[9164] = 12'h  c;
rom[9165] = 12'h  c;
rom[9166] = 12'h  c;
rom[9167] = 12'h  c;
rom[9168] = 12'h  c;
rom[9169] = 12'h  c;
rom[9170] = 12'h  c;
rom[9171] = 12'h  c;
rom[9172] = 12'h  c;
rom[9173] = 12'h  c;
rom[9174] = 12'h  c;
rom[9175] = 12'h88e;
rom[9176] = 12'hfff;
rom[9177] = 12'hfff;
rom[9178] = 12'hfff;
rom[9179] = 12'hfff;
rom[9180] = 12'hfff;
rom[9181] = 12'hfff;
rom[9182] = 12'hfff;
rom[9183] = 12'hfff;
rom[9184] = 12'hfff;
rom[9185] = 12'hfff;
rom[9186] = 12'hfff;
rom[9187] = 12'hfff;
rom[9188] = 12'hfff;
rom[9189] = 12'hfff;
rom[9190] = 12'hfff;
rom[9191] = 12'hfff;
rom[9192] = 12'hfff;
rom[9193] = 12'hfff;
rom[9194] = 12'hfff;
rom[9195] = 12'hfff;
rom[9196] = 12'hfff;
rom[9197] = 12'hfff;
rom[9198] = 12'hfff;
rom[9199] = 12'hfff;
rom[9200] = 12'hfff;
rom[9201] = 12'hfff;
rom[9202] = 12'hfff;
rom[9203] = 12'hfff;
rom[9204] = 12'hfff;
rom[9205] = 12'hfff;
rom[9206] = 12'hfff;
rom[9207] = 12'heef;
rom[9208] = 12'h44d;
rom[9209] = 12'h  c;
rom[9210] = 12'h  c;
rom[9211] = 12'h  c;
rom[9212] = 12'h  c;
rom[9213] = 12'h  c;
rom[9214] = 12'h  c;
rom[9215] = 12'h  c;
rom[9216] = 12'hfff;
rom[9217] = 12'hfff;
rom[9218] = 12'hfff;
rom[9219] = 12'hfff;
rom[9220] = 12'hfff;
rom[9221] = 12'hfff;
rom[9222] = 12'hfff;
rom[9223] = 12'hfff;
rom[9224] = 12'hfff;
rom[9225] = 12'hfff;
rom[9226] = 12'hfff;
rom[9227] = 12'hfff;
rom[9228] = 12'hfff;
rom[9229] = 12'hfff;
rom[9230] = 12'hfff;
rom[9231] = 12'hfff;
rom[9232] = 12'hfff;
rom[9233] = 12'hfff;
rom[9234] = 12'hfff;
rom[9235] = 12'hfff;
rom[9236] = 12'hfff;
rom[9237] = 12'hfff;
rom[9238] = 12'hfff;
rom[9239] = 12'hfff;
rom[9240] = 12'hfff;
rom[9241] = 12'hfff;
rom[9242] = 12'hfff;
rom[9243] = 12'hfff;
rom[9244] = 12'hfff;
rom[9245] = 12'hfff;
rom[9246] = 12'hfff;
rom[9247] = 12'hfff;
rom[9248] = 12'hfff;
rom[9249] = 12'hfff;
rom[9250] = 12'hfff;
rom[9251] = 12'hfff;
rom[9252] = 12'hfff;
rom[9253] = 12'hfff;
rom[9254] = 12'hfff;
rom[9255] = 12'hfff;
rom[9256] = 12'hfff;
rom[9257] = 12'hfff;
rom[9258] = 12'hfff;
rom[9259] = 12'heef;
rom[9260] = 12'h11d;
rom[9261] = 12'h  c;
rom[9262] = 12'h  c;
rom[9263] = 12'h  c;
rom[9264] = 12'h  c;
rom[9265] = 12'h  c;
rom[9266] = 12'h  c;
rom[9267] = 12'h  c;
rom[9268] = 12'h  c;
rom[9269] = 12'h  c;
rom[9270] = 12'h  c;
rom[9271] = 12'h  c;
rom[9272] = 12'h  c;
rom[9273] = 12'h  c;
rom[9274] = 12'h11d;
rom[9275] = 12'hbbf;
rom[9276] = 12'hfff;
rom[9277] = 12'hfff;
rom[9278] = 12'hfff;
rom[9279] = 12'hfff;
rom[9280] = 12'hfff;
rom[9281] = 12'hfff;
rom[9282] = 12'hfff;
rom[9283] = 12'hfff;
rom[9284] = 12'hfff;
rom[9285] = 12'hfff;
rom[9286] = 12'hfff;
rom[9287] = 12'hfff;
rom[9288] = 12'hfff;
rom[9289] = 12'hbbf;
rom[9290] = 12'h11d;
rom[9291] = 12'h  c;
rom[9292] = 12'h  c;
rom[9293] = 12'h  c;
rom[9294] = 12'h  c;
rom[9295] = 12'h  c;
rom[9296] = 12'h  c;
rom[9297] = 12'h  c;
rom[9298] = 12'h  c;
rom[9299] = 12'h  c;
rom[9300] = 12'h  c;
rom[9301] = 12'h  c;
rom[9302] = 12'h  c;
rom[9303] = 12'h  c;
rom[9304] = 12'h55d;
rom[9305] = 12'h77e;
rom[9306] = 12'haae;
rom[9307] = 12'hccf;
rom[9308] = 12'heef;
rom[9309] = 12'hfff;
rom[9310] = 12'hfff;
rom[9311] = 12'hfff;
rom[9312] = 12'hfff;
rom[9313] = 12'hfff;
rom[9314] = 12'hfff;
rom[9315] = 12'hfff;
rom[9316] = 12'hfff;
rom[9317] = 12'hfff;
rom[9318] = 12'hfff;
rom[9319] = 12'hfff;
rom[9320] = 12'hfff;
rom[9321] = 12'hfff;
rom[9322] = 12'hfff;
rom[9323] = 12'hfff;
rom[9324] = 12'hfff;
rom[9325] = 12'hfff;
rom[9326] = 12'hfff;
rom[9327] = 12'hfff;
rom[9328] = 12'hfff;
rom[9329] = 12'hfff;
rom[9330] = 12'heef;
rom[9331] = 12'hccf;
rom[9332] = 12'haae;
rom[9333] = 12'h77e;
rom[9334] = 12'h55d;
rom[9335] = 12'h11c;
rom[9336] = 12'h  c;
rom[9337] = 12'h  c;
rom[9338] = 12'h  c;
rom[9339] = 12'h  c;
rom[9340] = 12'h  c;
rom[9341] = 12'h  c;
rom[9342] = 12'h11d;
rom[9343] = 12'hccf;
rom[9344] = 12'hfff;
rom[9345] = 12'hfff;
rom[9346] = 12'hfff;
rom[9347] = 12'hfff;
rom[9348] = 12'hfff;
rom[9349] = 12'hfff;
rom[9350] = 12'hfff;
rom[9351] = 12'hfff;
rom[9352] = 12'hfff;
rom[9353] = 12'hfff;
rom[9354] = 12'hfff;
rom[9355] = 12'hfff;
rom[9356] = 12'hfff;
rom[9357] = 12'hfff;
rom[9358] = 12'hfff;
rom[9359] = 12'hfff;
rom[9360] = 12'hfff;
rom[9361] = 12'hfff;
rom[9362] = 12'hfff;
rom[9363] = 12'hfff;
rom[9364] = 12'hfff;
rom[9365] = 12'hfff;
rom[9366] = 12'hfff;
rom[9367] = 12'hfff;
rom[9368] = 12'hfff;
rom[9369] = 12'hfff;
rom[9370] = 12'hfff;
rom[9371] = 12'hfff;
rom[9372] = 12'hfff;
rom[9373] = 12'hfff;
rom[9374] = 12'hfff;
rom[9375] = 12'hfff;
rom[9376] = 12'hfff;
rom[9377] = 12'hfff;
rom[9378] = 12'hfff;
rom[9379] = 12'hfff;
rom[9380] = 12'hfff;
rom[9381] = 12'hfff;
rom[9382] = 12'hfff;
rom[9383] = 12'hfff;
rom[9384] = 12'hfff;
rom[9385] = 12'hfff;
rom[9386] = 12'hfff;
rom[9387] = 12'h99e;
rom[9388] = 12'h  c;
rom[9389] = 12'h  c;
rom[9390] = 12'h  c;
rom[9391] = 12'h  c;
rom[9392] = 12'h  c;
rom[9393] = 12'h  c;
rom[9394] = 12'h  c;
rom[9395] = 12'h  c;
rom[9396] = 12'h  c;
rom[9397] = 12'h  c;
rom[9398] = 12'h  c;
rom[9399] = 12'h  c;
rom[9400] = 12'h  c;
rom[9401] = 12'h  c;
rom[9402] = 12'h  c;
rom[9403] = 12'h  c;
rom[9404] = 12'haae;
rom[9405] = 12'hfff;
rom[9406] = 12'hfff;
rom[9407] = 12'hfff;
rom[9408] = 12'hfff;
rom[9409] = 12'hfff;
rom[9410] = 12'hfff;
rom[9411] = 12'hfff;
rom[9412] = 12'hfff;
rom[9413] = 12'hfff;
rom[9414] = 12'hfff;
rom[9415] = 12'hfff;
rom[9416] = 12'hfff;
rom[9417] = 12'hfff;
rom[9418] = 12'heef;
rom[9419] = 12'h99e;
rom[9420] = 12'h77e;
rom[9421] = 12'h77e;
rom[9422] = 12'h88e;
rom[9423] = 12'h55d;
rom[9424] = 12'h11d;
rom[9425] = 12'h  c;
rom[9426] = 12'h  c;
rom[9427] = 12'h  c;
rom[9428] = 12'h  c;
rom[9429] = 12'h  c;
rom[9430] = 12'h  c;
rom[9431] = 12'h  c;
rom[9432] = 12'h  c;
rom[9433] = 12'h  c;
rom[9434] = 12'h  c;
rom[9435] = 12'h  c;
rom[9436] = 12'h  c;
rom[9437] = 12'h  c;
rom[9438] = 12'h  c;
rom[9439] = 12'h11d;
rom[9440] = 12'h22d;
rom[9441] = 12'h33d;
rom[9442] = 12'h44d;
rom[9443] = 12'h44d;
rom[9444] = 12'h44d;
rom[9445] = 12'h55d;
rom[9446] = 12'h55d;
rom[9447] = 12'h55d;
rom[9448] = 12'h55d;
rom[9449] = 12'h55d;
rom[9450] = 12'h44d;
rom[9451] = 12'h44d;
rom[9452] = 12'h44d;
rom[9453] = 12'h33d;
rom[9454] = 12'h22d;
rom[9455] = 12'h11d;
rom[9456] = 12'h  c;
rom[9457] = 12'h  c;
rom[9458] = 12'h  c;
rom[9459] = 12'h  c;
rom[9460] = 12'h  c;
rom[9461] = 12'h  c;
rom[9462] = 12'h  c;
rom[9463] = 12'h  c;
rom[9464] = 12'h  c;
rom[9465] = 12'h  c;
rom[9466] = 12'h  c;
rom[9467] = 12'h  c;
rom[9468] = 12'h  c;
rom[9469] = 12'h22d;
rom[9470] = 12'hddf;
rom[9471] = 12'hfff;
rom[9472] = 12'hfff;
rom[9473] = 12'hfff;
rom[9474] = 12'hfff;
rom[9475] = 12'hfff;
rom[9476] = 12'hfff;
rom[9477] = 12'hfff;
rom[9478] = 12'hfff;
rom[9479] = 12'hfff;
rom[9480] = 12'hfff;
rom[9481] = 12'hfff;
rom[9482] = 12'hfff;
rom[9483] = 12'hfff;
rom[9484] = 12'hfff;
rom[9485] = 12'hfff;
rom[9486] = 12'hfff;
rom[9487] = 12'hfff;
rom[9488] = 12'hfff;
rom[9489] = 12'hfff;
rom[9490] = 12'hfff;
rom[9491] = 12'hfff;
rom[9492] = 12'hfff;
rom[9493] = 12'hfff;
rom[9494] = 12'hfff;
rom[9495] = 12'hfff;
rom[9496] = 12'hfff;
rom[9497] = 12'hfff;
rom[9498] = 12'hfff;
rom[9499] = 12'hfff;
rom[9500] = 12'hfff;
rom[9501] = 12'hfff;
rom[9502] = 12'h99e;
rom[9503] = 12'h55d;
rom[9504] = 12'h33d;
rom[9505] = 12'h22d;
rom[9506] = 12'h22d;
rom[9507] = 12'h11d;
rom[9508] = 12'h11c;
rom[9509] = 12'h11c;
rom[9510] = 12'h11c;
rom[9511] = 12'h11c;
rom[9512] = 12'h11d;
rom[9513] = 12'h22d;
rom[9514] = 12'h22d;
rom[9515] = 12'h11d;
rom[9516] = 12'h  c;
rom[9517] = 12'h  c;
rom[9518] = 12'h  c;
rom[9519] = 12'h  c;
rom[9520] = 12'h  c;
rom[9521] = 12'h  c;
rom[9522] = 12'h  c;
rom[9523] = 12'h  c;
rom[9524] = 12'h  c;
rom[9525] = 12'h  c;
rom[9526] = 12'h  c;
rom[9527] = 12'h  c;
rom[9528] = 12'h  c;
rom[9529] = 12'h  c;
rom[9530] = 12'h  c;
rom[9531] = 12'h  c;
rom[9532] = 12'h  c;
rom[9533] = 12'hbbf;
rom[9534] = 12'hfff;
rom[9535] = 12'hfff;
rom[9536] = 12'hfff;
rom[9537] = 12'hfff;
rom[9538] = 12'hfff;
rom[9539] = 12'hfff;
rom[9540] = 12'hfff;
rom[9541] = 12'hfff;
rom[9542] = 12'hfff;
rom[9543] = 12'hfff;
rom[9544] = 12'hfff;
rom[9545] = 12'hfff;
rom[9546] = 12'hfff;
rom[9547] = 12'hfff;
rom[9548] = 12'hfff;
rom[9549] = 12'hfff;
rom[9550] = 12'hfff;
rom[9551] = 12'hfff;
rom[9552] = 12'hddf;
rom[9553] = 12'h44d;
rom[9554] = 12'h  c;
rom[9555] = 12'h  c;
rom[9556] = 12'h  c;
rom[9557] = 12'h  c;
rom[9558] = 12'h  c;
rom[9559] = 12'h  c;
rom[9560] = 12'h  c;
rom[9561] = 12'h  c;
rom[9562] = 12'h  c;
rom[9563] = 12'h  c;
rom[9564] = 12'h  c;
rom[9565] = 12'h  c;
rom[9566] = 12'h  c;
rom[9567] = 12'h  c;
rom[9568] = 12'h  c;
rom[9569] = 12'h  c;
rom[9570] = 12'h  c;
rom[9571] = 12'h  c;
rom[9572] = 12'h  c;
rom[9573] = 12'h  c;
rom[9574] = 12'h  c;
rom[9575] = 12'h  c;
rom[9576] = 12'h  c;
rom[9577] = 12'h  c;
rom[9578] = 12'h  c;
rom[9579] = 12'h  c;
rom[9580] = 12'h  c;
rom[9581] = 12'h  c;
rom[9582] = 12'h  c;
rom[9583] = 12'h  c;
rom[9584] = 12'h  c;
rom[9585] = 12'h  c;
rom[9586] = 12'h  c;
rom[9587] = 12'h  c;
rom[9588] = 12'h  c;
rom[9589] = 12'h  c;
rom[9590] = 12'h  c;
rom[9591] = 12'h  c;
rom[9592] = 12'h  c;
rom[9593] = 12'h  c;
rom[9594] = 12'h  c;
rom[9595] = 12'h11d;
rom[9596] = 12'h99e;
rom[9597] = 12'hfff;
rom[9598] = 12'hfff;
rom[9599] = 12'hfff;
rom[9600] = 12'hfff;
rom[9601] = 12'hfff;
rom[9602] = 12'hfff;
rom[9603] = 12'hfff;
rom[9604] = 12'hfff;
rom[9605] = 12'hfff;
rom[9606] = 12'hfff;
rom[9607] = 12'hfff;
rom[9608] = 12'hfff;
rom[9609] = 12'hfff;
rom[9610] = 12'hfff;
rom[9611] = 12'hfff;
rom[9612] = 12'hfff;
rom[9613] = 12'hfff;
rom[9614] = 12'hfff;
rom[9615] = 12'hfff;
rom[9616] = 12'hfff;
rom[9617] = 12'hfff;
rom[9618] = 12'hfff;
rom[9619] = 12'hfff;
rom[9620] = 12'hfff;
rom[9621] = 12'hfff;
rom[9622] = 12'hfff;
rom[9623] = 12'hfff;
rom[9624] = 12'hfff;
rom[9625] = 12'hfff;
rom[9626] = 12'hfff;
rom[9627] = 12'haae;
rom[9628] = 12'h99e;
rom[9629] = 12'h33d;
rom[9630] = 12'h  c;
rom[9631] = 12'h  c;
rom[9632] = 12'h  c;
rom[9633] = 12'h  c;
rom[9634] = 12'h  c;
rom[9635] = 12'h  c;
rom[9636] = 12'h  c;
rom[9637] = 12'h  c;
rom[9638] = 12'h  c;
rom[9639] = 12'h  c;
rom[9640] = 12'h  c;
rom[9641] = 12'h  c;
rom[9642] = 12'h  c;
rom[9643] = 12'h  c;
rom[9644] = 12'h  c;
rom[9645] = 12'h  c;
rom[9646] = 12'h  c;
rom[9647] = 12'h  c;
rom[9648] = 12'h  c;
rom[9649] = 12'h  c;
rom[9650] = 12'h  c;
rom[9651] = 12'h  c;
rom[9652] = 12'h  c;
rom[9653] = 12'h  c;
rom[9654] = 12'h  c;
rom[9655] = 12'h  c;
rom[9656] = 12'h  c;
rom[9657] = 12'h  c;
rom[9658] = 12'h  c;
rom[9659] = 12'h  c;
rom[9660] = 12'h  c;
rom[9661] = 12'h11d;
rom[9662] = 12'heef;
rom[9663] = 12'hfff;
rom[9664] = 12'hfff;
rom[9665] = 12'hfff;
rom[9666] = 12'hfff;
rom[9667] = 12'hfff;
rom[9668] = 12'hfff;
rom[9669] = 12'hfff;
rom[9670] = 12'hfff;
rom[9671] = 12'hfff;
rom[9672] = 12'hfff;
rom[9673] = 12'hfff;
rom[9674] = 12'hfff;
rom[9675] = 12'hfff;
rom[9676] = 12'hfff;
rom[9677] = 12'hfff;
rom[9678] = 12'hfff;
rom[9679] = 12'hfff;
rom[9680] = 12'hfff;
rom[9681] = 12'heef;
rom[9682] = 12'h99e;
rom[9683] = 12'h66e;
rom[9684] = 12'h  c;
rom[9685] = 12'h  c;
rom[9686] = 12'h  c;
rom[9687] = 12'h  c;
rom[9688] = 12'h  c;
rom[9689] = 12'h  c;
rom[9690] = 12'h  c;
rom[9691] = 12'h  c;
rom[9692] = 12'h  c;
rom[9693] = 12'h  c;
rom[9694] = 12'h  c;
rom[9695] = 12'h  c;
rom[9696] = 12'h  c;
rom[9697] = 12'h  c;
rom[9698] = 12'h  c;
rom[9699] = 12'h  c;
rom[9700] = 12'h  c;
rom[9701] = 12'h  c;
rom[9702] = 12'h  c;
rom[9703] = 12'h  c;
rom[9704] = 12'h  c;
rom[9705] = 12'h  c;
rom[9706] = 12'h  c;
rom[9707] = 12'h  c;
rom[9708] = 12'h  c;
rom[9709] = 12'h  c;
rom[9710] = 12'h  c;
rom[9711] = 12'h  c;
rom[9712] = 12'h  c;
rom[9713] = 12'h  c;
rom[9714] = 12'h  c;
rom[9715] = 12'h  c;
rom[9716] = 12'h  c;
rom[9717] = 12'h  c;
rom[9718] = 12'h  c;
rom[9719] = 12'h  c;
rom[9720] = 12'h  c;
rom[9721] = 12'h  c;
rom[9722] = 12'h33d;
rom[9723] = 12'heef;
rom[9724] = 12'hfff;
rom[9725] = 12'hfff;
rom[9726] = 12'hfff;
rom[9727] = 12'hfff;
rom[9728] = 12'hfff;
rom[9729] = 12'hfff;
rom[9730] = 12'hfff;
rom[9731] = 12'hfff;
rom[9732] = 12'hfff;
rom[9733] = 12'hfff;
rom[9734] = 12'hfff;
rom[9735] = 12'hfff;
rom[9736] = 12'hfff;
rom[9737] = 12'hfff;
rom[9738] = 12'hfff;
rom[9739] = 12'hfff;
rom[9740] = 12'hfff;
rom[9741] = 12'hfff;
rom[9742] = 12'hfff;
rom[9743] = 12'hfff;
rom[9744] = 12'hfff;
rom[9745] = 12'hfff;
rom[9746] = 12'hfff;
rom[9747] = 12'hfff;
rom[9748] = 12'hfff;
rom[9749] = 12'hfff;
rom[9750] = 12'hfff;
rom[9751] = 12'hfff;
rom[9752] = 12'hbbf;
rom[9753] = 12'h55d;
rom[9754] = 12'h  c;
rom[9755] = 12'h  c;
rom[9756] = 12'h  c;
rom[9757] = 12'h  c;
rom[9758] = 12'h  c;
rom[9759] = 12'h  c;
rom[9760] = 12'h  c;
rom[9761] = 12'h  c;
rom[9762] = 12'h  c;
rom[9763] = 12'h  c;
rom[9764] = 12'h  c;
rom[9765] = 12'h  c;
rom[9766] = 12'h  c;
rom[9767] = 12'h  c;
rom[9768] = 12'h  c;
rom[9769] = 12'h  c;
rom[9770] = 12'h  c;
rom[9771] = 12'h  c;
rom[9772] = 12'h  c;
rom[9773] = 12'h  c;
rom[9774] = 12'h  c;
rom[9775] = 12'h  c;
rom[9776] = 12'h  c;
rom[9777] = 12'h  c;
rom[9778] = 12'h44d;
rom[9779] = 12'hbbf;
rom[9780] = 12'hccf;
rom[9781] = 12'hccf;
rom[9782] = 12'hccf;
rom[9783] = 12'hccf;
rom[9784] = 12'h44d;
rom[9785] = 12'h  c;
rom[9786] = 12'h  c;
rom[9787] = 12'h  c;
rom[9788] = 12'h  c;
rom[9789] = 12'h  c;
rom[9790] = 12'h77e;
rom[9791] = 12'hfff;
rom[9792] = 12'hfff;
rom[9793] = 12'hfff;
rom[9794] = 12'hfff;
rom[9795] = 12'hfff;
rom[9796] = 12'hfff;
rom[9797] = 12'hfff;
rom[9798] = 12'hfff;
rom[9799] = 12'hfff;
rom[9800] = 12'hfff;
rom[9801] = 12'hfff;
rom[9802] = 12'hfff;
rom[9803] = 12'hfff;
rom[9804] = 12'hfff;
rom[9805] = 12'hfff;
rom[9806] = 12'hfff;
rom[9807] = 12'hfff;
rom[9808] = 12'hfff;
rom[9809] = 12'hfff;
rom[9810] = 12'hfff;
rom[9811] = 12'hfff;
rom[9812] = 12'haae;
rom[9813] = 12'h  c;
rom[9814] = 12'h  c;
rom[9815] = 12'h  c;
rom[9816] = 12'h  c;
rom[9817] = 12'h  c;
rom[9818] = 12'h  c;
rom[9819] = 12'h  c;
rom[9820] = 12'h  c;
rom[9821] = 12'h  c;
rom[9822] = 12'h  c;
rom[9823] = 12'h  c;
rom[9824] = 12'h  c;
rom[9825] = 12'h  c;
rom[9826] = 12'h  c;
rom[9827] = 12'h  c;
rom[9828] = 12'h  c;
rom[9829] = 12'h  c;
rom[9830] = 12'h  c;
rom[9831] = 12'h  c;
rom[9832] = 12'h  c;
rom[9833] = 12'h  c;
rom[9834] = 12'h  c;
rom[9835] = 12'h  c;
rom[9836] = 12'h  c;
rom[9837] = 12'h  c;
rom[9838] = 12'h  c;
rom[9839] = 12'h  c;
rom[9840] = 12'h  c;
rom[9841] = 12'h  c;
rom[9842] = 12'h  c;
rom[9843] = 12'h  c;
rom[9844] = 12'h  c;
rom[9845] = 12'h  c;
rom[9846] = 12'h  c;
rom[9847] = 12'h  c;
rom[9848] = 12'h11d;
rom[9849] = 12'h77e;
rom[9850] = 12'hfff;
rom[9851] = 12'hfff;
rom[9852] = 12'hfff;
rom[9853] = 12'hfff;
rom[9854] = 12'hfff;
rom[9855] = 12'hfff;
rom[9856] = 12'hfff;
rom[9857] = 12'hfff;
rom[9858] = 12'hfff;
rom[9859] = 12'hfff;
rom[9860] = 12'hfff;
rom[9861] = 12'hfff;
rom[9862] = 12'hfff;
rom[9863] = 12'hfff;
rom[9864] = 12'hfff;
rom[9865] = 12'hfff;
rom[9866] = 12'hfff;
rom[9867] = 12'hfff;
rom[9868] = 12'hfff;
rom[9869] = 12'hfff;
rom[9870] = 12'hfff;
rom[9871] = 12'hfff;
rom[9872] = 12'hfff;
rom[9873] = 12'hfff;
rom[9874] = 12'hfff;
rom[9875] = 12'hfff;
rom[9876] = 12'hfff;
rom[9877] = 12'hfff;
rom[9878] = 12'heef;
rom[9879] = 12'h33d;
rom[9880] = 12'h  c;
rom[9881] = 12'h  c;
rom[9882] = 12'h  c;
rom[9883] = 12'h  c;
rom[9884] = 12'h  c;
rom[9885] = 12'h  c;
rom[9886] = 12'h  c;
rom[9887] = 12'h  c;
rom[9888] = 12'h  c;
rom[9889] = 12'h  c;
rom[9890] = 12'h  c;
rom[9891] = 12'h  c;
rom[9892] = 12'h  c;
rom[9893] = 12'h  c;
rom[9894] = 12'h  c;
rom[9895] = 12'h  c;
rom[9896] = 12'h  c;
rom[9897] = 12'h  c;
rom[9898] = 12'h  c;
rom[9899] = 12'h  c;
rom[9900] = 12'h  c;
rom[9901] = 12'h  c;
rom[9902] = 12'h  c;
rom[9903] = 12'h  c;
rom[9904] = 12'h  c;
rom[9905] = 12'h  c;
rom[9906] = 12'h  c;
rom[9907] = 12'h11d;
rom[9908] = 12'heef;
rom[9909] = 12'hfff;
rom[9910] = 12'hfff;
rom[9911] = 12'hfff;
rom[9912] = 12'hfff;
rom[9913] = 12'h55d;
rom[9914] = 12'h  c;
rom[9915] = 12'h  c;
rom[9916] = 12'h  c;
rom[9917] = 12'h  c;
rom[9918] = 12'h22d;
rom[9919] = 12'hfff;
rom[9920] = 12'hfff;
rom[9921] = 12'hfff;
rom[9922] = 12'hfff;
rom[9923] = 12'hfff;
rom[9924] = 12'hfff;
rom[9925] = 12'hfff;
rom[9926] = 12'hfff;
rom[9927] = 12'hfff;
rom[9928] = 12'hfff;
rom[9929] = 12'hfff;
rom[9930] = 12'hfff;
rom[9931] = 12'hfff;
rom[9932] = 12'hfff;
rom[9933] = 12'hfff;
rom[9934] = 12'hfff;
rom[9935] = 12'hfff;
rom[9936] = 12'hfff;
rom[9937] = 12'hfff;
rom[9938] = 12'hfff;
rom[9939] = 12'hfff;
rom[9940] = 12'hfff;
rom[9941] = 12'hbbf;
rom[9942] = 12'h11c;
rom[9943] = 12'h  c;
rom[9944] = 12'h  c;
rom[9945] = 12'h  c;
rom[9946] = 12'h  c;
rom[9947] = 12'h  c;
rom[9948] = 12'h  c;
rom[9949] = 12'h  c;
rom[9950] = 12'h  c;
rom[9951] = 12'h  c;
rom[9952] = 12'h  c;
rom[9953] = 12'h  c;
rom[9954] = 12'h  c;
rom[9955] = 12'h  c;
rom[9956] = 12'h  c;
rom[9957] = 12'h  c;
rom[9958] = 12'h  c;
rom[9959] = 12'h  c;
rom[9960] = 12'h  c;
rom[9961] = 12'h  c;
rom[9962] = 12'h  c;
rom[9963] = 12'h  c;
rom[9964] = 12'h  c;
rom[9965] = 12'h  c;
rom[9966] = 12'h  c;
rom[9967] = 12'h  c;
rom[9968] = 12'h  c;
rom[9969] = 12'h  c;
rom[9970] = 12'h11d;
rom[9971] = 12'h22d;
rom[9972] = 12'h55d;
rom[9973] = 12'h77e;
rom[9974] = 12'h99e;
rom[9975] = 12'hccf;
rom[9976] = 12'hfff;
rom[9977] = 12'hfff;
rom[9978] = 12'hfff;
rom[9979] = 12'hfff;
rom[9980] = 12'hfff;
rom[9981] = 12'hfff;
rom[9982] = 12'hfff;
rom[9983] = 12'hfff;
rom[9984] = 12'hfff;
rom[9985] = 12'hfff;
rom[9986] = 12'hfff;
rom[9987] = 12'hfff;
rom[9988] = 12'hfff;
rom[9989] = 12'hfff;
rom[9990] = 12'hfff;
rom[9991] = 12'hfff;
rom[9992] = 12'hfff;
rom[9993] = 12'hfff;
rom[9994] = 12'hfff;
rom[9995] = 12'hfff;
rom[9996] = 12'hfff;
rom[9997] = 12'hfff;
rom[9998] = 12'hfff;
rom[9999] = 12'hfff;
rom[10000] = 12'hfff;
rom[10001] = 12'hfff;
rom[10002] = 12'hfff;
rom[10003] = 12'hfff;
rom[10004] = 12'hfff;
rom[10005] = 12'hfff;
rom[10006] = 12'h44d;
rom[10007] = 12'h  c;
rom[10008] = 12'h  c;
rom[10009] = 12'h  c;
rom[10010] = 12'h  c;
rom[10011] = 12'h  c;
rom[10012] = 12'h  c;
rom[10013] = 12'h  c;
rom[10014] = 12'h  c;
rom[10015] = 12'h  c;
rom[10016] = 12'h  c;
rom[10017] = 12'h  c;
rom[10018] = 12'h  c;
rom[10019] = 12'h  c;
rom[10020] = 12'h  c;
rom[10021] = 12'h  c;
rom[10022] = 12'h  c;
rom[10023] = 12'h  c;
rom[10024] = 12'h  c;
rom[10025] = 12'h  c;
rom[10026] = 12'h  c;
rom[10027] = 12'h  c;
rom[10028] = 12'h  c;
rom[10029] = 12'h  c;
rom[10030] = 12'h  c;
rom[10031] = 12'h  c;
rom[10032] = 12'h  c;
rom[10033] = 12'h  c;
rom[10034] = 12'h  c;
rom[10035] = 12'h  c;
rom[10036] = 12'h99e;
rom[10037] = 12'hfff;
rom[10038] = 12'hfff;
rom[10039] = 12'hfff;
rom[10040] = 12'hfff;
rom[10041] = 12'heef;
rom[10042] = 12'h  c;
rom[10043] = 12'h  c;
rom[10044] = 12'h  c;
rom[10045] = 12'h  c;
rom[10046] = 12'h  c;
rom[10047] = 12'hfff;
rom[10048] = 12'hfff;
rom[10049] = 12'hfff;
rom[10050] = 12'hfff;
rom[10051] = 12'hfff;
rom[10052] = 12'hfff;
rom[10053] = 12'hfff;
rom[10054] = 12'hfff;
rom[10055] = 12'hfff;
rom[10056] = 12'hfff;
rom[10057] = 12'hfff;
rom[10058] = 12'hfff;
rom[10059] = 12'hfff;
rom[10060] = 12'hfff;
rom[10061] = 12'hfff;
rom[10062] = 12'hfff;
rom[10063] = 12'hfff;
rom[10064] = 12'hfff;
rom[10065] = 12'hfff;
rom[10066] = 12'hfff;
rom[10067] = 12'hfff;
rom[10068] = 12'hfff;
rom[10069] = 12'hfff;
rom[10070] = 12'hddf;
rom[10071] = 12'h22d;
rom[10072] = 12'h  c;
rom[10073] = 12'h  c;
rom[10074] = 12'h  c;
rom[10075] = 12'h  c;
rom[10076] = 12'h  c;
rom[10077] = 12'h88e;
rom[10078] = 12'hfff;
rom[10079] = 12'heef;
rom[10080] = 12'hddf;
rom[10081] = 12'hccf;
rom[10082] = 12'hbbf;
rom[10083] = 12'hbbf;
rom[10084] = 12'hbbf;
rom[10085] = 12'haae;
rom[10086] = 12'haae;
rom[10087] = 12'haae;
rom[10088] = 12'haae;
rom[10089] = 12'haae;
rom[10090] = 12'hbbf;
rom[10091] = 12'hbbf;
rom[10092] = 12'hbbf;
rom[10093] = 12'hccf;
rom[10094] = 12'hddf;
rom[10095] = 12'heef;
rom[10096] = 12'hfff;
rom[10097] = 12'hfff;
rom[10098] = 12'hfff;
rom[10099] = 12'hfff;
rom[10100] = 12'hfff;
rom[10101] = 12'hfff;
rom[10102] = 12'hfff;
rom[10103] = 12'hfff;
rom[10104] = 12'hfff;
rom[10105] = 12'hfff;
rom[10106] = 12'hfff;
rom[10107] = 12'hfff;
rom[10108] = 12'hfff;
rom[10109] = 12'hfff;
rom[10110] = 12'hfff;
rom[10111] = 12'hfff;
rom[10112] = 12'hfff;
rom[10113] = 12'hfff;
rom[10114] = 12'hfff;
rom[10115] = 12'hfff;
rom[10116] = 12'hfff;
rom[10117] = 12'hfff;
rom[10118] = 12'hfff;
rom[10119] = 12'hfff;
rom[10120] = 12'hfff;
rom[10121] = 12'hfff;
rom[10122] = 12'hfff;
rom[10123] = 12'hfff;
rom[10124] = 12'hfff;
rom[10125] = 12'hfff;
rom[10126] = 12'hfff;
rom[10127] = 12'hfff;
rom[10128] = 12'hfff;
rom[10129] = 12'hfff;
rom[10130] = 12'hfff;
rom[10131] = 12'hfff;
rom[10132] = 12'hfff;
rom[10133] = 12'heef;
rom[10134] = 12'h  c;
rom[10135] = 12'h  c;
rom[10136] = 12'h  c;
rom[10137] = 12'h  c;
rom[10138] = 12'h  c;
rom[10139] = 12'h  c;
rom[10140] = 12'h  c;
rom[10141] = 12'h  c;
rom[10142] = 12'h33d;
rom[10143] = 12'h99e;
rom[10144] = 12'hccf;
rom[10145] = 12'hddf;
rom[10146] = 12'hddf;
rom[10147] = 12'heef;
rom[10148] = 12'heef;
rom[10149] = 12'heef;
rom[10150] = 12'heef;
rom[10151] = 12'heef;
rom[10152] = 12'heef;
rom[10153] = 12'hddf;
rom[10154] = 12'hddf;
rom[10155] = 12'hccf;
rom[10156] = 12'h99e;
rom[10157] = 12'h33d;
rom[10158] = 12'h  c;
rom[10159] = 12'h  c;
rom[10160] = 12'h  c;
rom[10161] = 12'h  c;
rom[10162] = 12'h  c;
rom[10163] = 12'h  c;
rom[10164] = 12'h99e;
rom[10165] = 12'hfff;
rom[10166] = 12'hfff;
rom[10167] = 12'hfff;
rom[10168] = 12'hfff;
rom[10169] = 12'hfff;
rom[10170] = 12'h11d;
rom[10171] = 12'h  c;
rom[10172] = 12'h  c;
rom[10173] = 12'h  c;
rom[10174] = 12'h  c;
rom[10175] = 12'hddf;
rom[10176] = 12'hfff;
rom[10177] = 12'hfff;
rom[10178] = 12'hfff;
rom[10179] = 12'hfff;
rom[10180] = 12'hfff;
rom[10181] = 12'hfff;
rom[10182] = 12'hfff;
rom[10183] = 12'hfff;
rom[10184] = 12'hfff;
rom[10185] = 12'hfff;
rom[10186] = 12'hfff;
rom[10187] = 12'hfff;
rom[10188] = 12'hfff;
rom[10189] = 12'hfff;
rom[10190] = 12'hfff;
rom[10191] = 12'hfff;
rom[10192] = 12'hfff;
rom[10193] = 12'hfff;
rom[10194] = 12'hfff;
rom[10195] = 12'hfff;
rom[10196] = 12'hfff;
rom[10197] = 12'hfff;
rom[10198] = 12'hfff;
rom[10199] = 12'hfff;
rom[10200] = 12'h66e;
rom[10201] = 12'h  c;
rom[10202] = 12'h  c;
rom[10203] = 12'h  c;
rom[10204] = 12'h  c;
rom[10205] = 12'h66e;
rom[10206] = 12'heef;
rom[10207] = 12'hfff;
rom[10208] = 12'hfff;
rom[10209] = 12'hfff;
rom[10210] = 12'hfff;
rom[10211] = 12'hfff;
rom[10212] = 12'hfff;
rom[10213] = 12'hfff;
rom[10214] = 12'hfff;
rom[10215] = 12'hfff;
rom[10216] = 12'hfff;
rom[10217] = 12'hfff;
rom[10218] = 12'hfff;
rom[10219] = 12'hfff;
rom[10220] = 12'hfff;
rom[10221] = 12'hfff;
rom[10222] = 12'hfff;
rom[10223] = 12'hfff;
rom[10224] = 12'hfff;
rom[10225] = 12'hfff;
rom[10226] = 12'hfff;
rom[10227] = 12'hfff;
rom[10228] = 12'hfff;
rom[10229] = 12'hfff;
rom[10230] = 12'hfff;
rom[10231] = 12'hfff;
rom[10232] = 12'hfff;
rom[10233] = 12'hfff;
rom[10234] = 12'hfff;
rom[10235] = 12'hfff;
rom[10236] = 12'hfff;
rom[10237] = 12'hfff;
rom[10238] = 12'hfff;
rom[10239] = 12'hfff;
rom[10240] = 12'hfff;
rom[10241] = 12'hfff;
rom[10242] = 12'hfff;
rom[10243] = 12'hfff;
rom[10244] = 12'hfff;
rom[10245] = 12'hfff;
rom[10246] = 12'hfff;
rom[10247] = 12'hfff;
rom[10248] = 12'hfff;
rom[10249] = 12'hfff;
rom[10250] = 12'hfff;
rom[10251] = 12'hfff;
rom[10252] = 12'hfff;
rom[10253] = 12'hfff;
rom[10254] = 12'hfff;
rom[10255] = 12'hfff;
rom[10256] = 12'hfff;
rom[10257] = 12'hfff;
rom[10258] = 12'hfff;
rom[10259] = 12'hfff;
rom[10260] = 12'heef;
rom[10261] = 12'h44d;
rom[10262] = 12'h  c;
rom[10263] = 12'h  c;
rom[10264] = 12'h  c;
rom[10265] = 12'h  c;
rom[10266] = 12'h  c;
rom[10267] = 12'h33d;
rom[10268] = 12'h99e;
rom[10269] = 12'haae;
rom[10270] = 12'hfff;
rom[10271] = 12'hfff;
rom[10272] = 12'hfff;
rom[10273] = 12'hfff;
rom[10274] = 12'hfff;
rom[10275] = 12'hfff;
rom[10276] = 12'hfff;
rom[10277] = 12'hfff;
rom[10278] = 12'hfff;
rom[10279] = 12'hfff;
rom[10280] = 12'hfff;
rom[10281] = 12'hfff;
rom[10282] = 12'hfff;
rom[10283] = 12'hfff;
rom[10284] = 12'hfff;
rom[10285] = 12'hfff;
rom[10286] = 12'haae;
rom[10287] = 12'h99e;
rom[10288] = 12'h22d;
rom[10289] = 12'h  c;
rom[10290] = 12'h  c;
rom[10291] = 12'h11d;
rom[10292] = 12'heef;
rom[10293] = 12'hfff;
rom[10294] = 12'hfff;
rom[10295] = 12'hfff;
rom[10296] = 12'hfff;
rom[10297] = 12'hfff;
rom[10298] = 12'h33d;
rom[10299] = 12'h  c;
rom[10300] = 12'h  c;
rom[10301] = 12'h  c;
rom[10302] = 12'h  c;
rom[10303] = 12'hccf;
rom[10304] = 12'hfff;
rom[10305] = 12'hfff;
rom[10306] = 12'hfff;
rom[10307] = 12'hfff;
rom[10308] = 12'hfff;
rom[10309] = 12'hfff;
rom[10310] = 12'hfff;
rom[10311] = 12'hfff;
rom[10312] = 12'hfff;
rom[10313] = 12'hfff;
rom[10314] = 12'hfff;
rom[10315] = 12'hfff;
rom[10316] = 12'hfff;
rom[10317] = 12'hfff;
rom[10318] = 12'hfff;
rom[10319] = 12'hfff;
rom[10320] = 12'hfff;
rom[10321] = 12'hfff;
rom[10322] = 12'hfff;
rom[10323] = 12'hfff;
rom[10324] = 12'hfff;
rom[10325] = 12'hfff;
rom[10326] = 12'hfff;
rom[10327] = 12'hfff;
rom[10328] = 12'h99e;
rom[10329] = 12'h  c;
rom[10330] = 12'h  c;
rom[10331] = 12'h  c;
rom[10332] = 12'h  c;
rom[10333] = 12'h22d;
rom[10334] = 12'h88e;
rom[10335] = 12'hfff;
rom[10336] = 12'hfff;
rom[10337] = 12'hfff;
rom[10338] = 12'hfff;
rom[10339] = 12'hfff;
rom[10340] = 12'hfff;
rom[10341] = 12'hfff;
rom[10342] = 12'hfff;
rom[10343] = 12'hfff;
rom[10344] = 12'hfff;
rom[10345] = 12'hfff;
rom[10346] = 12'hfff;
rom[10347] = 12'hfff;
rom[10348] = 12'hfff;
rom[10349] = 12'hfff;
rom[10350] = 12'hfff;
rom[10351] = 12'hfff;
rom[10352] = 12'hfff;
rom[10353] = 12'hfff;
rom[10354] = 12'hfff;
rom[10355] = 12'hfff;
rom[10356] = 12'hfff;
rom[10357] = 12'hfff;
rom[10358] = 12'hfff;
rom[10359] = 12'hfff;
rom[10360] = 12'hfff;
rom[10361] = 12'hfff;
rom[10362] = 12'hfff;
rom[10363] = 12'hfff;
rom[10364] = 12'hfff;
rom[10365] = 12'hfff;
rom[10366] = 12'hfff;
rom[10367] = 12'hfff;
rom[10368] = 12'hfff;
rom[10369] = 12'hfff;
rom[10370] = 12'hfff;
rom[10371] = 12'hfff;
rom[10372] = 12'hfff;
rom[10373] = 12'hfff;
rom[10374] = 12'hfff;
rom[10375] = 12'hfff;
rom[10376] = 12'hfff;
rom[10377] = 12'hfff;
rom[10378] = 12'hfff;
rom[10379] = 12'hfff;
rom[10380] = 12'hfff;
rom[10381] = 12'hfff;
rom[10382] = 12'hfff;
rom[10383] = 12'hfff;
rom[10384] = 12'hfff;
rom[10385] = 12'hfff;
rom[10386] = 12'hfff;
rom[10387] = 12'heef;
rom[10388] = 12'h11d;
rom[10389] = 12'h  c;
rom[10390] = 12'h  c;
rom[10391] = 12'h  c;
rom[10392] = 12'h  c;
rom[10393] = 12'h11d;
rom[10394] = 12'hbbf;
rom[10395] = 12'hfff;
rom[10396] = 12'hfff;
rom[10397] = 12'hfff;
rom[10398] = 12'hfff;
rom[10399] = 12'hfff;
rom[10400] = 12'hfff;
rom[10401] = 12'hfff;
rom[10402] = 12'hfff;
rom[10403] = 12'hfff;
rom[10404] = 12'hfff;
rom[10405] = 12'hfff;
rom[10406] = 12'hfff;
rom[10407] = 12'hfff;
rom[10408] = 12'hfff;
rom[10409] = 12'hfff;
rom[10410] = 12'hfff;
rom[10411] = 12'hfff;
rom[10412] = 12'hfff;
rom[10413] = 12'hfff;
rom[10414] = 12'hfff;
rom[10415] = 12'hfff;
rom[10416] = 12'heef;
rom[10417] = 12'h99e;
rom[10418] = 12'h99e;
rom[10419] = 12'heef;
rom[10420] = 12'hfff;
rom[10421] = 12'hfff;
rom[10422] = 12'hfff;
rom[10423] = 12'hfff;
rom[10424] = 12'hfff;
rom[10425] = 12'hfff;
rom[10426] = 12'h44d;
rom[10427] = 12'h  c;
rom[10428] = 12'h  c;
rom[10429] = 12'h  c;
rom[10430] = 12'h  c;
rom[10431] = 12'hbbf;
rom[10432] = 12'hfff;
rom[10433] = 12'hfff;
rom[10434] = 12'hfff;
rom[10435] = 12'hfff;
rom[10436] = 12'hfff;
rom[10437] = 12'hfff;
rom[10438] = 12'hfff;
rom[10439] = 12'hfff;
rom[10440] = 12'hfff;
rom[10441] = 12'hfff;
rom[10442] = 12'hfff;
rom[10443] = 12'hfff;
rom[10444] = 12'hfff;
rom[10445] = 12'hfff;
rom[10446] = 12'hfff;
rom[10447] = 12'hfff;
rom[10448] = 12'hfff;
rom[10449] = 12'hfff;
rom[10450] = 12'hfff;
rom[10451] = 12'hfff;
rom[10452] = 12'hfff;
rom[10453] = 12'hfff;
rom[10454] = 12'hfff;
rom[10455] = 12'hfff;
rom[10456] = 12'heef;
rom[10457] = 12'h11d;
rom[10458] = 12'h  c;
rom[10459] = 12'h  c;
rom[10460] = 12'h  c;
rom[10461] = 12'h  c;
rom[10462] = 12'h  c;
rom[10463] = 12'h99e;
rom[10464] = 12'hfff;
rom[10465] = 12'hfff;
rom[10466] = 12'hfff;
rom[10467] = 12'hfff;
rom[10468] = 12'hfff;
rom[10469] = 12'hfff;
rom[10470] = 12'hfff;
rom[10471] = 12'hfff;
rom[10472] = 12'hfff;
rom[10473] = 12'hfff;
rom[10474] = 12'hfff;
rom[10475] = 12'hfff;
rom[10476] = 12'hfff;
rom[10477] = 12'hfff;
rom[10478] = 12'hfff;
rom[10479] = 12'hfff;
rom[10480] = 12'hfff;
rom[10481] = 12'hfff;
rom[10482] = 12'hfff;
rom[10483] = 12'hfff;
rom[10484] = 12'hfff;
rom[10485] = 12'hfff;
rom[10486] = 12'hfff;
rom[10487] = 12'hfff;
rom[10488] = 12'hfff;
rom[10489] = 12'hfff;
rom[10490] = 12'hfff;
rom[10491] = 12'hfff;
rom[10492] = 12'hfff;
rom[10493] = 12'hfff;
rom[10494] = 12'hfff;
rom[10495] = 12'hfff;
rom[10496] = 12'hfff;
rom[10497] = 12'hfff;
rom[10498] = 12'hfff;
rom[10499] = 12'hfff;
rom[10500] = 12'hfff;
rom[10501] = 12'hfff;
rom[10502] = 12'hfff;
rom[10503] = 12'hfff;
rom[10504] = 12'hfff;
rom[10505] = 12'hfff;
rom[10506] = 12'hfff;
rom[10507] = 12'hfff;
rom[10508] = 12'hfff;
rom[10509] = 12'hfff;
rom[10510] = 12'hfff;
rom[10511] = 12'hfff;
rom[10512] = 12'hfff;
rom[10513] = 12'hfff;
rom[10514] = 12'hfff;
rom[10515] = 12'h99e;
rom[10516] = 12'h  c;
rom[10517] = 12'h  c;
rom[10518] = 12'h  c;
rom[10519] = 12'h  c;
rom[10520] = 12'h  c;
rom[10521] = 12'h88e;
rom[10522] = 12'hfff;
rom[10523] = 12'hfff;
rom[10524] = 12'hfff;
rom[10525] = 12'hfff;
rom[10526] = 12'hfff;
rom[10527] = 12'hfff;
rom[10528] = 12'hfff;
rom[10529] = 12'hfff;
rom[10530] = 12'hfff;
rom[10531] = 12'hfff;
rom[10532] = 12'hfff;
rom[10533] = 12'hfff;
rom[10534] = 12'hfff;
rom[10535] = 12'hfff;
rom[10536] = 12'hfff;
rom[10537] = 12'hfff;
rom[10538] = 12'hfff;
rom[10539] = 12'hfff;
rom[10540] = 12'hfff;
rom[10541] = 12'hfff;
rom[10542] = 12'hfff;
rom[10543] = 12'hfff;
rom[10544] = 12'hfff;
rom[10545] = 12'hfff;
rom[10546] = 12'hfff;
rom[10547] = 12'hfff;
rom[10548] = 12'hfff;
rom[10549] = 12'hfff;
rom[10550] = 12'hfff;
rom[10551] = 12'hfff;
rom[10552] = 12'hfff;
rom[10553] = 12'hfff;
rom[10554] = 12'h55d;
rom[10555] = 12'h  c;
rom[10556] = 12'h  c;
rom[10557] = 12'h  c;
rom[10558] = 12'h  c;
rom[10559] = 12'haae;
rom[10560] = 12'hfff;
rom[10561] = 12'hfff;
rom[10562] = 12'hfff;
rom[10563] = 12'hfff;
rom[10564] = 12'hfff;
rom[10565] = 12'hfff;
rom[10566] = 12'hfff;
rom[10567] = 12'hfff;
rom[10568] = 12'hfff;
rom[10569] = 12'hfff;
rom[10570] = 12'hfff;
rom[10571] = 12'hfff;
rom[10572] = 12'hfff;
rom[10573] = 12'hfff;
rom[10574] = 12'hfff;
rom[10575] = 12'hfff;
rom[10576] = 12'hfff;
rom[10577] = 12'hfff;
rom[10578] = 12'hfff;
rom[10579] = 12'hfff;
rom[10580] = 12'hfff;
rom[10581] = 12'hfff;
rom[10582] = 12'hfff;
rom[10583] = 12'hfff;
rom[10584] = 12'hfff;
rom[10585] = 12'hddf;
rom[10586] = 12'h11d;
rom[10587] = 12'h  c;
rom[10588] = 12'h  c;
rom[10589] = 12'h  c;
rom[10590] = 12'h  c;
rom[10591] = 12'h88e;
rom[10592] = 12'hfff;
rom[10593] = 12'hfff;
rom[10594] = 12'hfff;
rom[10595] = 12'hfff;
rom[10596] = 12'hfff;
rom[10597] = 12'hfff;
rom[10598] = 12'hfff;
rom[10599] = 12'hfff;
rom[10600] = 12'hfff;
rom[10601] = 12'hfff;
rom[10602] = 12'hfff;
rom[10603] = 12'hfff;
rom[10604] = 12'hfff;
rom[10605] = 12'hfff;
rom[10606] = 12'hfff;
rom[10607] = 12'hfff;
rom[10608] = 12'hfff;
rom[10609] = 12'hfff;
rom[10610] = 12'hfff;
rom[10611] = 12'hfff;
rom[10612] = 12'hfff;
rom[10613] = 12'hfff;
rom[10614] = 12'hfff;
rom[10615] = 12'hfff;
rom[10616] = 12'hfff;
rom[10617] = 12'hfff;
rom[10618] = 12'hfff;
rom[10619] = 12'hfff;
rom[10620] = 12'hfff;
rom[10621] = 12'hfff;
rom[10622] = 12'hfff;
rom[10623] = 12'hfff;
rom[10624] = 12'hfff;
rom[10625] = 12'hfff;
rom[10626] = 12'hfff;
rom[10627] = 12'hfff;
rom[10628] = 12'hfff;
rom[10629] = 12'hfff;
rom[10630] = 12'hfff;
rom[10631] = 12'hfff;
rom[10632] = 12'hfff;
rom[10633] = 12'hfff;
rom[10634] = 12'hfff;
rom[10635] = 12'hfff;
rom[10636] = 12'hfff;
rom[10637] = 12'hfff;
rom[10638] = 12'hfff;
rom[10639] = 12'hfff;
rom[10640] = 12'hfff;
rom[10641] = 12'hfff;
rom[10642] = 12'heef;
rom[10643] = 12'h22d;
rom[10644] = 12'h  c;
rom[10645] = 12'h  c;
rom[10646] = 12'h  c;
rom[10647] = 12'h  c;
rom[10648] = 12'h  c;
rom[10649] = 12'haae;
rom[10650] = 12'hfff;
rom[10651] = 12'hfff;
rom[10652] = 12'hfff;
rom[10653] = 12'hfff;
rom[10654] = 12'hfff;
rom[10655] = 12'hfff;
rom[10656] = 12'hfff;
rom[10657] = 12'hfff;
rom[10658] = 12'hfff;
rom[10659] = 12'hfff;
rom[10660] = 12'hfff;
rom[10661] = 12'hfff;
rom[10662] = 12'hfff;
rom[10663] = 12'hfff;
rom[10664] = 12'hfff;
rom[10665] = 12'hfff;
rom[10666] = 12'hfff;
rom[10667] = 12'hfff;
rom[10668] = 12'hfff;
rom[10669] = 12'hfff;
rom[10670] = 12'hfff;
rom[10671] = 12'hfff;
rom[10672] = 12'hfff;
rom[10673] = 12'hfff;
rom[10674] = 12'hfff;
rom[10675] = 12'hfff;
rom[10676] = 12'hfff;
rom[10677] = 12'hfff;
rom[10678] = 12'hfff;
rom[10679] = 12'hfff;
rom[10680] = 12'hfff;
rom[10681] = 12'hfff;
rom[10682] = 12'h66d;
rom[10683] = 12'h  c;
rom[10684] = 12'h  c;
rom[10685] = 12'h  c;
rom[10686] = 12'h  c;
rom[10687] = 12'h99e;
rom[10688] = 12'hfff;
rom[10689] = 12'hfff;
rom[10690] = 12'hfff;
rom[10691] = 12'hfff;
rom[10692] = 12'hfff;
rom[10693] = 12'hfff;
rom[10694] = 12'hfff;
rom[10695] = 12'hfff;
rom[10696] = 12'hfff;
rom[10697] = 12'hfff;
rom[10698] = 12'hfff;
rom[10699] = 12'hfff;
rom[10700] = 12'hfff;
rom[10701] = 12'hfff;
rom[10702] = 12'hfff;
rom[10703] = 12'hfff;
rom[10704] = 12'hfff;
rom[10705] = 12'hfff;
rom[10706] = 12'hfff;
rom[10707] = 12'hfff;
rom[10708] = 12'hfff;
rom[10709] = 12'hfff;
rom[10710] = 12'hfff;
rom[10711] = 12'hfff;
rom[10712] = 12'hfff;
rom[10713] = 12'hfff;
rom[10714] = 12'hbbe;
rom[10715] = 12'h11d;
rom[10716] = 12'h  c;
rom[10717] = 12'h  c;
rom[10718] = 12'h  c;
rom[10719] = 12'h55d;
rom[10720] = 12'hfff;
rom[10721] = 12'hfff;
rom[10722] = 12'hfff;
rom[10723] = 12'hfff;
rom[10724] = 12'hfff;
rom[10725] = 12'hfff;
rom[10726] = 12'hfff;
rom[10727] = 12'hfff;
rom[10728] = 12'hfff;
rom[10729] = 12'hfff;
rom[10730] = 12'hfff;
rom[10731] = 12'hfff;
rom[10732] = 12'hfff;
rom[10733] = 12'hfff;
rom[10734] = 12'hfff;
rom[10735] = 12'hfff;
rom[10736] = 12'hfff;
rom[10737] = 12'hfff;
rom[10738] = 12'hfff;
rom[10739] = 12'hfff;
rom[10740] = 12'hfff;
rom[10741] = 12'hfff;
rom[10742] = 12'hfff;
rom[10743] = 12'hfff;
rom[10744] = 12'hfff;
rom[10745] = 12'hfff;
rom[10746] = 12'hfff;
rom[10747] = 12'hfff;
rom[10748] = 12'hfff;
rom[10749] = 12'hfff;
rom[10750] = 12'hfff;
rom[10751] = 12'hfff;
rom[10752] = 12'hfff;
rom[10753] = 12'hfff;
rom[10754] = 12'hfff;
rom[10755] = 12'hfff;
rom[10756] = 12'hfff;
rom[10757] = 12'hfff;
rom[10758] = 12'hfff;
rom[10759] = 12'hfff;
rom[10760] = 12'hfff;
rom[10761] = 12'hfff;
rom[10762] = 12'hfff;
rom[10763] = 12'hfff;
rom[10764] = 12'hfff;
rom[10765] = 12'hfff;
rom[10766] = 12'hfff;
rom[10767] = 12'hfff;
rom[10768] = 12'hfff;
rom[10769] = 12'hfff;
rom[10770] = 12'h88e;
rom[10771] = 12'h  c;
rom[10772] = 12'h  c;
rom[10773] = 12'h  c;
rom[10774] = 12'h  c;
rom[10775] = 12'h  c;
rom[10776] = 12'h11d;
rom[10777] = 12'heef;
rom[10778] = 12'hfff;
rom[10779] = 12'hfff;
rom[10780] = 12'hfff;
rom[10781] = 12'hfff;
rom[10782] = 12'hfff;
rom[10783] = 12'hfff;
rom[10784] = 12'hfff;
rom[10785] = 12'hfff;
rom[10786] = 12'hfff;
rom[10787] = 12'hfff;
rom[10788] = 12'hfff;
rom[10789] = 12'hfff;
rom[10790] = 12'hfff;
rom[10791] = 12'hfff;
rom[10792] = 12'hfff;
rom[10793] = 12'hfff;
rom[10794] = 12'hfff;
rom[10795] = 12'hfff;
rom[10796] = 12'hfff;
rom[10797] = 12'hfff;
rom[10798] = 12'hfff;
rom[10799] = 12'hfff;
rom[10800] = 12'hfff;
rom[10801] = 12'hfff;
rom[10802] = 12'hfff;
rom[10803] = 12'hfff;
rom[10804] = 12'hfff;
rom[10805] = 12'hfff;
rom[10806] = 12'hfff;
rom[10807] = 12'hfff;
rom[10808] = 12'hfff;
rom[10809] = 12'hfff;
rom[10810] = 12'h66e;
rom[10811] = 12'h  c;
rom[10812] = 12'h  c;
rom[10813] = 12'h  c;
rom[10814] = 12'h  c;
rom[10815] = 12'h99e;
rom[10816] = 12'hfff;
rom[10817] = 12'hfff;
rom[10818] = 12'hfff;
rom[10819] = 12'hfff;
rom[10820] = 12'hfff;
rom[10821] = 12'hfff;
rom[10822] = 12'hfff;
rom[10823] = 12'hfff;
rom[10824] = 12'hfff;
rom[10825] = 12'hfff;
rom[10826] = 12'hfff;
rom[10827] = 12'hfff;
rom[10828] = 12'hfff;
rom[10829] = 12'hfff;
rom[10830] = 12'hfff;
rom[10831] = 12'hfff;
rom[10832] = 12'hfff;
rom[10833] = 12'hfff;
rom[10834] = 12'hfff;
rom[10835] = 12'hfff;
rom[10836] = 12'hfff;
rom[10837] = 12'hfff;
rom[10838] = 12'hfff;
rom[10839] = 12'hfff;
rom[10840] = 12'hfff;
rom[10841] = 12'hfff;
rom[10842] = 12'hddf;
rom[10843] = 12'h11d;
rom[10844] = 12'h  c;
rom[10845] = 12'h  c;
rom[10846] = 12'h  c;
rom[10847] = 12'h11d;
rom[10848] = 12'hddf;
rom[10849] = 12'hfff;
rom[10850] = 12'hfff;
rom[10851] = 12'hfff;
rom[10852] = 12'hfff;
rom[10853] = 12'hfff;
rom[10854] = 12'hfff;
rom[10855] = 12'hfff;
rom[10856] = 12'hfff;
rom[10857] = 12'hfff;
rom[10858] = 12'hfff;
rom[10859] = 12'hfff;
rom[10860] = 12'hfff;
rom[10861] = 12'hfff;
rom[10862] = 12'hfff;
rom[10863] = 12'hfff;
rom[10864] = 12'hfff;
rom[10865] = 12'hfff;
rom[10866] = 12'hfff;
rom[10867] = 12'hfff;
rom[10868] = 12'hfff;
rom[10869] = 12'hfff;
rom[10870] = 12'hfff;
rom[10871] = 12'hfff;
rom[10872] = 12'hfff;
rom[10873] = 12'hfff;
rom[10874] = 12'hfff;
rom[10875] = 12'hfff;
rom[10876] = 12'hfff;
rom[10877] = 12'hfff;
rom[10878] = 12'hfff;
rom[10879] = 12'hfff;
rom[10880] = 12'hfff;
rom[10881] = 12'hfff;
rom[10882] = 12'hfff;
rom[10883] = 12'hfff;
rom[10884] = 12'hfff;
rom[10885] = 12'hfff;
rom[10886] = 12'hfff;
rom[10887] = 12'hfff;
rom[10888] = 12'hfff;
rom[10889] = 12'hfff;
rom[10890] = 12'hfff;
rom[10891] = 12'hfff;
rom[10892] = 12'hfff;
rom[10893] = 12'hfff;
rom[10894] = 12'hfff;
rom[10895] = 12'hfff;
rom[10896] = 12'hfff;
rom[10897] = 12'hfff;
rom[10898] = 12'h33d;
rom[10899] = 12'h  c;
rom[10900] = 12'h  c;
rom[10901] = 12'h  c;
rom[10902] = 12'h11d;
rom[10903] = 12'h44d;
rom[10904] = 12'heef;
rom[10905] = 12'hfff;
rom[10906] = 12'hfff;
rom[10907] = 12'hfff;
rom[10908] = 12'hfff;
rom[10909] = 12'hfff;
rom[10910] = 12'hfff;
rom[10911] = 12'hfff;
rom[10912] = 12'hfff;
rom[10913] = 12'hfff;
rom[10914] = 12'hfff;
rom[10915] = 12'hfff;
rom[10916] = 12'hfff;
rom[10917] = 12'hfff;
rom[10918] = 12'hfff;
rom[10919] = 12'hfff;
rom[10920] = 12'hfff;
rom[10921] = 12'hfff;
rom[10922] = 12'hfff;
rom[10923] = 12'hfff;
rom[10924] = 12'hfff;
rom[10925] = 12'hfff;
rom[10926] = 12'hfff;
rom[10927] = 12'hfff;
rom[10928] = 12'hfff;
rom[10929] = 12'hfff;
rom[10930] = 12'hfff;
rom[10931] = 12'hfff;
rom[10932] = 12'hfff;
rom[10933] = 12'hfff;
rom[10934] = 12'hfff;
rom[10935] = 12'hfff;
rom[10936] = 12'hfff;
rom[10937] = 12'hfff;
rom[10938] = 12'h66e;
rom[10939] = 12'h  c;
rom[10940] = 12'h  c;
rom[10941] = 12'h  c;
rom[10942] = 12'h  c;
rom[10943] = 12'h99e;
rom[10944] = 12'hfff;
rom[10945] = 12'hfff;
rom[10946] = 12'hfff;
rom[10947] = 12'hfff;
rom[10948] = 12'hfff;
rom[10949] = 12'hfff;
rom[10950] = 12'hfff;
rom[10951] = 12'hfff;
rom[10952] = 12'hfff;
rom[10953] = 12'hfff;
rom[10954] = 12'hfff;
rom[10955] = 12'hfff;
rom[10956] = 12'hfff;
rom[10957] = 12'hfff;
rom[10958] = 12'hfff;
rom[10959] = 12'hfff;
rom[10960] = 12'hfff;
rom[10961] = 12'hfff;
rom[10962] = 12'hfff;
rom[10963] = 12'hfff;
rom[10964] = 12'hfff;
rom[10965] = 12'hfff;
rom[10966] = 12'hfff;
rom[10967] = 12'hfff;
rom[10968] = 12'hfff;
rom[10969] = 12'hfff;
rom[10970] = 12'hfff;
rom[10971] = 12'h66e;
rom[10972] = 12'h  c;
rom[10973] = 12'h  c;
rom[10974] = 12'h  c;
rom[10975] = 12'h  c;
rom[10976] = 12'h88e;
rom[10977] = 12'heef;
rom[10978] = 12'hfff;
rom[10979] = 12'hfff;
rom[10980] = 12'hfff;
rom[10981] = 12'hfff;
rom[10982] = 12'hfff;
rom[10983] = 12'hfff;
rom[10984] = 12'hfff;
rom[10985] = 12'hfff;
rom[10986] = 12'hfff;
rom[10987] = 12'hfff;
rom[10988] = 12'hfff;
rom[10989] = 12'hfff;
rom[10990] = 12'hfff;
rom[10991] = 12'hfff;
rom[10992] = 12'hfff;
rom[10993] = 12'hfff;
rom[10994] = 12'hfff;
rom[10995] = 12'hfff;
rom[10996] = 12'hfff;
rom[10997] = 12'hfff;
rom[10998] = 12'hfff;
rom[10999] = 12'hfff;
rom[11000] = 12'hfff;
rom[11001] = 12'hfff;
rom[11002] = 12'hfff;
rom[11003] = 12'hfff;
rom[11004] = 12'hfff;
rom[11005] = 12'hfff;
rom[11006] = 12'hfff;
rom[11007] = 12'hfff;
rom[11008] = 12'hfff;
rom[11009] = 12'hfff;
rom[11010] = 12'hfff;
rom[11011] = 12'hfff;
rom[11012] = 12'hfff;
rom[11013] = 12'hfff;
rom[11014] = 12'hfff;
rom[11015] = 12'hfff;
rom[11016] = 12'hfff;
rom[11017] = 12'hfff;
rom[11018] = 12'hfff;
rom[11019] = 12'hfff;
rom[11020] = 12'hfff;
rom[11021] = 12'hfff;
rom[11022] = 12'hfff;
rom[11023] = 12'hfff;
rom[11024] = 12'hfff;
rom[11025] = 12'hfff;
rom[11026] = 12'h11d;
rom[11027] = 12'h  c;
rom[11028] = 12'h  c;
rom[11029] = 12'h  c;
rom[11030] = 12'h  c;
rom[11031] = 12'hddf;
rom[11032] = 12'hfff;
rom[11033] = 12'hfff;
rom[11034] = 12'hfff;
rom[11035] = 12'hfff;
rom[11036] = 12'hfff;
rom[11037] = 12'hfff;
rom[11038] = 12'hfff;
rom[11039] = 12'hfff;
rom[11040] = 12'hfff;
rom[11041] = 12'hfff;
rom[11042] = 12'hfff;
rom[11043] = 12'hfff;
rom[11044] = 12'hfff;
rom[11045] = 12'hfff;
rom[11046] = 12'hfff;
rom[11047] = 12'hfff;
rom[11048] = 12'hfff;
rom[11049] = 12'hfff;
rom[11050] = 12'hfff;
rom[11051] = 12'hfff;
rom[11052] = 12'hfff;
rom[11053] = 12'hfff;
rom[11054] = 12'hfff;
rom[11055] = 12'hfff;
rom[11056] = 12'hfff;
rom[11057] = 12'hfff;
rom[11058] = 12'hfff;
rom[11059] = 12'hfff;
rom[11060] = 12'hfff;
rom[11061] = 12'hfff;
rom[11062] = 12'hfff;
rom[11063] = 12'hfff;
rom[11064] = 12'hfff;
rom[11065] = 12'hfff;
rom[11066] = 12'h66e;
rom[11067] = 12'h  c;
rom[11068] = 12'h  c;
rom[11069] = 12'h  c;
rom[11070] = 12'h  c;
rom[11071] = 12'h99e;
rom[11072] = 12'hfff;
rom[11073] = 12'hfff;
rom[11074] = 12'hfff;
rom[11075] = 12'hfff;
rom[11076] = 12'hfff;
rom[11077] = 12'hfff;
rom[11078] = 12'hfff;
rom[11079] = 12'hfff;
rom[11080] = 12'hfff;
rom[11081] = 12'hfff;
rom[11082] = 12'hfff;
rom[11083] = 12'hfff;
rom[11084] = 12'hfff;
rom[11085] = 12'hfff;
rom[11086] = 12'hfff;
rom[11087] = 12'hfff;
rom[11088] = 12'hfff;
rom[11089] = 12'hfff;
rom[11090] = 12'hfff;
rom[11091] = 12'hfff;
rom[11092] = 12'hfff;
rom[11093] = 12'hfff;
rom[11094] = 12'hfff;
rom[11095] = 12'hfff;
rom[11096] = 12'hfff;
rom[11097] = 12'hfff;
rom[11098] = 12'hfff;
rom[11099] = 12'h99e;
rom[11100] = 12'h  c;
rom[11101] = 12'h  c;
rom[11102] = 12'h  c;
rom[11103] = 12'h  c;
rom[11104] = 12'h22d;
rom[11105] = 12'h44d;
rom[11106] = 12'hfff;
rom[11107] = 12'hfff;
rom[11108] = 12'hfff;
rom[11109] = 12'hfff;
rom[11110] = 12'hfff;
rom[11111] = 12'hfff;
rom[11112] = 12'hfff;
rom[11113] = 12'hfff;
rom[11114] = 12'hfff;
rom[11115] = 12'hfff;
rom[11116] = 12'hfff;
rom[11117] = 12'hfff;
rom[11118] = 12'hfff;
rom[11119] = 12'hfff;
rom[11120] = 12'hfff;
rom[11121] = 12'hfff;
rom[11122] = 12'hfff;
rom[11123] = 12'hfff;
rom[11124] = 12'hfff;
rom[11125] = 12'hfff;
rom[11126] = 12'hfff;
rom[11127] = 12'hfff;
rom[11128] = 12'hfff;
rom[11129] = 12'hfff;
rom[11130] = 12'hfff;
rom[11131] = 12'hfff;
rom[11132] = 12'hfff;
rom[11133] = 12'hfff;
rom[11134] = 12'hfff;
rom[11135] = 12'hfff;
rom[11136] = 12'hfff;
rom[11137] = 12'hfff;
rom[11138] = 12'hfff;
rom[11139] = 12'hfff;
rom[11140] = 12'hfff;
rom[11141] = 12'hfff;
rom[11142] = 12'hfff;
rom[11143] = 12'hfff;
rom[11144] = 12'hfff;
rom[11145] = 12'hfff;
rom[11146] = 12'hfff;
rom[11147] = 12'hfff;
rom[11148] = 12'hfff;
rom[11149] = 12'hfff;
rom[11150] = 12'hfff;
rom[11151] = 12'hfff;
rom[11152] = 12'hfff;
rom[11153] = 12'hfff;
rom[11154] = 12'h  c;
rom[11155] = 12'h  c;
rom[11156] = 12'h  c;
rom[11157] = 12'h  c;
rom[11158] = 12'h  c;
rom[11159] = 12'hfff;
rom[11160] = 12'hfff;
rom[11161] = 12'hfff;
rom[11162] = 12'hfff;
rom[11163] = 12'hfff;
rom[11164] = 12'hfff;
rom[11165] = 12'hfff;
rom[11166] = 12'hfff;
rom[11167] = 12'hfff;
rom[11168] = 12'hfff;
rom[11169] = 12'hfff;
rom[11170] = 12'hfff;
rom[11171] = 12'hfff;
rom[11172] = 12'hfff;
rom[11173] = 12'hfff;
rom[11174] = 12'hfff;
rom[11175] = 12'hfff;
rom[11176] = 12'hfff;
rom[11177] = 12'hfff;
rom[11178] = 12'hfff;
rom[11179] = 12'hfff;
rom[11180] = 12'hfff;
rom[11181] = 12'hfff;
rom[11182] = 12'hfff;
rom[11183] = 12'hfff;
rom[11184] = 12'hfff;
rom[11185] = 12'hfff;
rom[11186] = 12'hfff;
rom[11187] = 12'hfff;
rom[11188] = 12'hfff;
rom[11189] = 12'hfff;
rom[11190] = 12'hfff;
rom[11191] = 12'hfff;
rom[11192] = 12'hfff;
rom[11193] = 12'hfff;
rom[11194] = 12'h66e;
rom[11195] = 12'h  c;
rom[11196] = 12'h  c;
rom[11197] = 12'h  c;
rom[11198] = 12'h  c;
rom[11199] = 12'h99e;
rom[11200] = 12'hfff;
rom[11201] = 12'hfff;
rom[11202] = 12'hfff;
rom[11203] = 12'hfff;
rom[11204] = 12'hfff;
rom[11205] = 12'hfff;
rom[11206] = 12'hfff;
rom[11207] = 12'hfff;
rom[11208] = 12'hfff;
rom[11209] = 12'hfff;
rom[11210] = 12'hfff;
rom[11211] = 12'hfff;
rom[11212] = 12'hfff;
rom[11213] = 12'hfff;
rom[11214] = 12'hfff;
rom[11215] = 12'hfff;
rom[11216] = 12'hfff;
rom[11217] = 12'hfff;
rom[11218] = 12'hfff;
rom[11219] = 12'hfff;
rom[11220] = 12'hfff;
rom[11221] = 12'hfff;
rom[11222] = 12'hfff;
rom[11223] = 12'hfff;
rom[11224] = 12'hfff;
rom[11225] = 12'hfff;
rom[11226] = 12'hfff;
rom[11227] = 12'heef;
rom[11228] = 12'h11d;
rom[11229] = 12'h  c;
rom[11230] = 12'h  c;
rom[11231] = 12'h  c;
rom[11232] = 12'h  c;
rom[11233] = 12'h  c;
rom[11234] = 12'h88e;
rom[11235] = 12'hfff;
rom[11236] = 12'hfff;
rom[11237] = 12'hfff;
rom[11238] = 12'hfff;
rom[11239] = 12'hfff;
rom[11240] = 12'hfff;
rom[11241] = 12'hfff;
rom[11242] = 12'hfff;
rom[11243] = 12'hfff;
rom[11244] = 12'hfff;
rom[11245] = 12'hfff;
rom[11246] = 12'hfff;
rom[11247] = 12'hfff;
rom[11248] = 12'hfff;
rom[11249] = 12'hfff;
rom[11250] = 12'hfff;
rom[11251] = 12'hfff;
rom[11252] = 12'hfff;
rom[11253] = 12'hfff;
rom[11254] = 12'hfff;
rom[11255] = 12'hfff;
rom[11256] = 12'hfff;
rom[11257] = 12'hfff;
rom[11258] = 12'hfff;
rom[11259] = 12'hfff;
rom[11260] = 12'hfff;
rom[11261] = 12'hfff;
rom[11262] = 12'hfff;
rom[11263] = 12'hfff;
rom[11264] = 12'hfff;
rom[11265] = 12'hfff;
rom[11266] = 12'hfff;
rom[11267] = 12'hfff;
rom[11268] = 12'hfff;
rom[11269] = 12'hfff;
rom[11270] = 12'hfff;
rom[11271] = 12'hfff;
rom[11272] = 12'hfff;
rom[11273] = 12'hfff;
rom[11274] = 12'hfff;
rom[11275] = 12'hfff;
rom[11276] = 12'hfff;
rom[11277] = 12'hfff;
rom[11278] = 12'hfff;
rom[11279] = 12'hfff;
rom[11280] = 12'hfff;
rom[11281] = 12'hfff;
rom[11282] = 12'h  c;
rom[11283] = 12'h  c;
rom[11284] = 12'h  c;
rom[11285] = 12'h  c;
rom[11286] = 12'h  c;
rom[11287] = 12'hfff;
rom[11288] = 12'hfff;
rom[11289] = 12'hfff;
rom[11290] = 12'hfff;
rom[11291] = 12'hfff;
rom[11292] = 12'hfff;
rom[11293] = 12'hfff;
rom[11294] = 12'hfff;
rom[11295] = 12'hfff;
rom[11296] = 12'hfff;
rom[11297] = 12'hfff;
rom[11298] = 12'hfff;
rom[11299] = 12'hfff;
rom[11300] = 12'hfff;
rom[11301] = 12'hfff;
rom[11302] = 12'hfff;
rom[11303] = 12'hfff;
rom[11304] = 12'hfff;
rom[11305] = 12'hfff;
rom[11306] = 12'hfff;
rom[11307] = 12'hfff;
rom[11308] = 12'hfff;
rom[11309] = 12'hfff;
rom[11310] = 12'hfff;
rom[11311] = 12'hfff;
rom[11312] = 12'hfff;
rom[11313] = 12'hfff;
rom[11314] = 12'hfff;
rom[11315] = 12'hfff;
rom[11316] = 12'hfff;
rom[11317] = 12'hfff;
rom[11318] = 12'hfff;
rom[11319] = 12'hfff;
rom[11320] = 12'hfff;
rom[11321] = 12'hfff;
rom[11322] = 12'h55d;
rom[11323] = 12'h  c;
rom[11324] = 12'h  c;
rom[11325] = 12'h  c;
rom[11326] = 12'h  c;
rom[11327] = 12'haae;
rom[11328] = 12'hfff;
rom[11329] = 12'hfff;
rom[11330] = 12'hfff;
rom[11331] = 12'hfff;
rom[11332] = 12'hfff;
rom[11333] = 12'hfff;
rom[11334] = 12'hfff;
rom[11335] = 12'hfff;
rom[11336] = 12'hfff;
rom[11337] = 12'hfff;
rom[11338] = 12'hfff;
rom[11339] = 12'hfff;
rom[11340] = 12'hfff;
rom[11341] = 12'hfff;
rom[11342] = 12'hfff;
rom[11343] = 12'hfff;
rom[11344] = 12'hfff;
rom[11345] = 12'hfff;
rom[11346] = 12'hfff;
rom[11347] = 12'hfff;
rom[11348] = 12'hfff;
rom[11349] = 12'hfff;
rom[11350] = 12'hfff;
rom[11351] = 12'hfff;
rom[11352] = 12'hfff;
rom[11353] = 12'hfff;
rom[11354] = 12'hfff;
rom[11355] = 12'hfff;
rom[11356] = 12'hddf;
rom[11357] = 12'h11d;
rom[11358] = 12'h  c;
rom[11359] = 12'h  c;
rom[11360] = 12'h  c;
rom[11361] = 12'h  c;
rom[11362] = 12'h  c;
rom[11363] = 12'heef;
rom[11364] = 12'hfff;
rom[11365] = 12'hfff;
rom[11366] = 12'hfff;
rom[11367] = 12'hfff;
rom[11368] = 12'hfff;
rom[11369] = 12'hfff;
rom[11370] = 12'hfff;
rom[11371] = 12'hfff;
rom[11372] = 12'hfff;
rom[11373] = 12'hfff;
rom[11374] = 12'hfff;
rom[11375] = 12'hfff;
rom[11376] = 12'hfff;
rom[11377] = 12'hfff;
rom[11378] = 12'hfff;
rom[11379] = 12'hfff;
rom[11380] = 12'hfff;
rom[11381] = 12'hfff;
rom[11382] = 12'hfff;
rom[11383] = 12'hfff;
rom[11384] = 12'hfff;
rom[11385] = 12'hfff;
rom[11386] = 12'hfff;
rom[11387] = 12'hfff;
rom[11388] = 12'hfff;
rom[11389] = 12'hfff;
rom[11390] = 12'hfff;
rom[11391] = 12'hfff;
rom[11392] = 12'hfff;
rom[11393] = 12'hfff;
rom[11394] = 12'hfff;
rom[11395] = 12'hfff;
rom[11396] = 12'hfff;
rom[11397] = 12'hfff;
rom[11398] = 12'hfff;
rom[11399] = 12'hfff;
rom[11400] = 12'hfff;
rom[11401] = 12'hfff;
rom[11402] = 12'hfff;
rom[11403] = 12'hfff;
rom[11404] = 12'hfff;
rom[11405] = 12'hfff;
rom[11406] = 12'hfff;
rom[11407] = 12'hfff;
rom[11408] = 12'hfff;
rom[11409] = 12'heef;
rom[11410] = 12'h  c;
rom[11411] = 12'h  c;
rom[11412] = 12'h  c;
rom[11413] = 12'h  c;
rom[11414] = 12'h11d;
rom[11415] = 12'hfff;
rom[11416] = 12'hfff;
rom[11417] = 12'hfff;
rom[11418] = 12'hfff;
rom[11419] = 12'hfff;
rom[11420] = 12'hfff;
rom[11421] = 12'hfff;
rom[11422] = 12'hfff;
rom[11423] = 12'hfff;
rom[11424] = 12'hfff;
rom[11425] = 12'hfff;
rom[11426] = 12'hfff;
rom[11427] = 12'hfff;
rom[11428] = 12'hfff;
rom[11429] = 12'hfff;
rom[11430] = 12'hfff;
rom[11431] = 12'hfff;
rom[11432] = 12'hfff;
rom[11433] = 12'hfff;
rom[11434] = 12'hfff;
rom[11435] = 12'hfff;
rom[11436] = 12'hfff;
rom[11437] = 12'hfff;
rom[11438] = 12'hfff;
rom[11439] = 12'hfff;
rom[11440] = 12'hfff;
rom[11441] = 12'hfff;
rom[11442] = 12'hfff;
rom[11443] = 12'hfff;
rom[11444] = 12'hfff;
rom[11445] = 12'hfff;
rom[11446] = 12'hfff;
rom[11447] = 12'hfff;
rom[11448] = 12'hfff;
rom[11449] = 12'hfff;
rom[11450] = 12'h44d;
rom[11451] = 12'h  c;
rom[11452] = 12'h  c;
rom[11453] = 12'h  c;
rom[11454] = 12'h  c;
rom[11455] = 12'hbbe;
rom[11456] = 12'hfff;
rom[11457] = 12'hfff;
rom[11458] = 12'hfff;
rom[11459] = 12'hfff;
rom[11460] = 12'hfff;
rom[11461] = 12'hfff;
rom[11462] = 12'hfff;
rom[11463] = 12'hfff;
rom[11464] = 12'hfff;
rom[11465] = 12'hfff;
rom[11466] = 12'hfff;
rom[11467] = 12'hfff;
rom[11468] = 12'hfff;
rom[11469] = 12'hfff;
rom[11470] = 12'hfff;
rom[11471] = 12'hfff;
rom[11472] = 12'hfff;
rom[11473] = 12'hfff;
rom[11474] = 12'hfff;
rom[11475] = 12'hfff;
rom[11476] = 12'hfff;
rom[11477] = 12'hfff;
rom[11478] = 12'hfff;
rom[11479] = 12'hfff;
rom[11480] = 12'hfff;
rom[11481] = 12'hfff;
rom[11482] = 12'hfff;
rom[11483] = 12'hfff;
rom[11484] = 12'hfff;
rom[11485] = 12'heef;
rom[11486] = 12'h11d;
rom[11487] = 12'h  c;
rom[11488] = 12'h  c;
rom[11489] = 12'h  c;
rom[11490] = 12'h  c;
rom[11491] = 12'h88e;
rom[11492] = 12'hfff;
rom[11493] = 12'hfff;
rom[11494] = 12'hfff;
rom[11495] = 12'hfff;
rom[11496] = 12'hfff;
rom[11497] = 12'hfff;
rom[11498] = 12'hfff;
rom[11499] = 12'hfff;
rom[11500] = 12'hfff;
rom[11501] = 12'hfff;
rom[11502] = 12'hfff;
rom[11503] = 12'hfff;
rom[11504] = 12'hfff;
rom[11505] = 12'hfff;
rom[11506] = 12'hfff;
rom[11507] = 12'hfff;
rom[11508] = 12'hfff;
rom[11509] = 12'hfff;
rom[11510] = 12'hfff;
rom[11511] = 12'hfff;
rom[11512] = 12'hfff;
rom[11513] = 12'hfff;
rom[11514] = 12'hfff;
rom[11515] = 12'hfff;
rom[11516] = 12'hfff;
rom[11517] = 12'hfff;
rom[11518] = 12'hfff;
rom[11519] = 12'hfff;
rom[11520] = 12'hfff;
rom[11521] = 12'hfff;
rom[11522] = 12'hfff;
rom[11523] = 12'hfff;
rom[11524] = 12'hfff;
rom[11525] = 12'hfff;
rom[11526] = 12'hfff;
rom[11527] = 12'hfff;
rom[11528] = 12'hfff;
rom[11529] = 12'hfff;
rom[11530] = 12'hfff;
rom[11531] = 12'hfff;
rom[11532] = 12'hfff;
rom[11533] = 12'hfff;
rom[11534] = 12'hfff;
rom[11535] = 12'hfff;
rom[11536] = 12'hfff;
rom[11537] = 12'heef;
rom[11538] = 12'h  c;
rom[11539] = 12'h  c;
rom[11540] = 12'h  c;
rom[11541] = 12'h  c;
rom[11542] = 12'h11d;
rom[11543] = 12'hfff;
rom[11544] = 12'hfff;
rom[11545] = 12'hfff;
rom[11546] = 12'hfff;
rom[11547] = 12'hfff;
rom[11548] = 12'hfff;
rom[11549] = 12'hfff;
rom[11550] = 12'hfff;
rom[11551] = 12'hfff;
rom[11552] = 12'hfff;
rom[11553] = 12'hfff;
rom[11554] = 12'hfff;
rom[11555] = 12'hfff;
rom[11556] = 12'hfff;
rom[11557] = 12'hfff;
rom[11558] = 12'hfff;
rom[11559] = 12'hfff;
rom[11560] = 12'hfff;
rom[11561] = 12'hfff;
rom[11562] = 12'hfff;
rom[11563] = 12'hfff;
rom[11564] = 12'hfff;
rom[11565] = 12'hfff;
rom[11566] = 12'hfff;
rom[11567] = 12'hfff;
rom[11568] = 12'hfff;
rom[11569] = 12'hfff;
rom[11570] = 12'hfff;
rom[11571] = 12'hfff;
rom[11572] = 12'hfff;
rom[11573] = 12'hfff;
rom[11574] = 12'hfff;
rom[11575] = 12'hfff;
rom[11576] = 12'hfff;
rom[11577] = 12'hfff;
rom[11578] = 12'h44d;
rom[11579] = 12'h  c;
rom[11580] = 12'h  c;
rom[11581] = 12'h  c;
rom[11582] = 12'h  c;
rom[11583] = 12'hbbf;
rom[11584] = 12'hfff;
rom[11585] = 12'hfff;
rom[11586] = 12'hfff;
rom[11587] = 12'hfff;
rom[11588] = 12'hfff;
rom[11589] = 12'hfff;
rom[11590] = 12'hfff;
rom[11591] = 12'hfff;
rom[11592] = 12'hfff;
rom[11593] = 12'hfff;
rom[11594] = 12'hfff;
rom[11595] = 12'hfff;
rom[11596] = 12'hfff;
rom[11597] = 12'hfff;
rom[11598] = 12'hfff;
rom[11599] = 12'hfff;
rom[11600] = 12'hfff;
rom[11601] = 12'hfff;
rom[11602] = 12'hfff;
rom[11603] = 12'hfff;
rom[11604] = 12'hfff;
rom[11605] = 12'hfff;
rom[11606] = 12'hfff;
rom[11607] = 12'hfff;
rom[11608] = 12'hfff;
rom[11609] = 12'hfff;
rom[11610] = 12'hfff;
rom[11611] = 12'hfff;
rom[11612] = 12'hfff;
rom[11613] = 12'hfff;
rom[11614] = 12'h88e;
rom[11615] = 12'h  c;
rom[11616] = 12'h  c;
rom[11617] = 12'h  c;
rom[11618] = 12'h  c;
rom[11619] = 12'h11d;
rom[11620] = 12'heef;
rom[11621] = 12'hfff;
rom[11622] = 12'hfff;
rom[11623] = 12'hfff;
rom[11624] = 12'hfff;
rom[11625] = 12'hfff;
rom[11626] = 12'hfff;
rom[11627] = 12'hfff;
rom[11628] = 12'hfff;
rom[11629] = 12'hfff;
rom[11630] = 12'hfff;
rom[11631] = 12'hfff;
rom[11632] = 12'hfff;
rom[11633] = 12'hfff;
rom[11634] = 12'hfff;
rom[11635] = 12'hfff;
rom[11636] = 12'hfff;
rom[11637] = 12'hfff;
rom[11638] = 12'hfff;
rom[11639] = 12'hfff;
rom[11640] = 12'hfff;
rom[11641] = 12'hfff;
rom[11642] = 12'hfff;
rom[11643] = 12'hfff;
rom[11644] = 12'hfff;
rom[11645] = 12'hfff;
rom[11646] = 12'hfff;
rom[11647] = 12'hfff;
rom[11648] = 12'hfff;
rom[11649] = 12'hfff;
rom[11650] = 12'hfff;
rom[11651] = 12'hfff;
rom[11652] = 12'hfff;
rom[11653] = 12'hfff;
rom[11654] = 12'hfff;
rom[11655] = 12'hfff;
rom[11656] = 12'hfff;
rom[11657] = 12'hfff;
rom[11658] = 12'hfff;
rom[11659] = 12'hfff;
rom[11660] = 12'hfff;
rom[11661] = 12'hfff;
rom[11662] = 12'hfff;
rom[11663] = 12'hfff;
rom[11664] = 12'hfff;
rom[11665] = 12'heef;
rom[11666] = 12'h  c;
rom[11667] = 12'h  c;
rom[11668] = 12'h  c;
rom[11669] = 12'h  c;
rom[11670] = 12'h11d;
rom[11671] = 12'hfff;
rom[11672] = 12'hfff;
rom[11673] = 12'hfff;
rom[11674] = 12'hfff;
rom[11675] = 12'hfff;
rom[11676] = 12'hfff;
rom[11677] = 12'hfff;
rom[11678] = 12'hfff;
rom[11679] = 12'hfff;
rom[11680] = 12'hfff;
rom[11681] = 12'hfff;
rom[11682] = 12'hfff;
rom[11683] = 12'hfff;
rom[11684] = 12'hfff;
rom[11685] = 12'hfff;
rom[11686] = 12'hfff;
rom[11687] = 12'hfff;
rom[11688] = 12'hfff;
rom[11689] = 12'hfff;
rom[11690] = 12'hfff;
rom[11691] = 12'hfff;
rom[11692] = 12'hfff;
rom[11693] = 12'hfff;
rom[11694] = 12'hfff;
rom[11695] = 12'hfff;
rom[11696] = 12'hfff;
rom[11697] = 12'hfff;
rom[11698] = 12'hfff;
rom[11699] = 12'hfff;
rom[11700] = 12'hfff;
rom[11701] = 12'hfff;
rom[11702] = 12'hfff;
rom[11703] = 12'hfff;
rom[11704] = 12'hfff;
rom[11705] = 12'hfff;
rom[11706] = 12'h33d;
rom[11707] = 12'h  c;
rom[11708] = 12'h  c;
rom[11709] = 12'h  c;
rom[11710] = 12'h  c;
rom[11711] = 12'hccf;
rom[11712] = 12'hfff;
rom[11713] = 12'hfff;
rom[11714] = 12'hfff;
rom[11715] = 12'hfff;
rom[11716] = 12'hfff;
rom[11717] = 12'hfff;
rom[11718] = 12'hfff;
rom[11719] = 12'hfff;
rom[11720] = 12'hfff;
rom[11721] = 12'hfff;
rom[11722] = 12'hfff;
rom[11723] = 12'hfff;
rom[11724] = 12'hfff;
rom[11725] = 12'hfff;
rom[11726] = 12'hfff;
rom[11727] = 12'hfff;
rom[11728] = 12'hfff;
rom[11729] = 12'hfff;
rom[11730] = 12'hfff;
rom[11731] = 12'hfff;
rom[11732] = 12'hfff;
rom[11733] = 12'hfff;
rom[11734] = 12'hfff;
rom[11735] = 12'hfff;
rom[11736] = 12'hfff;
rom[11737] = 12'hfff;
rom[11738] = 12'hfff;
rom[11739] = 12'hfff;
rom[11740] = 12'hfff;
rom[11741] = 12'hfff;
rom[11742] = 12'heef;
rom[11743] = 12'h  c;
rom[11744] = 12'h  c;
rom[11745] = 12'h  c;
rom[11746] = 12'h  c;
rom[11747] = 12'h  c;
rom[11748] = 12'h33d;
rom[11749] = 12'hfff;
rom[11750] = 12'hfff;
rom[11751] = 12'hfff;
rom[11752] = 12'hfff;
rom[11753] = 12'hfff;
rom[11754] = 12'hfff;
rom[11755] = 12'hfff;
rom[11756] = 12'hfff;
rom[11757] = 12'hfff;
rom[11758] = 12'hfff;
rom[11759] = 12'hfff;
rom[11760] = 12'hfff;
rom[11761] = 12'hfff;
rom[11762] = 12'hfff;
rom[11763] = 12'hfff;
rom[11764] = 12'hfff;
rom[11765] = 12'hfff;
rom[11766] = 12'hfff;
rom[11767] = 12'hfff;
rom[11768] = 12'hfff;
rom[11769] = 12'hfff;
rom[11770] = 12'hfff;
rom[11771] = 12'hfff;
rom[11772] = 12'hfff;
rom[11773] = 12'hfff;
rom[11774] = 12'hfff;
rom[11775] = 12'hfff;
rom[11776] = 12'hfff;
rom[11777] = 12'hfff;
rom[11778] = 12'hfff;
rom[11779] = 12'hfff;
rom[11780] = 12'hfff;
rom[11781] = 12'hfff;
rom[11782] = 12'hfff;
rom[11783] = 12'hfff;
rom[11784] = 12'hfff;
rom[11785] = 12'hfff;
rom[11786] = 12'hfff;
rom[11787] = 12'hfff;
rom[11788] = 12'hfff;
rom[11789] = 12'hfff;
rom[11790] = 12'hfff;
rom[11791] = 12'hfff;
rom[11792] = 12'hfff;
rom[11793] = 12'heef;
rom[11794] = 12'h  c;
rom[11795] = 12'h  c;
rom[11796] = 12'h  c;
rom[11797] = 12'h  c;
rom[11798] = 12'h11d;
rom[11799] = 12'hfff;
rom[11800] = 12'hfff;
rom[11801] = 12'hfff;
rom[11802] = 12'hfff;
rom[11803] = 12'hfff;
rom[11804] = 12'hfff;
rom[11805] = 12'hfff;
rom[11806] = 12'hfff;
rom[11807] = 12'hfff;
rom[11808] = 12'hfff;
rom[11809] = 12'hfff;
rom[11810] = 12'hfff;
rom[11811] = 12'hfff;
rom[11812] = 12'hfff;
rom[11813] = 12'hfff;
rom[11814] = 12'hfff;
rom[11815] = 12'hfff;
rom[11816] = 12'hfff;
rom[11817] = 12'hfff;
rom[11818] = 12'hfff;
rom[11819] = 12'hfff;
rom[11820] = 12'hfff;
rom[11821] = 12'hfff;
rom[11822] = 12'hfff;
rom[11823] = 12'hfff;
rom[11824] = 12'hfff;
rom[11825] = 12'hfff;
rom[11826] = 12'hfff;
rom[11827] = 12'hfff;
rom[11828] = 12'hfff;
rom[11829] = 12'hfff;
rom[11830] = 12'hfff;
rom[11831] = 12'hfff;
rom[11832] = 12'hfff;
rom[11833] = 12'hfff;
rom[11834] = 12'h22d;
rom[11835] = 12'h  c;
rom[11836] = 12'h  c;
rom[11837] = 12'h  c;
rom[11838] = 12'h  c;
rom[11839] = 12'hddf;
rom[11840] = 12'hfff;
rom[11841] = 12'hfff;
rom[11842] = 12'hfff;
rom[11843] = 12'hfff;
rom[11844] = 12'hfff;
rom[11845] = 12'hfff;
rom[11846] = 12'hfff;
rom[11847] = 12'hfff;
rom[11848] = 12'hfff;
rom[11849] = 12'hfff;
rom[11850] = 12'hfff;
rom[11851] = 12'hfff;
rom[11852] = 12'hfff;
rom[11853] = 12'hfff;
rom[11854] = 12'hfff;
rom[11855] = 12'hfff;
rom[11856] = 12'hfff;
rom[11857] = 12'hfff;
rom[11858] = 12'hfff;
rom[11859] = 12'hfff;
rom[11860] = 12'hfff;
rom[11861] = 12'hfff;
rom[11862] = 12'hfff;
rom[11863] = 12'hfff;
rom[11864] = 12'hfff;
rom[11865] = 12'hfff;
rom[11866] = 12'hfff;
rom[11867] = 12'hfff;
rom[11868] = 12'hfff;
rom[11869] = 12'hfff;
rom[11870] = 12'hfff;
rom[11871] = 12'h88e;
rom[11872] = 12'h  c;
rom[11873] = 12'h  c;
rom[11874] = 12'h  c;
rom[11875] = 12'h  c;
rom[11876] = 12'h  c;
rom[11877] = 12'h22d;
rom[11878] = 12'hfff;
rom[11879] = 12'hfff;
rom[11880] = 12'hfff;
rom[11881] = 12'hfff;
rom[11882] = 12'hfff;
rom[11883] = 12'hfff;
rom[11884] = 12'hfff;
rom[11885] = 12'hfff;
rom[11886] = 12'hfff;
rom[11887] = 12'hfff;
rom[11888] = 12'hfff;
rom[11889] = 12'hfff;
rom[11890] = 12'hfff;
rom[11891] = 12'hfff;
rom[11892] = 12'hfff;
rom[11893] = 12'hfff;
rom[11894] = 12'hfff;
rom[11895] = 12'hfff;
rom[11896] = 12'hfff;
rom[11897] = 12'hfff;
rom[11898] = 12'hfff;
rom[11899] = 12'hfff;
rom[11900] = 12'hfff;
rom[11901] = 12'hfff;
rom[11902] = 12'hfff;
rom[11903] = 12'hfff;
rom[11904] = 12'hfff;
rom[11905] = 12'hfff;
rom[11906] = 12'hfff;
rom[11907] = 12'hfff;
rom[11908] = 12'hfff;
rom[11909] = 12'hfff;
rom[11910] = 12'hfff;
rom[11911] = 12'hfff;
rom[11912] = 12'hfff;
rom[11913] = 12'hfff;
rom[11914] = 12'hfff;
rom[11915] = 12'hfff;
rom[11916] = 12'hfff;
rom[11917] = 12'hfff;
rom[11918] = 12'hfff;
rom[11919] = 12'hfff;
rom[11920] = 12'hfff;
rom[11921] = 12'hfff;
rom[11922] = 12'h  c;
rom[11923] = 12'h  c;
rom[11924] = 12'h  c;
rom[11925] = 12'h  c;
rom[11926] = 12'h  c;
rom[11927] = 12'hfff;
rom[11928] = 12'hfff;
rom[11929] = 12'hfff;
rom[11930] = 12'hfff;
rom[11931] = 12'hfff;
rom[11932] = 12'hfff;
rom[11933] = 12'hfff;
rom[11934] = 12'hfff;
rom[11935] = 12'hfff;
rom[11936] = 12'hfff;
rom[11937] = 12'hfff;
rom[11938] = 12'hfff;
rom[11939] = 12'hfff;
rom[11940] = 12'hfff;
rom[11941] = 12'hfff;
rom[11942] = 12'hfff;
rom[11943] = 12'hfff;
rom[11944] = 12'hfff;
rom[11945] = 12'hfff;
rom[11946] = 12'hfff;
rom[11947] = 12'hfff;
rom[11948] = 12'hfff;
rom[11949] = 12'hfff;
rom[11950] = 12'hfff;
rom[11951] = 12'hfff;
rom[11952] = 12'hfff;
rom[11953] = 12'hfff;
rom[11954] = 12'hfff;
rom[11955] = 12'hfff;
rom[11956] = 12'hfff;
rom[11957] = 12'hfff;
rom[11958] = 12'hfff;
rom[11959] = 12'hfff;
rom[11960] = 12'hfff;
rom[11961] = 12'hfff;
rom[11962] = 12'h22d;
rom[11963] = 12'h  c;
rom[11964] = 12'h  c;
rom[11965] = 12'h  c;
rom[11966] = 12'h  c;
rom[11967] = 12'hddf;
rom[11968] = 12'hfff;
rom[11969] = 12'hfff;
rom[11970] = 12'hfff;
rom[11971] = 12'hfff;
rom[11972] = 12'hfff;
rom[11973] = 12'hfff;
rom[11974] = 12'hfff;
rom[11975] = 12'hfff;
rom[11976] = 12'hfff;
rom[11977] = 12'hfff;
rom[11978] = 12'hfff;
rom[11979] = 12'hfff;
rom[11980] = 12'hfff;
rom[11981] = 12'hfff;
rom[11982] = 12'hfff;
rom[11983] = 12'hfff;
rom[11984] = 12'hfff;
rom[11985] = 12'hfff;
rom[11986] = 12'hfff;
rom[11987] = 12'hfff;
rom[11988] = 12'hfff;
rom[11989] = 12'hfff;
rom[11990] = 12'hfff;
rom[11991] = 12'hfff;
rom[11992] = 12'hfff;
rom[11993] = 12'hfff;
rom[11994] = 12'hfff;
rom[11995] = 12'hfff;
rom[11996] = 12'hfff;
rom[11997] = 12'hfff;
rom[11998] = 12'hfff;
rom[11999] = 12'hfff;
rom[12000] = 12'h22d;
rom[12001] = 12'h  c;
rom[12002] = 12'h  c;
rom[12003] = 12'h  c;
rom[12004] = 12'h  c;
rom[12005] = 12'h  c;
rom[12006] = 12'h99e;
rom[12007] = 12'hfff;
rom[12008] = 12'hfff;
rom[12009] = 12'hfff;
rom[12010] = 12'hfff;
rom[12011] = 12'hfff;
rom[12012] = 12'hfff;
rom[12013] = 12'hfff;
rom[12014] = 12'hfff;
rom[12015] = 12'hfff;
rom[12016] = 12'hfff;
rom[12017] = 12'hfff;
rom[12018] = 12'hfff;
rom[12019] = 12'hfff;
rom[12020] = 12'hfff;
rom[12021] = 12'hfff;
rom[12022] = 12'hfff;
rom[12023] = 12'hfff;
rom[12024] = 12'hfff;
rom[12025] = 12'hfff;
rom[12026] = 12'hfff;
rom[12027] = 12'hfff;
rom[12028] = 12'hfff;
rom[12029] = 12'hfff;
rom[12030] = 12'hfff;
rom[12031] = 12'hfff;
rom[12032] = 12'hfff;
rom[12033] = 12'hfff;
rom[12034] = 12'hfff;
rom[12035] = 12'hfff;
rom[12036] = 12'hfff;
rom[12037] = 12'hfff;
rom[12038] = 12'hfff;
rom[12039] = 12'hfff;
rom[12040] = 12'hfff;
rom[12041] = 12'hfff;
rom[12042] = 12'hfff;
rom[12043] = 12'hfff;
rom[12044] = 12'hfff;
rom[12045] = 12'hfff;
rom[12046] = 12'hfff;
rom[12047] = 12'hfff;
rom[12048] = 12'hfff;
rom[12049] = 12'hfff;
rom[12050] = 12'h  c;
rom[12051] = 12'h  c;
rom[12052] = 12'h  c;
rom[12053] = 12'h  c;
rom[12054] = 12'h  c;
rom[12055] = 12'hfff;
rom[12056] = 12'hfff;
rom[12057] = 12'hfff;
rom[12058] = 12'hfff;
rom[12059] = 12'hfff;
rom[12060] = 12'hfff;
rom[12061] = 12'hfff;
rom[12062] = 12'hfff;
rom[12063] = 12'hfff;
rom[12064] = 12'hfff;
rom[12065] = 12'hfff;
rom[12066] = 12'hfff;
rom[12067] = 12'hfff;
rom[12068] = 12'hfff;
rom[12069] = 12'hfff;
rom[12070] = 12'hfff;
rom[12071] = 12'hfff;
rom[12072] = 12'hfff;
rom[12073] = 12'hfff;
rom[12074] = 12'hfff;
rom[12075] = 12'hfff;
rom[12076] = 12'hfff;
rom[12077] = 12'hfff;
rom[12078] = 12'hfff;
rom[12079] = 12'hfff;
rom[12080] = 12'hfff;
rom[12081] = 12'hfff;
rom[12082] = 12'hfff;
rom[12083] = 12'hfff;
rom[12084] = 12'hfff;
rom[12085] = 12'hfff;
rom[12086] = 12'hfff;
rom[12087] = 12'hfff;
rom[12088] = 12'hfff;
rom[12089] = 12'hfff;
rom[12090] = 12'h  c;
rom[12091] = 12'h  c;
rom[12092] = 12'h  c;
rom[12093] = 12'h  c;
rom[12094] = 12'h  c;
rom[12095] = 12'heef;
rom[12096] = 12'hfff;
rom[12097] = 12'hfff;
rom[12098] = 12'hfff;
rom[12099] = 12'hfff;
rom[12100] = 12'hfff;
rom[12101] = 12'hfff;
rom[12102] = 12'hfff;
rom[12103] = 12'hfff;
rom[12104] = 12'hfff;
rom[12105] = 12'hfff;
rom[12106] = 12'hfff;
rom[12107] = 12'hfff;
rom[12108] = 12'hfff;
rom[12109] = 12'hfff;
rom[12110] = 12'hfff;
rom[12111] = 12'hfff;
rom[12112] = 12'hfff;
rom[12113] = 12'hfff;
rom[12114] = 12'hfff;
rom[12115] = 12'hfff;
rom[12116] = 12'hfff;
rom[12117] = 12'hfff;
rom[12118] = 12'hfff;
rom[12119] = 12'hfff;
rom[12120] = 12'hfff;
rom[12121] = 12'hfff;
rom[12122] = 12'hfff;
rom[12123] = 12'hfff;
rom[12124] = 12'hfff;
rom[12125] = 12'hfff;
rom[12126] = 12'hfff;
rom[12127] = 12'hfff;
rom[12128] = 12'hfff;
rom[12129] = 12'h33d;
rom[12130] = 12'h  c;
rom[12131] = 12'h  c;
rom[12132] = 12'h  c;
rom[12133] = 12'h  c;
rom[12134] = 12'h22d;
rom[12135] = 12'hfff;
rom[12136] = 12'hfff;
rom[12137] = 12'hfff;
rom[12138] = 12'hfff;
rom[12139] = 12'hfff;
rom[12140] = 12'hfff;
rom[12141] = 12'hfff;
rom[12142] = 12'hfff;
rom[12143] = 12'hfff;
rom[12144] = 12'hfff;
rom[12145] = 12'hfff;
rom[12146] = 12'hfff;
rom[12147] = 12'hfff;
rom[12148] = 12'hfff;
rom[12149] = 12'hfff;
rom[12150] = 12'hfff;
rom[12151] = 12'hfff;
rom[12152] = 12'hfff;
rom[12153] = 12'hfff;
rom[12154] = 12'hfff;
rom[12155] = 12'hfff;
rom[12156] = 12'hfff;
rom[12157] = 12'hfff;
rom[12158] = 12'hfff;
rom[12159] = 12'hfff;
rom[12160] = 12'hfff;
rom[12161] = 12'hfff;
rom[12162] = 12'hfff;
rom[12163] = 12'hfff;
rom[12164] = 12'hfff;
rom[12165] = 12'hfff;
rom[12166] = 12'hfff;
rom[12167] = 12'hfff;
rom[12168] = 12'hfff;
rom[12169] = 12'hfff;
rom[12170] = 12'hfff;
rom[12171] = 12'hfff;
rom[12172] = 12'hfff;
rom[12173] = 12'hfff;
rom[12174] = 12'hfff;
rom[12175] = 12'hfff;
rom[12176] = 12'hfff;
rom[12177] = 12'hfff;
rom[12178] = 12'h11d;
rom[12179] = 12'h  c;
rom[12180] = 12'h  c;
rom[12181] = 12'h  c;
rom[12182] = 12'h  c;
rom[12183] = 12'hddf;
rom[12184] = 12'hfff;
rom[12185] = 12'hfff;
rom[12186] = 12'hfff;
rom[12187] = 12'hfff;
rom[12188] = 12'hfff;
rom[12189] = 12'hfff;
rom[12190] = 12'hfff;
rom[12191] = 12'hfff;
rom[12192] = 12'hfff;
rom[12193] = 12'hfff;
rom[12194] = 12'hfff;
rom[12195] = 12'hfff;
rom[12196] = 12'hfff;
rom[12197] = 12'hfff;
rom[12198] = 12'hfff;
rom[12199] = 12'hfff;
rom[12200] = 12'hfff;
rom[12201] = 12'hfff;
rom[12202] = 12'hfff;
rom[12203] = 12'hfff;
rom[12204] = 12'hfff;
rom[12205] = 12'hfff;
rom[12206] = 12'hfff;
rom[12207] = 12'hfff;
rom[12208] = 12'hfff;
rom[12209] = 12'hfff;
rom[12210] = 12'hfff;
rom[12211] = 12'hfff;
rom[12212] = 12'hfff;
rom[12213] = 12'hfff;
rom[12214] = 12'hfff;
rom[12215] = 12'hfff;
rom[12216] = 12'hfff;
rom[12217] = 12'heef;
rom[12218] = 12'h  c;
rom[12219] = 12'h  c;
rom[12220] = 12'h  c;
rom[12221] = 12'h  c;
rom[12222] = 12'h  c;
rom[12223] = 12'hfff;
rom[12224] = 12'hfff;
rom[12225] = 12'hfff;
rom[12226] = 12'hfff;
rom[12227] = 12'hfff;
rom[12228] = 12'hfff;
rom[12229] = 12'hfff;
rom[12230] = 12'hfff;
rom[12231] = 12'hfff;
rom[12232] = 12'hfff;
rom[12233] = 12'hfff;
rom[12234] = 12'hfff;
rom[12235] = 12'hfff;
rom[12236] = 12'hfff;
rom[12237] = 12'hfff;
rom[12238] = 12'hfff;
rom[12239] = 12'hfff;
rom[12240] = 12'hfff;
rom[12241] = 12'hfff;
rom[12242] = 12'hfff;
rom[12243] = 12'hfff;
rom[12244] = 12'hfff;
rom[12245] = 12'hfff;
rom[12246] = 12'hfff;
rom[12247] = 12'hfff;
rom[12248] = 12'hfff;
rom[12249] = 12'hfff;
rom[12250] = 12'hfff;
rom[12251] = 12'hfff;
rom[12252] = 12'hfff;
rom[12253] = 12'hfff;
rom[12254] = 12'hfff;
rom[12255] = 12'hfff;
rom[12256] = 12'hfff;
rom[12257] = 12'heef;
rom[12258] = 12'h11d;
rom[12259] = 12'h  c;
rom[12260] = 12'h  c;
rom[12261] = 12'h  c;
rom[12262] = 12'h  c;
rom[12263] = 12'hbbf;
rom[12264] = 12'hfff;
rom[12265] = 12'hfff;
rom[12266] = 12'hfff;
rom[12267] = 12'hfff;
rom[12268] = 12'hfff;
rom[12269] = 12'hfff;
rom[12270] = 12'hfff;
rom[12271] = 12'hfff;
rom[12272] = 12'hfff;
rom[12273] = 12'hfff;
rom[12274] = 12'hfff;
rom[12275] = 12'hfff;
rom[12276] = 12'hfff;
rom[12277] = 12'hfff;
rom[12278] = 12'hfff;
rom[12279] = 12'hfff;
rom[12280] = 12'hfff;
rom[12281] = 12'hfff;
rom[12282] = 12'hfff;
rom[12283] = 12'hfff;
rom[12284] = 12'hfff;
rom[12285] = 12'hfff;
rom[12286] = 12'hfff;
rom[12287] = 12'hfff;
rom[12288] = 12'hfff;
rom[12289] = 12'hfff;
rom[12290] = 12'hfff;
rom[12291] = 12'hfff;
rom[12292] = 12'hfff;
rom[12293] = 12'hfff;
rom[12294] = 12'hfff;
rom[12295] = 12'hfff;
rom[12296] = 12'hfff;
rom[12297] = 12'hfff;
rom[12298] = 12'hfff;
rom[12299] = 12'hfff;
rom[12300] = 12'hfff;
rom[12301] = 12'hfff;
rom[12302] = 12'hfff;
rom[12303] = 12'hfff;
rom[12304] = 12'hfff;
rom[12305] = 12'hfff;
rom[12306] = 12'h33d;
rom[12307] = 12'h  c;
rom[12308] = 12'h  c;
rom[12309] = 12'h  c;
rom[12310] = 12'h  c;
rom[12311] = 12'h55d;
rom[12312] = 12'hfff;
rom[12313] = 12'hfff;
rom[12314] = 12'hfff;
rom[12315] = 12'hfff;
rom[12316] = 12'hfff;
rom[12317] = 12'hfff;
rom[12318] = 12'hfff;
rom[12319] = 12'hfff;
rom[12320] = 12'hfff;
rom[12321] = 12'hfff;
rom[12322] = 12'hfff;
rom[12323] = 12'hfff;
rom[12324] = 12'hfff;
rom[12325] = 12'hfff;
rom[12326] = 12'hfff;
rom[12327] = 12'hfff;
rom[12328] = 12'hfff;
rom[12329] = 12'hfff;
rom[12330] = 12'hfff;
rom[12331] = 12'hfff;
rom[12332] = 12'hfff;
rom[12333] = 12'hfff;
rom[12334] = 12'hfff;
rom[12335] = 12'hfff;
rom[12336] = 12'hfff;
rom[12337] = 12'hfff;
rom[12338] = 12'hfff;
rom[12339] = 12'hfff;
rom[12340] = 12'hfff;
rom[12341] = 12'hfff;
rom[12342] = 12'hfff;
rom[12343] = 12'hfff;
rom[12344] = 12'hfff;
rom[12345] = 12'hccf;
rom[12346] = 12'h  c;
rom[12347] = 12'h  c;
rom[12348] = 12'h  c;
rom[12349] = 12'h  c;
rom[12350] = 12'h22d;
rom[12351] = 12'hfff;
rom[12352] = 12'hfff;
rom[12353] = 12'hfff;
rom[12354] = 12'hfff;
rom[12355] = 12'hfff;
rom[12356] = 12'hfff;
rom[12357] = 12'hfff;
rom[12358] = 12'hfff;
rom[12359] = 12'hfff;
rom[12360] = 12'hfff;
rom[12361] = 12'hfff;
rom[12362] = 12'hfff;
rom[12363] = 12'hfff;
rom[12364] = 12'hfff;
rom[12365] = 12'hfff;
rom[12366] = 12'hfff;
rom[12367] = 12'hfff;
rom[12368] = 12'hfff;
rom[12369] = 12'hfff;
rom[12370] = 12'hfff;
rom[12371] = 12'hfff;
rom[12372] = 12'hfff;
rom[12373] = 12'hfff;
rom[12374] = 12'hfff;
rom[12375] = 12'hfff;
rom[12376] = 12'hfff;
rom[12377] = 12'hfff;
rom[12378] = 12'hfff;
rom[12379] = 12'hfff;
rom[12380] = 12'hfff;
rom[12381] = 12'hfff;
rom[12382] = 12'hfff;
rom[12383] = 12'hfff;
rom[12384] = 12'hfff;
rom[12385] = 12'hfff;
rom[12386] = 12'h99e;
rom[12387] = 12'h  c;
rom[12388] = 12'h  c;
rom[12389] = 12'h  c;
rom[12390] = 12'h  c;
rom[12391] = 12'h66e;
rom[12392] = 12'hfff;
rom[12393] = 12'hfff;
rom[12394] = 12'hfff;
rom[12395] = 12'hfff;
rom[12396] = 12'hfff;
rom[12397] = 12'hfff;
rom[12398] = 12'hfff;
rom[12399] = 12'hfff;
rom[12400] = 12'hfff;
rom[12401] = 12'hfff;
rom[12402] = 12'hfff;
rom[12403] = 12'hfff;
rom[12404] = 12'hfff;
rom[12405] = 12'hfff;
rom[12406] = 12'hfff;
rom[12407] = 12'hfff;
rom[12408] = 12'hfff;
rom[12409] = 12'hfff;
rom[12410] = 12'hfff;
rom[12411] = 12'hfff;
rom[12412] = 12'hfff;
rom[12413] = 12'hfff;
rom[12414] = 12'hfff;
rom[12415] = 12'hfff;
rom[12416] = 12'hfff;
rom[12417] = 12'hfff;
rom[12418] = 12'hfff;
rom[12419] = 12'hfff;
rom[12420] = 12'hfff;
rom[12421] = 12'hfff;
rom[12422] = 12'hfff;
rom[12423] = 12'hfff;
rom[12424] = 12'hfff;
rom[12425] = 12'hfff;
rom[12426] = 12'hfff;
rom[12427] = 12'hfff;
rom[12428] = 12'hfff;
rom[12429] = 12'hfff;
rom[12430] = 12'hfff;
rom[12431] = 12'hfff;
rom[12432] = 12'hfff;
rom[12433] = 12'hfff;
rom[12434] = 12'h88e;
rom[12435] = 12'h  c;
rom[12436] = 12'h  c;
rom[12437] = 12'h  c;
rom[12438] = 12'h  c;
rom[12439] = 12'h  c;
rom[12440] = 12'h44d;
rom[12441] = 12'h77e;
rom[12442] = 12'h66e;
rom[12443] = 12'h99e;
rom[12444] = 12'heef;
rom[12445] = 12'hfff;
rom[12446] = 12'hfff;
rom[12447] = 12'hfff;
rom[12448] = 12'hfff;
rom[12449] = 12'hfff;
rom[12450] = 12'hfff;
rom[12451] = 12'hfff;
rom[12452] = 12'hfff;
rom[12453] = 12'hfff;
rom[12454] = 12'hfff;
rom[12455] = 12'hfff;
rom[12456] = 12'hfff;
rom[12457] = 12'hfff;
rom[12458] = 12'hfff;
rom[12459] = 12'hfff;
rom[12460] = 12'hfff;
rom[12461] = 12'hfff;
rom[12462] = 12'hfff;
rom[12463] = 12'hfff;
rom[12464] = 12'hfff;
rom[12465] = 12'hfff;
rom[12466] = 12'hfff;
rom[12467] = 12'hfff;
rom[12468] = 12'hfff;
rom[12469] = 12'hfff;
rom[12470] = 12'hfff;
rom[12471] = 12'hfff;
rom[12472] = 12'hfff;
rom[12473] = 12'h99e;
rom[12474] = 12'h11d;
rom[12475] = 12'h  c;
rom[12476] = 12'h  c;
rom[12477] = 12'h  c;
rom[12478] = 12'h55d;
rom[12479] = 12'hfff;
rom[12480] = 12'hfff;
rom[12481] = 12'hfff;
rom[12482] = 12'hfff;
rom[12483] = 12'hfff;
rom[12484] = 12'hfff;
rom[12485] = 12'hfff;
rom[12486] = 12'hfff;
rom[12487] = 12'hfff;
rom[12488] = 12'hfff;
rom[12489] = 12'hfff;
rom[12490] = 12'hfff;
rom[12491] = 12'hfff;
rom[12492] = 12'hfff;
rom[12493] = 12'hfff;
rom[12494] = 12'hfff;
rom[12495] = 12'hfff;
rom[12496] = 12'hfff;
rom[12497] = 12'hfff;
rom[12498] = 12'hfff;
rom[12499] = 12'hfff;
rom[12500] = 12'hfff;
rom[12501] = 12'hfff;
rom[12502] = 12'hfff;
rom[12503] = 12'hfff;
rom[12504] = 12'hfff;
rom[12505] = 12'hfff;
rom[12506] = 12'hfff;
rom[12507] = 12'hfff;
rom[12508] = 12'hfff;
rom[12509] = 12'hfff;
rom[12510] = 12'hfff;
rom[12511] = 12'hfff;
rom[12512] = 12'hfff;
rom[12513] = 12'hfff;
rom[12514] = 12'hddf;
rom[12515] = 12'h  c;
rom[12516] = 12'h  c;
rom[12517] = 12'h  c;
rom[12518] = 12'h  c;
rom[12519] = 12'h  c;
rom[12520] = 12'h99e;
rom[12521] = 12'hfff;
rom[12522] = 12'hfff;
rom[12523] = 12'hfff;
rom[12524] = 12'hfff;
rom[12525] = 12'hfff;
rom[12526] = 12'hfff;
rom[12527] = 12'hfff;
rom[12528] = 12'hfff;
rom[12529] = 12'hfff;
rom[12530] = 12'hfff;
rom[12531] = 12'hfff;
rom[12532] = 12'hfff;
rom[12533] = 12'hfff;
rom[12534] = 12'hfff;
rom[12535] = 12'hfff;
rom[12536] = 12'hfff;
rom[12537] = 12'hfff;
rom[12538] = 12'hfff;
rom[12539] = 12'hfff;
rom[12540] = 12'hfff;
rom[12541] = 12'hfff;
rom[12542] = 12'hfff;
rom[12543] = 12'hfff;
rom[12544] = 12'hfff;
rom[12545] = 12'hfff;
rom[12546] = 12'hfff;
rom[12547] = 12'hfff;
rom[12548] = 12'hfff;
rom[12549] = 12'hfff;
rom[12550] = 12'hfff;
rom[12551] = 12'hfff;
rom[12552] = 12'hfff;
rom[12553] = 12'hfff;
rom[12554] = 12'hfff;
rom[12555] = 12'hfff;
rom[12556] = 12'hfff;
rom[12557] = 12'hfff;
rom[12558] = 12'hfff;
rom[12559] = 12'hfff;
rom[12560] = 12'hfff;
rom[12561] = 12'hfff;
rom[12562] = 12'heef;
rom[12563] = 12'h11d;
rom[12564] = 12'h  c;
rom[12565] = 12'h  c;
rom[12566] = 12'h  c;
rom[12567] = 12'h  c;
rom[12568] = 12'h  c;
rom[12569] = 12'h11c;
rom[12570] = 12'h  c;
rom[12571] = 12'h  c;
rom[12572] = 12'h11d;
rom[12573] = 12'h77e;
rom[12574] = 12'h77e;
rom[12575] = 12'hccf;
rom[12576] = 12'hfff;
rom[12577] = 12'hfff;
rom[12578] = 12'hfff;
rom[12579] = 12'hfff;
rom[12580] = 12'hfff;
rom[12581] = 12'hfff;
rom[12582] = 12'hfff;
rom[12583] = 12'hfff;
rom[12584] = 12'hfff;
rom[12585] = 12'hfff;
rom[12586] = 12'hfff;
rom[12587] = 12'hfff;
rom[12588] = 12'hfff;
rom[12589] = 12'hfff;
rom[12590] = 12'hfff;
rom[12591] = 12'hfff;
rom[12592] = 12'hfff;
rom[12593] = 12'hfff;
rom[12594] = 12'hfff;
rom[12595] = 12'hfff;
rom[12596] = 12'hfff;
rom[12597] = 12'hfff;
rom[12598] = 12'hfff;
rom[12599] = 12'hfff;
rom[12600] = 12'hccf;
rom[12601] = 12'h44d;
rom[12602] = 12'h11d;
rom[12603] = 12'h  c;
rom[12604] = 12'h  c;
rom[12605] = 12'h  c;
rom[12606] = 12'h99e;
rom[12607] = 12'hfff;
rom[12608] = 12'hfff;
rom[12609] = 12'hfff;
rom[12610] = 12'hfff;
rom[12611] = 12'hfff;
rom[12612] = 12'hfff;
rom[12613] = 12'hfff;
rom[12614] = 12'hfff;
rom[12615] = 12'hfff;
rom[12616] = 12'hfff;
rom[12617] = 12'hfff;
rom[12618] = 12'hfff;
rom[12619] = 12'hfff;
rom[12620] = 12'hfff;
rom[12621] = 12'hfff;
rom[12622] = 12'hfff;
rom[12623] = 12'hfff;
rom[12624] = 12'hfff;
rom[12625] = 12'hfff;
rom[12626] = 12'hfff;
rom[12627] = 12'hfff;
rom[12628] = 12'hfff;
rom[12629] = 12'hfff;
rom[12630] = 12'hfff;
rom[12631] = 12'hfff;
rom[12632] = 12'hfff;
rom[12633] = 12'hfff;
rom[12634] = 12'hfff;
rom[12635] = 12'hfff;
rom[12636] = 12'hfff;
rom[12637] = 12'hfff;
rom[12638] = 12'hfff;
rom[12639] = 12'hfff;
rom[12640] = 12'hfff;
rom[12641] = 12'hfff;
rom[12642] = 12'hfff;
rom[12643] = 12'h44d;
rom[12644] = 12'h  c;
rom[12645] = 12'h  c;
rom[12646] = 12'h  c;
rom[12647] = 12'h  c;
rom[12648] = 12'h11d;
rom[12649] = 12'heef;
rom[12650] = 12'hfff;
rom[12651] = 12'hfff;
rom[12652] = 12'hfff;
rom[12653] = 12'hfff;
rom[12654] = 12'hfff;
rom[12655] = 12'hfff;
rom[12656] = 12'hfff;
rom[12657] = 12'hfff;
rom[12658] = 12'hfff;
rom[12659] = 12'hfff;
rom[12660] = 12'hfff;
rom[12661] = 12'hfff;
rom[12662] = 12'hfff;
rom[12663] = 12'hfff;
rom[12664] = 12'hfff;
rom[12665] = 12'hfff;
rom[12666] = 12'hfff;
rom[12667] = 12'hfff;
rom[12668] = 12'hfff;
rom[12669] = 12'hfff;
rom[12670] = 12'hfff;
rom[12671] = 12'hfff;
rom[12672] = 12'hfff;
rom[12673] = 12'hfff;
rom[12674] = 12'hfff;
rom[12675] = 12'hfff;
rom[12676] = 12'hfff;
rom[12677] = 12'hfff;
rom[12678] = 12'hfff;
rom[12679] = 12'hfff;
rom[12680] = 12'hfff;
rom[12681] = 12'hfff;
rom[12682] = 12'hfff;
rom[12683] = 12'hfff;
rom[12684] = 12'hfff;
rom[12685] = 12'hfff;
rom[12686] = 12'hfff;
rom[12687] = 12'hfff;
rom[12688] = 12'hfff;
rom[12689] = 12'hfff;
rom[12690] = 12'hfff;
rom[12691] = 12'hbbf;
rom[12692] = 12'h  c;
rom[12693] = 12'h  c;
rom[12694] = 12'h  c;
rom[12695] = 12'h  c;
rom[12696] = 12'h  c;
rom[12697] = 12'h  c;
rom[12698] = 12'h  c;
rom[12699] = 12'h  c;
rom[12700] = 12'h  c;
rom[12701] = 12'h  c;
rom[12702] = 12'h  c;
rom[12703] = 12'h  c;
rom[12704] = 12'h44d;
rom[12705] = 12'hbbf;
rom[12706] = 12'hddf;
rom[12707] = 12'hfff;
rom[12708] = 12'hfff;
rom[12709] = 12'hfff;
rom[12710] = 12'hfff;
rom[12711] = 12'hfff;
rom[12712] = 12'hfff;
rom[12713] = 12'hfff;
rom[12714] = 12'hfff;
rom[12715] = 12'hfff;
rom[12716] = 12'hfff;
rom[12717] = 12'hfff;
rom[12718] = 12'hfff;
rom[12719] = 12'hfff;
rom[12720] = 12'hfff;
rom[12721] = 12'hfff;
rom[12722] = 12'hfff;
rom[12723] = 12'hfff;
rom[12724] = 12'hfff;
rom[12725] = 12'hfff;
rom[12726] = 12'hddf;
rom[12727] = 12'h44d;
rom[12728] = 12'h  c;
rom[12729] = 12'h  c;
rom[12730] = 12'h  c;
rom[12731] = 12'h  c;
rom[12732] = 12'h  c;
rom[12733] = 12'h44d;
rom[12734] = 12'hfff;
rom[12735] = 12'hfff;
rom[12736] = 12'hfff;
rom[12737] = 12'hfff;
rom[12738] = 12'hfff;
rom[12739] = 12'hfff;
rom[12740] = 12'hfff;
rom[12741] = 12'hfff;
rom[12742] = 12'hfff;
rom[12743] = 12'hfff;
rom[12744] = 12'hfff;
rom[12745] = 12'hfff;
rom[12746] = 12'hfff;
rom[12747] = 12'hfff;
rom[12748] = 12'hfff;
rom[12749] = 12'hfff;
rom[12750] = 12'hfff;
rom[12751] = 12'hfff;
rom[12752] = 12'hfff;
rom[12753] = 12'hfff;
rom[12754] = 12'hfff;
rom[12755] = 12'hfff;
rom[12756] = 12'hfff;
rom[12757] = 12'hfff;
rom[12758] = 12'hfff;
rom[12759] = 12'hfff;
rom[12760] = 12'hfff;
rom[12761] = 12'hfff;
rom[12762] = 12'hfff;
rom[12763] = 12'hfff;
rom[12764] = 12'hfff;
rom[12765] = 12'hfff;
rom[12766] = 12'hfff;
rom[12767] = 12'hfff;
rom[12768] = 12'hfff;
rom[12769] = 12'hfff;
rom[12770] = 12'hfff;
rom[12771] = 12'haae;
rom[12772] = 12'h11d;
rom[12773] = 12'h  c;
rom[12774] = 12'h  c;
rom[12775] = 12'h  c;
rom[12776] = 12'h  c;
rom[12777] = 12'h99e;
rom[12778] = 12'hfff;
rom[12779] = 12'hfff;
rom[12780] = 12'hfff;
rom[12781] = 12'hfff;
rom[12782] = 12'hfff;
rom[12783] = 12'hfff;
rom[12784] = 12'hfff;
rom[12785] = 12'hfff;
rom[12786] = 12'hfff;
rom[12787] = 12'hfff;
rom[12788] = 12'hfff;
rom[12789] = 12'hfff;
rom[12790] = 12'hfff;
rom[12791] = 12'hfff;
rom[12792] = 12'hfff;
rom[12793] = 12'hfff;
rom[12794] = 12'hfff;
rom[12795] = 12'hfff;
rom[12796] = 12'hfff;
rom[12797] = 12'hfff;
rom[12798] = 12'hfff;
rom[12799] = 12'hfff;
rom[12800] = 12'hfff;
rom[12801] = 12'hfff;
rom[12802] = 12'hfff;
rom[12803] = 12'hfff;
rom[12804] = 12'hfff;
rom[12805] = 12'hfff;
rom[12806] = 12'hfff;
rom[12807] = 12'hfff;
rom[12808] = 12'hfff;
rom[12809] = 12'hfff;
rom[12810] = 12'hfff;
rom[12811] = 12'hfff;
rom[12812] = 12'hfff;
rom[12813] = 12'hfff;
rom[12814] = 12'hfff;
rom[12815] = 12'hfff;
rom[12816] = 12'hfff;
rom[12817] = 12'hfff;
rom[12818] = 12'hfff;
rom[12819] = 12'hfff;
rom[12820] = 12'haae;
rom[12821] = 12'h  c;
rom[12822] = 12'h  c;
rom[12823] = 12'h  c;
rom[12824] = 12'h  c;
rom[12825] = 12'h  c;
rom[12826] = 12'h  c;
rom[12827] = 12'h  c;
rom[12828] = 12'h  c;
rom[12829] = 12'h11d;
rom[12830] = 12'h  c;
rom[12831] = 12'h  c;
rom[12832] = 12'h  c;
rom[12833] = 12'h11d;
rom[12834] = 12'h  c;
rom[12835] = 12'h44d;
rom[12836] = 12'h77e;
rom[12837] = 12'h77e;
rom[12838] = 12'haae;
rom[12839] = 12'hfff;
rom[12840] = 12'hfff;
rom[12841] = 12'hfff;
rom[12842] = 12'hfff;
rom[12843] = 12'hfff;
rom[12844] = 12'hfff;
rom[12845] = 12'hfff;
rom[12846] = 12'hfff;
rom[12847] = 12'hfff;
rom[12848] = 12'hfff;
rom[12849] = 12'hfff;
rom[12850] = 12'hfff;
rom[12851] = 12'hfff;
rom[12852] = 12'hfff;
rom[12853] = 12'hccf;
rom[12854] = 12'h  c;
rom[12855] = 12'h  c;
rom[12856] = 12'h  c;
rom[12857] = 12'h  c;
rom[12858] = 12'h  c;
rom[12859] = 12'h  c;
rom[12860] = 12'h  c;
rom[12861] = 12'h99e;
rom[12862] = 12'hfff;
rom[12863] = 12'hfff;
rom[12864] = 12'hfff;
rom[12865] = 12'hfff;
rom[12866] = 12'hfff;
rom[12867] = 12'hfff;
rom[12868] = 12'hfff;
rom[12869] = 12'hfff;
rom[12870] = 12'hfff;
rom[12871] = 12'hfff;
rom[12872] = 12'hfff;
rom[12873] = 12'hfff;
rom[12874] = 12'hfff;
rom[12875] = 12'hfff;
rom[12876] = 12'hfff;
rom[12877] = 12'hfff;
rom[12878] = 12'hfff;
rom[12879] = 12'hfff;
rom[12880] = 12'hfff;
rom[12881] = 12'hfff;
rom[12882] = 12'hfff;
rom[12883] = 12'hfff;
rom[12884] = 12'hfff;
rom[12885] = 12'hfff;
rom[12886] = 12'hfff;
rom[12887] = 12'hfff;
rom[12888] = 12'hfff;
rom[12889] = 12'hfff;
rom[12890] = 12'hfff;
rom[12891] = 12'hfff;
rom[12892] = 12'hfff;
rom[12893] = 12'hfff;
rom[12894] = 12'hfff;
rom[12895] = 12'hfff;
rom[12896] = 12'hfff;
rom[12897] = 12'hfff;
rom[12898] = 12'hfff;
rom[12899] = 12'h99e;
rom[12900] = 12'h  c;
rom[12901] = 12'h  c;
rom[12902] = 12'h  c;
rom[12903] = 12'h  c;
rom[12904] = 12'h  c;
rom[12905] = 12'h66e;
rom[12906] = 12'hfff;
rom[12907] = 12'hfff;
rom[12908] = 12'hfff;
rom[12909] = 12'hfff;
rom[12910] = 12'hfff;
rom[12911] = 12'hfff;
rom[12912] = 12'hfff;
rom[12913] = 12'hfff;
rom[12914] = 12'hfff;
rom[12915] = 12'hfff;
rom[12916] = 12'hfff;
rom[12917] = 12'hfff;
rom[12918] = 12'hfff;
rom[12919] = 12'hfff;
rom[12920] = 12'hfff;
rom[12921] = 12'hfff;
rom[12922] = 12'hfff;
rom[12923] = 12'hfff;
rom[12924] = 12'hfff;
rom[12925] = 12'hfff;
rom[12926] = 12'hfff;
rom[12927] = 12'hfff;
rom[12928] = 12'hfff;
rom[12929] = 12'hfff;
rom[12930] = 12'hfff;
rom[12931] = 12'hfff;
rom[12932] = 12'hfff;
rom[12933] = 12'hfff;
rom[12934] = 12'hfff;
rom[12935] = 12'hfff;
rom[12936] = 12'hfff;
rom[12937] = 12'hfff;
rom[12938] = 12'hfff;
rom[12939] = 12'hfff;
rom[12940] = 12'hfff;
rom[12941] = 12'hfff;
rom[12942] = 12'hfff;
rom[12943] = 12'hfff;
rom[12944] = 12'hfff;
rom[12945] = 12'hfff;
rom[12946] = 12'hfff;
rom[12947] = 12'hfff;
rom[12948] = 12'hfff;
rom[12949] = 12'hbbf;
rom[12950] = 12'h11d;
rom[12951] = 12'h  c;
rom[12952] = 12'h  c;
rom[12953] = 12'h  c;
rom[12954] = 12'h  c;
rom[12955] = 12'h  c;
rom[12956] = 12'h  c;
rom[12957] = 12'h  c;
rom[12958] = 12'h  c;
rom[12959] = 12'h  c;
rom[12960] = 12'h  c;
rom[12961] = 12'h  c;
rom[12962] = 12'h  c;
rom[12963] = 12'h  c;
rom[12964] = 12'h11c;
rom[12965] = 12'h  c;
rom[12966] = 12'h  c;
rom[12967] = 12'h44d;
rom[12968] = 12'heef;
rom[12969] = 12'hfff;
rom[12970] = 12'hfff;
rom[12971] = 12'hfff;
rom[12972] = 12'hfff;
rom[12973] = 12'hfff;
rom[12974] = 12'hfff;
rom[12975] = 12'hfff;
rom[12976] = 12'hfff;
rom[12977] = 12'hfff;
rom[12978] = 12'hfff;
rom[12979] = 12'hfff;
rom[12980] = 12'heef;
rom[12981] = 12'h11d;
rom[12982] = 12'h11d;
rom[12983] = 12'h  c;
rom[12984] = 12'h  c;
rom[12985] = 12'h  c;
rom[12986] = 12'h  c;
rom[12987] = 12'h  c;
rom[12988] = 12'h22d;
rom[12989] = 12'heef;
rom[12990] = 12'hfff;
rom[12991] = 12'hfff;
rom[12992] = 12'hfff;
rom[12993] = 12'hfff;
rom[12994] = 12'hfff;
rom[12995] = 12'hfff;
rom[12996] = 12'hfff;
rom[12997] = 12'hfff;
rom[12998] = 12'hfff;
rom[12999] = 12'hfff;
rom[13000] = 12'hfff;
rom[13001] = 12'hfff;
rom[13002] = 12'hfff;
rom[13003] = 12'hfff;
rom[13004] = 12'hfff;
rom[13005] = 12'hfff;
rom[13006] = 12'hfff;
rom[13007] = 12'hfff;
rom[13008] = 12'hfff;
rom[13009] = 12'hfff;
rom[13010] = 12'hfff;
rom[13011] = 12'hfff;
rom[13012] = 12'hfff;
rom[13013] = 12'hfff;
rom[13014] = 12'hfff;
rom[13015] = 12'hfff;
rom[13016] = 12'hfff;
rom[13017] = 12'hfff;
rom[13018] = 12'hfff;
rom[13019] = 12'hfff;
rom[13020] = 12'hfff;
rom[13021] = 12'hfff;
rom[13022] = 12'hfff;
rom[13023] = 12'hfff;
rom[13024] = 12'hfff;
rom[13025] = 12'hfff;
rom[13026] = 12'hfff;
rom[13027] = 12'heef;
rom[13028] = 12'h11d;
rom[13029] = 12'h  c;
rom[13030] = 12'h  c;
rom[13031] = 12'h  c;
rom[13032] = 12'h  c;
rom[13033] = 12'h66e;
rom[13034] = 12'hfff;
rom[13035] = 12'hfff;
rom[13036] = 12'hfff;
rom[13037] = 12'hfff;
rom[13038] = 12'hfff;
rom[13039] = 12'hfff;
rom[13040] = 12'hfff;
rom[13041] = 12'hfff;
rom[13042] = 12'hfff;
rom[13043] = 12'hfff;
rom[13044] = 12'hfff;
rom[13045] = 12'hfff;
rom[13046] = 12'hfff;
rom[13047] = 12'hfff;
rom[13048] = 12'hfff;
rom[13049] = 12'hfff;
rom[13050] = 12'hfff;
rom[13051] = 12'hfff;
rom[13052] = 12'hfff;
rom[13053] = 12'hfff;
rom[13054] = 12'hfff;
rom[13055] = 12'hfff;
rom[13056] = 12'hfff;
rom[13057] = 12'hfff;
rom[13058] = 12'hfff;
rom[13059] = 12'hfff;
rom[13060] = 12'hfff;
rom[13061] = 12'hfff;
rom[13062] = 12'hfff;
rom[13063] = 12'hfff;
rom[13064] = 12'hfff;
rom[13065] = 12'hfff;
rom[13066] = 12'hfff;
rom[13067] = 12'hfff;
rom[13068] = 12'hfff;
rom[13069] = 12'hfff;
rom[13070] = 12'hfff;
rom[13071] = 12'hfff;
rom[13072] = 12'hfff;
rom[13073] = 12'hfff;
rom[13074] = 12'hfff;
rom[13075] = 12'hfff;
rom[13076] = 12'hfff;
rom[13077] = 12'hfff;
rom[13078] = 12'heef;
rom[13079] = 12'h99e;
rom[13080] = 12'h77e;
rom[13081] = 12'h11d;
rom[13082] = 12'h  c;
rom[13083] = 12'h  c;
rom[13084] = 12'h  c;
rom[13085] = 12'h  c;
rom[13086] = 12'h  c;
rom[13087] = 12'h  c;
rom[13088] = 12'h  c;
rom[13089] = 12'h  c;
rom[13090] = 12'h  c;
rom[13091] = 12'h  c;
rom[13092] = 12'h  c;
rom[13093] = 12'h  c;
rom[13094] = 12'h  c;
rom[13095] = 12'h  c;
rom[13096] = 12'h  c;
rom[13097] = 12'h11d;
rom[13098] = 12'h33d;
rom[13099] = 12'h44d;
rom[13100] = 12'h55d;
rom[13101] = 12'h66e;
rom[13102] = 12'h77e;
rom[13103] = 12'h88e;
rom[13104] = 12'h88e;
rom[13105] = 12'h88e;
rom[13106] = 12'h77e;
rom[13107] = 12'h66e;
rom[13108] = 12'h33d;
rom[13109] = 12'h  c;
rom[13110] = 12'h  c;
rom[13111] = 12'h  c;
rom[13112] = 12'h  c;
rom[13113] = 12'h22d;
rom[13114] = 12'h  c;
rom[13115] = 12'h11d;
rom[13116] = 12'heef;
rom[13117] = 12'hfff;
rom[13118] = 12'hfff;
rom[13119] = 12'hfff;
rom[13120] = 12'hfff;
rom[13121] = 12'hfff;
rom[13122] = 12'hfff;
rom[13123] = 12'hfff;
rom[13124] = 12'hfff;
rom[13125] = 12'hfff;
rom[13126] = 12'hfff;
rom[13127] = 12'hfff;
rom[13128] = 12'hfff;
rom[13129] = 12'hfff;
rom[13130] = 12'hfff;
rom[13131] = 12'hfff;
rom[13132] = 12'hfff;
rom[13133] = 12'hfff;
rom[13134] = 12'hfff;
rom[13135] = 12'hfff;
rom[13136] = 12'hfff;
rom[13137] = 12'hfff;
rom[13138] = 12'hfff;
rom[13139] = 12'hfff;
rom[13140] = 12'hfff;
rom[13141] = 12'hfff;
rom[13142] = 12'hfff;
rom[13143] = 12'hfff;
rom[13144] = 12'hfff;
rom[13145] = 12'hfff;
rom[13146] = 12'hfff;
rom[13147] = 12'hfff;
rom[13148] = 12'hfff;
rom[13149] = 12'hfff;
rom[13150] = 12'hfff;
rom[13151] = 12'hfff;
rom[13152] = 12'hfff;
rom[13153] = 12'hfff;
rom[13154] = 12'hfff;
rom[13155] = 12'hfff;
rom[13156] = 12'h88e;
rom[13157] = 12'h  c;
rom[13158] = 12'h11d;
rom[13159] = 12'h  c;
rom[13160] = 12'h  c;
rom[13161] = 12'h77e;
rom[13162] = 12'hfff;
rom[13163] = 12'hfff;
rom[13164] = 12'hfff;
rom[13165] = 12'hfff;
rom[13166] = 12'hfff;
rom[13167] = 12'hfff;
rom[13168] = 12'hfff;
rom[13169] = 12'hfff;
rom[13170] = 12'hfff;
rom[13171] = 12'hfff;
rom[13172] = 12'hfff;
rom[13173] = 12'hfff;
rom[13174] = 12'hfff;
rom[13175] = 12'hfff;
rom[13176] = 12'hfff;
rom[13177] = 12'hfff;
rom[13178] = 12'hfff;
rom[13179] = 12'hfff;
rom[13180] = 12'hfff;
rom[13181] = 12'hfff;
rom[13182] = 12'hfff;
rom[13183] = 12'hfff;
rom[13184] = 12'hfff;
rom[13185] = 12'hfff;
rom[13186] = 12'hfff;
rom[13187] = 12'hfff;
rom[13188] = 12'hfff;
rom[13189] = 12'hfff;
rom[13190] = 12'hfff;
rom[13191] = 12'hfff;
rom[13192] = 12'hfff;
rom[13193] = 12'hfff;
rom[13194] = 12'hfff;
rom[13195] = 12'hfff;
rom[13196] = 12'hfff;
rom[13197] = 12'hfff;
rom[13198] = 12'hfff;
rom[13199] = 12'hfff;
rom[13200] = 12'hfff;
rom[13201] = 12'hfff;
rom[13202] = 12'hfff;
rom[13203] = 12'hfff;
rom[13204] = 12'hfff;
rom[13205] = 12'hfff;
rom[13206] = 12'hfff;
rom[13207] = 12'hfff;
rom[13208] = 12'hfff;
rom[13209] = 12'heef;
rom[13210] = 12'h99e;
rom[13211] = 12'h66e;
rom[13212] = 12'h66e;
rom[13213] = 12'h77e;
rom[13214] = 12'h33d;
rom[13215] = 12'h  c;
rom[13216] = 12'h  c;
rom[13217] = 12'h  c;
rom[13218] = 12'h  c;
rom[13219] = 12'h  c;
rom[13220] = 12'h  c;
rom[13221] = 12'h  c;
rom[13222] = 12'h  c;
rom[13223] = 12'h  c;
rom[13224] = 12'h  c;
rom[13225] = 12'h  c;
rom[13226] = 12'h  c;
rom[13227] = 12'h  c;
rom[13228] = 12'h  c;
rom[13229] = 12'h  c;
rom[13230] = 12'h  c;
rom[13231] = 12'h  c;
rom[13232] = 12'h  c;
rom[13233] = 12'h  c;
rom[13234] = 12'h  c;
rom[13235] = 12'h  c;
rom[13236] = 12'h  c;
rom[13237] = 12'h  c;
rom[13238] = 12'h  c;
rom[13239] = 12'h  c;
rom[13240] = 12'h  c;
rom[13241] = 12'h55d;
rom[13242] = 12'h99e;
rom[13243] = 12'heef;
rom[13244] = 12'hfff;
rom[13245] = 12'hfff;
rom[13246] = 12'hfff;
rom[13247] = 12'hfff;
rom[13248] = 12'hfff;
rom[13249] = 12'hfff;
rom[13250] = 12'hfff;
rom[13251] = 12'hfff;
rom[13252] = 12'hfff;
rom[13253] = 12'hfff;
rom[13254] = 12'hfff;
rom[13255] = 12'hfff;
rom[13256] = 12'hfff;
rom[13257] = 12'hfff;
rom[13258] = 12'hfff;
rom[13259] = 12'hfff;
rom[13260] = 12'hfff;
rom[13261] = 12'hfff;
rom[13262] = 12'hfff;
rom[13263] = 12'hfff;
rom[13264] = 12'hfff;
rom[13265] = 12'hfff;
rom[13266] = 12'hfff;
rom[13267] = 12'hfff;
rom[13268] = 12'hfff;
rom[13269] = 12'hfff;
rom[13270] = 12'hfff;
rom[13271] = 12'hfff;
rom[13272] = 12'hfff;
rom[13273] = 12'hfff;
rom[13274] = 12'hfff;
rom[13275] = 12'hfff;
rom[13276] = 12'hfff;
rom[13277] = 12'hfff;
rom[13278] = 12'hfff;
rom[13279] = 12'hfff;
rom[13280] = 12'hfff;
rom[13281] = 12'hfff;
rom[13282] = 12'hfff;
rom[13283] = 12'hfff;
rom[13284] = 12'h99e;
rom[13285] = 12'h  c;
rom[13286] = 12'h  c;
rom[13287] = 12'h  c;
rom[13288] = 12'h  c;
rom[13289] = 12'h99e;
rom[13290] = 12'hfff;
rom[13291] = 12'hfff;
rom[13292] = 12'hfff;
rom[13293] = 12'hfff;
rom[13294] = 12'hfff;
rom[13295] = 12'hfff;
rom[13296] = 12'hfff;
rom[13297] = 12'hfff;
rom[13298] = 12'hfff;
rom[13299] = 12'hfff;
rom[13300] = 12'hfff;
rom[13301] = 12'hfff;
rom[13302] = 12'hfff;
rom[13303] = 12'hfff;
rom[13304] = 12'hfff;
rom[13305] = 12'hfff;
rom[13306] = 12'hfff;
rom[13307] = 12'hfff;
rom[13308] = 12'hfff;
rom[13309] = 12'hfff;
rom[13310] = 12'hfff;
rom[13311] = 12'hfff;
rom[13312] = 12'hfff;
rom[13313] = 12'hfff;
rom[13314] = 12'hfff;
rom[13315] = 12'hfff;
rom[13316] = 12'hfff;
rom[13317] = 12'hfff;
rom[13318] = 12'hfff;
rom[13319] = 12'hfff;
rom[13320] = 12'hfff;
rom[13321] = 12'hfff;
rom[13322] = 12'hfff;
rom[13323] = 12'hfff;
rom[13324] = 12'hfff;
rom[13325] = 12'hfff;
rom[13326] = 12'hfff;
rom[13327] = 12'hfff;
rom[13328] = 12'hfff;
rom[13329] = 12'hfff;
rom[13330] = 12'hfff;
rom[13331] = 12'hfff;
rom[13332] = 12'hfff;
rom[13333] = 12'hfff;
rom[13334] = 12'hfff;
rom[13335] = 12'hfff;
rom[13336] = 12'hfff;
rom[13337] = 12'hfff;
rom[13338] = 12'hfff;
rom[13339] = 12'hfff;
rom[13340] = 12'hfff;
rom[13341] = 12'hfff;
rom[13342] = 12'heef;
rom[13343] = 12'h99e;
rom[13344] = 12'h88e;
rom[13345] = 12'h33d;
rom[13346] = 12'h  c;
rom[13347] = 12'h  c;
rom[13348] = 12'h  c;
rom[13349] = 12'h  c;
rom[13350] = 12'h  c;
rom[13351] = 12'h  c;
rom[13352] = 12'h  c;
rom[13353] = 12'h  c;
rom[13354] = 12'h  c;
rom[13355] = 12'h  c;
rom[13356] = 12'h  c;
rom[13357] = 12'h  c;
rom[13358] = 12'h  c;
rom[13359] = 12'h  c;
rom[13360] = 12'h  c;
rom[13361] = 12'h  c;
rom[13362] = 12'h  c;
rom[13363] = 12'h  c;
rom[13364] = 12'h  c;
rom[13365] = 12'h  c;
rom[13366] = 12'h  c;
rom[13367] = 12'h  c;
rom[13368] = 12'h  c;
rom[13369] = 12'h99e;
rom[13370] = 12'hfff;
rom[13371] = 12'hfff;
rom[13372] = 12'hfff;
rom[13373] = 12'hfff;
rom[13374] = 12'hfff;
rom[13375] = 12'hfff;
rom[13376] = 12'hfff;
rom[13377] = 12'hfff;
rom[13378] = 12'hfff;
rom[13379] = 12'hfff;
rom[13380] = 12'hfff;
rom[13381] = 12'hfff;
rom[13382] = 12'hfff;
rom[13383] = 12'hfff;
rom[13384] = 12'hfff;
rom[13385] = 12'hfff;
rom[13386] = 12'hfff;
rom[13387] = 12'hfff;
rom[13388] = 12'hfff;
rom[13389] = 12'hfff;
rom[13390] = 12'hfff;
rom[13391] = 12'hfff;
rom[13392] = 12'hfff;
rom[13393] = 12'hfff;
rom[13394] = 12'hfff;
rom[13395] = 12'hfff;
rom[13396] = 12'hfff;
rom[13397] = 12'hfff;
rom[13398] = 12'hfff;
rom[13399] = 12'hfff;
rom[13400] = 12'hfff;
rom[13401] = 12'hfff;
rom[13402] = 12'hfff;
rom[13403] = 12'hfff;
rom[13404] = 12'hfff;
rom[13405] = 12'hfff;
rom[13406] = 12'hfff;
rom[13407] = 12'hfff;
rom[13408] = 12'hfff;
rom[13409] = 12'hfff;
rom[13410] = 12'hfff;
rom[13411] = 12'hfff;
rom[13412] = 12'heef;
rom[13413] = 12'h11d;
rom[13414] = 12'h  c;
rom[13415] = 12'h  c;
rom[13416] = 12'h11d;
rom[13417] = 12'heef;
rom[13418] = 12'hfff;
rom[13419] = 12'hfff;
rom[13420] = 12'hfff;
rom[13421] = 12'hfff;
rom[13422] = 12'hfff;
rom[13423] = 12'hfff;
rom[13424] = 12'hfff;
rom[13425] = 12'hfff;
rom[13426] = 12'hfff;
rom[13427] = 12'hfff;
rom[13428] = 12'hfff;
rom[13429] = 12'hfff;
rom[13430] = 12'hfff;
rom[13431] = 12'hfff;
rom[13432] = 12'hfff;
rom[13433] = 12'hfff;
rom[13434] = 12'hfff;
rom[13435] = 12'hfff;
rom[13436] = 12'hfff;
rom[13437] = 12'hfff;
rom[13438] = 12'hfff;
rom[13439] = 12'hfff;
rom[13440] = 12'hfff;
rom[13441] = 12'hfff;
rom[13442] = 12'hfff;
rom[13443] = 12'hfff;
rom[13444] = 12'hfff;
rom[13445] = 12'hfff;
rom[13446] = 12'hfff;
rom[13447] = 12'hfff;
rom[13448] = 12'hfff;
rom[13449] = 12'hfff;
rom[13450] = 12'hfff;
rom[13451] = 12'hfff;
rom[13452] = 12'hfff;
rom[13453] = 12'hfff;
rom[13454] = 12'hfff;
rom[13455] = 12'hfff;
rom[13456] = 12'hfff;
rom[13457] = 12'hfff;
rom[13458] = 12'hfff;
rom[13459] = 12'hfff;
rom[13460] = 12'hfff;
rom[13461] = 12'hfff;
rom[13462] = 12'hfff;
rom[13463] = 12'hfff;
rom[13464] = 12'hfff;
rom[13465] = 12'hfff;
rom[13466] = 12'hfff;
rom[13467] = 12'hfff;
rom[13468] = 12'hfff;
rom[13469] = 12'hfff;
rom[13470] = 12'hfff;
rom[13471] = 12'hfff;
rom[13472] = 12'hfff;
rom[13473] = 12'heef;
rom[13474] = 12'h99e;
rom[13475] = 12'h77e;
rom[13476] = 12'h88e;
rom[13477] = 12'h33d;
rom[13478] = 12'h  c;
rom[13479] = 12'h  c;
rom[13480] = 12'h  c;
rom[13481] = 12'h  c;
rom[13482] = 12'h  c;
rom[13483] = 12'h  c;
rom[13484] = 12'h  c;
rom[13485] = 12'h  c;
rom[13486] = 12'h  c;
rom[13487] = 12'h  c;
rom[13488] = 12'h  c;
rom[13489] = 12'h  c;
rom[13490] = 12'h  c;
rom[13491] = 12'h  c;
rom[13492] = 12'h  c;
rom[13493] = 12'h  c;
rom[13494] = 12'h  c;
rom[13495] = 12'h  c;
rom[13496] = 12'h11d;
rom[13497] = 12'heef;
rom[13498] = 12'hfff;
rom[13499] = 12'hfff;
rom[13500] = 12'hfff;
rom[13501] = 12'hfff;
rom[13502] = 12'hfff;
rom[13503] = 12'hfff;
rom[13504] = 12'hfff;
rom[13505] = 12'hfff;
rom[13506] = 12'hfff;
rom[13507] = 12'hfff;
rom[13508] = 12'hfff;
rom[13509] = 12'hfff;
rom[13510] = 12'hfff;
rom[13511] = 12'hfff;
rom[13512] = 12'hfff;
rom[13513] = 12'hfff;
rom[13514] = 12'hfff;
rom[13515] = 12'hfff;
rom[13516] = 12'hfff;
rom[13517] = 12'hfff;
rom[13518] = 12'hfff;
rom[13519] = 12'hfff;
rom[13520] = 12'hfff;
rom[13521] = 12'hfff;
rom[13522] = 12'hfff;
rom[13523] = 12'hfff;
rom[13524] = 12'hfff;
rom[13525] = 12'hfff;
rom[13526] = 12'hfff;
rom[13527] = 12'hfff;
rom[13528] = 12'hfff;
rom[13529] = 12'hfff;
rom[13530] = 12'hfff;
rom[13531] = 12'hfff;
rom[13532] = 12'hfff;
rom[13533] = 12'hfff;
rom[13534] = 12'hfff;
rom[13535] = 12'hfff;
rom[13536] = 12'hfff;
rom[13537] = 12'hfff;
rom[13538] = 12'hfff;
rom[13539] = 12'hfff;
rom[13540] = 12'hfff;
rom[13541] = 12'heef;
rom[13542] = 12'h99e;
rom[13543] = 12'h99e;
rom[13544] = 12'heef;
rom[13545] = 12'hfff;
rom[13546] = 12'hfff;
rom[13547] = 12'hfff;
rom[13548] = 12'hfff;
rom[13549] = 12'hfff;
rom[13550] = 12'hfff;
rom[13551] = 12'hfff;
rom[13552] = 12'hfff;
rom[13553] = 12'hfff;
rom[13554] = 12'hfff;
rom[13555] = 12'hfff;
rom[13556] = 12'hfff;
rom[13557] = 12'hfff;
rom[13558] = 12'hfff;
rom[13559] = 12'hfff;
rom[13560] = 12'hfff;
rom[13561] = 12'hfff;
rom[13562] = 12'hfff;
rom[13563] = 12'hfff;
rom[13564] = 12'hfff;
rom[13565] = 12'hfff;
rom[13566] = 12'hfff;
rom[13567] = 12'hfff;
rom[13568] = 12'hfff;
rom[13569] = 12'hfff;
rom[13570] = 12'hfff;
rom[13571] = 12'hfff;
rom[13572] = 12'hfff;
rom[13573] = 12'hfff;
rom[13574] = 12'hfff;
rom[13575] = 12'hfff;
rom[13576] = 12'hfff;
rom[13577] = 12'hfff;
rom[13578] = 12'hfff;
rom[13579] = 12'hfff;
rom[13580] = 12'hfff;
rom[13581] = 12'hfff;
rom[13582] = 12'hfff;
rom[13583] = 12'hfff;
rom[13584] = 12'hfff;
rom[13585] = 12'hfff;
rom[13586] = 12'hfff;
rom[13587] = 12'hfff;
rom[13588] = 12'hfff;
rom[13589] = 12'hfff;
rom[13590] = 12'hfff;
rom[13591] = 12'hfff;
rom[13592] = 12'hfff;
rom[13593] = 12'hfff;
rom[13594] = 12'hfff;
rom[13595] = 12'hfff;
rom[13596] = 12'hfff;
rom[13597] = 12'hfff;
rom[13598] = 12'hfff;
rom[13599] = 12'hfff;
rom[13600] = 12'hfff;
rom[13601] = 12'hfff;
rom[13602] = 12'hfff;
rom[13603] = 12'hfff;
rom[13604] = 12'hfff;
rom[13605] = 12'hfff;
rom[13606] = 12'haae;
rom[13607] = 12'h33d;
rom[13608] = 12'h  c;
rom[13609] = 12'h  c;
rom[13610] = 12'h  c;
rom[13611] = 12'h  c;
rom[13612] = 12'h  c;
rom[13613] = 12'h  c;
rom[13614] = 12'h  c;
rom[13615] = 12'h  c;
rom[13616] = 12'h  c;
rom[13617] = 12'h  c;
rom[13618] = 12'h  c;
rom[13619] = 12'h  c;
rom[13620] = 12'h  c;
rom[13621] = 12'h  c;
rom[13622] = 12'h  c;
rom[13623] = 12'h44d;
rom[13624] = 12'hddf;
rom[13625] = 12'hfff;
rom[13626] = 12'hfff;
rom[13627] = 12'hfff;
rom[13628] = 12'hfff;
rom[13629] = 12'hfff;
rom[13630] = 12'hfff;
rom[13631] = 12'hfff;
rom[13632] = 12'hfff;
rom[13633] = 12'hfff;
rom[13634] = 12'hfff;
rom[13635] = 12'hfff;
rom[13636] = 12'hfff;
rom[13637] = 12'hfff;
rom[13638] = 12'hfff;
rom[13639] = 12'hfff;
rom[13640] = 12'hfff;
rom[13641] = 12'hfff;
rom[13642] = 12'hfff;
rom[13643] = 12'hfff;
rom[13644] = 12'hfff;
rom[13645] = 12'hfff;
rom[13646] = 12'hfff;
rom[13647] = 12'hfff;
rom[13648] = 12'hfff;
rom[13649] = 12'hfff;
rom[13650] = 12'hfff;
rom[13651] = 12'hfff;
rom[13652] = 12'hfff;
rom[13653] = 12'hfff;
rom[13654] = 12'hfff;
rom[13655] = 12'hfff;
rom[13656] = 12'hfff;
rom[13657] = 12'hfff;
rom[13658] = 12'hfff;
rom[13659] = 12'hfff;
rom[13660] = 12'hfff;
rom[13661] = 12'hfff;
rom[13662] = 12'hfff;
rom[13663] = 12'hfff;
rom[13664] = 12'hfff;
rom[13665] = 12'hfff;
rom[13666] = 12'hfff;
rom[13667] = 12'hfff;
rom[13668] = 12'hfff;
rom[13669] = 12'hfff;
rom[13670] = 12'hfff;
rom[13671] = 12'hfff;
rom[13672] = 12'hfff;
rom[13673] = 12'hfff;
rom[13674] = 12'hfff;
rom[13675] = 12'hfff;
rom[13676] = 12'hfff;
rom[13677] = 12'hfff;
rom[13678] = 12'hfff;
rom[13679] = 12'hfff;
rom[13680] = 12'hfff;
rom[13681] = 12'hfff;
rom[13682] = 12'hfff;
rom[13683] = 12'hfff;
rom[13684] = 12'hfff;
rom[13685] = 12'hfff;
rom[13686] = 12'hfff;
rom[13687] = 12'hfff;
rom[13688] = 12'hfff;
rom[13689] = 12'hfff;
rom[13690] = 12'hfff;
rom[13691] = 12'hfff;
rom[13692] = 12'hfff;
rom[13693] = 12'hfff;
rom[13694] = 12'hfff;
rom[13695] = 12'hfff;
rom[13696] = 12'hfff;
rom[13697] = 12'hfff;
rom[13698] = 12'hfff;
rom[13699] = 12'hfff;
rom[13700] = 12'hfff;
rom[13701] = 12'hfff;
rom[13702] = 12'hfff;
rom[13703] = 12'hfff;
rom[13704] = 12'hfff;
rom[13705] = 12'hfff;
rom[13706] = 12'hfff;
rom[13707] = 12'hfff;
rom[13708] = 12'hfff;
rom[13709] = 12'hfff;
rom[13710] = 12'hfff;
rom[13711] = 12'hfff;
rom[13712] = 12'hfff;
rom[13713] = 12'hfff;
rom[13714] = 12'hfff;
rom[13715] = 12'hfff;
rom[13716] = 12'hfff;
rom[13717] = 12'hfff;
rom[13718] = 12'hfff;
rom[13719] = 12'hfff;
rom[13720] = 12'hfff;
rom[13721] = 12'hfff;
rom[13722] = 12'hfff;
rom[13723] = 12'hfff;
rom[13724] = 12'hfff;
rom[13725] = 12'hfff;
rom[13726] = 12'hfff;
rom[13727] = 12'hfff;
rom[13728] = 12'hfff;
rom[13729] = 12'hfff;
rom[13730] = 12'hfff;
rom[13731] = 12'hfff;
rom[13732] = 12'hfff;
rom[13733] = 12'hfff;
rom[13734] = 12'hfff;
rom[13735] = 12'hfff;
rom[13736] = 12'hfff;
rom[13737] = 12'hddf;
rom[13738] = 12'hccf;
rom[13739] = 12'hbbf;
rom[13740] = 12'haae;
rom[13741] = 12'h99e;
rom[13742] = 12'h88e;
rom[13743] = 12'h77e;
rom[13744] = 12'h77e;
rom[13745] = 12'h77e;
rom[13746] = 12'h88e;
rom[13747] = 12'h99e;
rom[13748] = 12'haae;
rom[13749] = 12'hccf;
rom[13750] = 12'hfff;
rom[13751] = 12'hfff;
rom[13752] = 12'hfff;
rom[13753] = 12'hfff;
rom[13754] = 12'hfff;
rom[13755] = 12'hfff;
rom[13756] = 12'hfff;
rom[13757] = 12'hfff;
rom[13758] = 12'hfff;
rom[13759] = 12'hfff;
rom[13760] = 12'hfff;
rom[13761] = 12'hfff;
rom[13762] = 12'hfff;
rom[13763] = 12'hfff;
rom[13764] = 12'hfff;
rom[13765] = 12'hfff;
rom[13766] = 12'hfff;
rom[13767] = 12'hfff;
rom[13768] = 12'hfff;
rom[13769] = 12'hfff;
rom[13770] = 12'hfff;
rom[13771] = 12'hfff;
rom[13772] = 12'hfff;
rom[13773] = 12'hfff;
rom[13774] = 12'hfff;
rom[13775] = 12'hfff;
rom[13776] = 12'hfff;
rom[13777] = 12'hfff;
rom[13778] = 12'hfff;
rom[13779] = 12'hfff;
rom[13780] = 12'hfff;
rom[13781] = 12'hfff;
rom[13782] = 12'hfff;
rom[13783] = 12'hfff;
rom[13784] = 12'hfff;
rom[13785] = 12'hfff;
rom[13786] = 12'hfff;
rom[13787] = 12'hfff;
rom[13788] = 12'hfff;
rom[13789] = 12'hfff;
rom[13790] = 12'hfff;
rom[13791] = 12'hfff;
rom[13792] = 12'hfff;
rom[13793] = 12'hfff;
rom[13794] = 12'hfff;
rom[13795] = 12'hfff;
rom[13796] = 12'hfff;
rom[13797] = 12'hfff;
rom[13798] = 12'hfff;
rom[13799] = 12'hfff;
rom[13800] = 12'hfff;
rom[13801] = 12'hfff;
rom[13802] = 12'hfff;
rom[13803] = 12'hfff;
rom[13804] = 12'hfff;
rom[13805] = 12'hfff;
rom[13806] = 12'hfff;
rom[13807] = 12'hfff;
rom[13808] = 12'hfff;
rom[13809] = 12'hfff;
rom[13810] = 12'hfff;
rom[13811] = 12'hfff;
rom[13812] = 12'hfff;
rom[13813] = 12'hfff;
rom[13814] = 12'hfff;
rom[13815] = 12'hfff;
rom[13816] = 12'hfff;
rom[13817] = 12'hfff;
rom[13818] = 12'hfff;
rom[13819] = 12'hfff;
rom[13820] = 12'hfff;
rom[13821] = 12'hfff;
rom[13822] = 12'hfff;
rom[13823] = 12'hfff;
rom[13824] = 12'hfff;
rom[13825] = 12'hfff;
rom[13826] = 12'hfff;
rom[13827] = 12'hfff;
rom[13828] = 12'hfff;
rom[13829] = 12'hfff;
rom[13830] = 12'hfff;
rom[13831] = 12'hfff;
rom[13832] = 12'hfff;
rom[13833] = 12'hfff;
rom[13834] = 12'hfff;
rom[13835] = 12'hfff;
rom[13836] = 12'hfff;
rom[13837] = 12'hfff;
rom[13838] = 12'hfff;
rom[13839] = 12'hfff;
rom[13840] = 12'hfff;
rom[13841] = 12'hfff;
rom[13842] = 12'hfff;
rom[13843] = 12'hfff;
rom[13844] = 12'hfff;
rom[13845] = 12'hfff;
rom[13846] = 12'hfff;
rom[13847] = 12'hfff;
rom[13848] = 12'hfff;
rom[13849] = 12'hfff;
rom[13850] = 12'hfff;
rom[13851] = 12'hfff;
rom[13852] = 12'hfff;
rom[13853] = 12'hfff;
rom[13854] = 12'hfff;
rom[13855] = 12'hfff;
rom[13856] = 12'hfff;
rom[13857] = 12'hfff;
rom[13858] = 12'hfff;
rom[13859] = 12'hfff;
rom[13860] = 12'hfff;
rom[13861] = 12'hfff;
rom[13862] = 12'hfff;
rom[13863] = 12'hfff;
rom[13864] = 12'hfff;
rom[13865] = 12'hfff;
rom[13866] = 12'hfff;
rom[13867] = 12'hfff;
rom[13868] = 12'hfff;
rom[13869] = 12'hfff;
rom[13870] = 12'hfff;
rom[13871] = 12'hfff;
rom[13872] = 12'hfff;
rom[13873] = 12'hfff;
rom[13874] = 12'hfff;
rom[13875] = 12'hfff;
rom[13876] = 12'hfff;
rom[13877] = 12'hfff;
rom[13878] = 12'hfff;
rom[13879] = 12'hfff;
rom[13880] = 12'hfff;
rom[13881] = 12'hfff;
rom[13882] = 12'hfff;
rom[13883] = 12'hfff;
rom[13884] = 12'hfff;
rom[13885] = 12'hfff;
rom[13886] = 12'hfff;
rom[13887] = 12'hfff;
rom[13888] = 12'hfff;
rom[13889] = 12'hfff;
rom[13890] = 12'hfff;
rom[13891] = 12'hfff;
rom[13892] = 12'hfff;
rom[13893] = 12'hfff;
rom[13894] = 12'hfff;
rom[13895] = 12'hfff;
rom[13896] = 12'hfff;
rom[13897] = 12'hfff;
rom[13898] = 12'hfff;
rom[13899] = 12'hfff;
rom[13900] = 12'hfff;
rom[13901] = 12'hfff;
rom[13902] = 12'hfff;
rom[13903] = 12'hfff;
rom[13904] = 12'hfff;
rom[13905] = 12'hfff;
rom[13906] = 12'hfff;
rom[13907] = 12'hfff;
rom[13908] = 12'hfff;
rom[13909] = 12'hfff;
rom[13910] = 12'hfff;
rom[13911] = 12'hfff;
rom[13912] = 12'hfff;
rom[13913] = 12'hfff;
rom[13914] = 12'hfff;
rom[13915] = 12'hfff;
rom[13916] = 12'hfff;
rom[13917] = 12'hfff;
rom[13918] = 12'hfff;
rom[13919] = 12'hfff;
rom[13920] = 12'hfff;
rom[13921] = 12'hfff;
rom[13922] = 12'hfff;
rom[13923] = 12'hfff;
rom[13924] = 12'hfff;
rom[13925] = 12'hfff;
rom[13926] = 12'hfff;
rom[13927] = 12'hfff;
rom[13928] = 12'hfff;
rom[13929] = 12'hfff;
rom[13930] = 12'hfff;
rom[13931] = 12'hfff;
rom[13932] = 12'hfff;
rom[13933] = 12'hfff;
rom[13934] = 12'hfff;
rom[13935] = 12'hfff;
rom[13936] = 12'hfff;
rom[13937] = 12'hfff;
rom[13938] = 12'hfff;
rom[13939] = 12'hfff;
rom[13940] = 12'hfff;
rom[13941] = 12'hfff;
rom[13942] = 12'hfff;
rom[13943] = 12'hfff;
rom[13944] = 12'hfff;
rom[13945] = 12'hfff;
rom[13946] = 12'hfff;
rom[13947] = 12'hfff;
rom[13948] = 12'hfff;
rom[13949] = 12'hfff;
rom[13950] = 12'hfff;
rom[13951] = 12'hfff;
rom[13952] = 12'hfff;
rom[13953] = 12'hfff;
rom[13954] = 12'hfff;
rom[13955] = 12'hfff;
rom[13956] = 12'hfff;
rom[13957] = 12'hfff;
rom[13958] = 12'hfff;
rom[13959] = 12'hfff;
rom[13960] = 12'hfff;
rom[13961] = 12'hfff;
rom[13962] = 12'hfff;
rom[13963] = 12'hfff;
rom[13964] = 12'hfff;
rom[13965] = 12'hfff;
rom[13966] = 12'hfff;
rom[13967] = 12'hfff;
rom[13968] = 12'hfff;
rom[13969] = 12'hfff;
rom[13970] = 12'hfff;
rom[13971] = 12'hfff;
rom[13972] = 12'hfff;
rom[13973] = 12'hfff;
rom[13974] = 12'hfff;
rom[13975] = 12'hfff;
rom[13976] = 12'hfff;
rom[13977] = 12'hfff;
rom[13978] = 12'hfff;
rom[13979] = 12'hfff;
rom[13980] = 12'hfff;
rom[13981] = 12'hfff;
rom[13982] = 12'hfff;
rom[13983] = 12'hfff;
rom[13984] = 12'hfff;
rom[13985] = 12'hfff;
rom[13986] = 12'hfff;
rom[13987] = 12'hfff;
rom[13988] = 12'hfff;
rom[13989] = 12'hfff;
rom[13990] = 12'hfff;
rom[13991] = 12'hfff;
rom[13992] = 12'hfff;
rom[13993] = 12'hfff;
rom[13994] = 12'hfff;
rom[13995] = 12'hfff;
rom[13996] = 12'hfff;
rom[13997] = 12'hfff;
rom[13998] = 12'hfff;
rom[13999] = 12'hfff;
rom[14000] = 12'hfff;
rom[14001] = 12'hfff;
rom[14002] = 12'hfff;
rom[14003] = 12'hfff;
rom[14004] = 12'hfff;
rom[14005] = 12'hfff;
rom[14006] = 12'hfff;
rom[14007] = 12'hfff;
rom[14008] = 12'hfff;
rom[14009] = 12'hfff;
rom[14010] = 12'hfff;
rom[14011] = 12'hfff;
rom[14012] = 12'hfff;
rom[14013] = 12'hfff;
rom[14014] = 12'hfff;
rom[14015] = 12'hfff;
rom[14016] = 12'hfff;
rom[14017] = 12'hfff;
rom[14018] = 12'hfff;
rom[14019] = 12'hfff;
rom[14020] = 12'hfff;
rom[14021] = 12'hfff;
rom[14022] = 12'hfff;
rom[14023] = 12'hfff;
rom[14024] = 12'hfff;
rom[14025] = 12'hfff;
rom[14026] = 12'hfff;
rom[14027] = 12'hfff;
rom[14028] = 12'hfff;
rom[14029] = 12'hfff;
rom[14030] = 12'hfff;
rom[14031] = 12'hfff;
rom[14032] = 12'hfff;
rom[14033] = 12'hfff;
rom[14034] = 12'hfff;
rom[14035] = 12'hfff;
rom[14036] = 12'hfff;
rom[14037] = 12'hfff;
rom[14038] = 12'hfff;
rom[14039] = 12'hfff;
rom[14040] = 12'hfff;
rom[14041] = 12'hfff;
rom[14042] = 12'hfff;
rom[14043] = 12'hfff;
rom[14044] = 12'hfff;
rom[14045] = 12'hfff;
rom[14046] = 12'hfff;
rom[14047] = 12'hfff;
rom[14048] = 12'hfff;
rom[14049] = 12'hfff;
rom[14050] = 12'hfff;
rom[14051] = 12'hfff;
rom[14052] = 12'hfff;
rom[14053] = 12'hfff;
rom[14054] = 12'hfff;
rom[14055] = 12'hfff;
rom[14056] = 12'hfff;
rom[14057] = 12'hfff;
rom[14058] = 12'hfff;
rom[14059] = 12'hfff;
rom[14060] = 12'hfff;
rom[14061] = 12'hfff;
rom[14062] = 12'hfff;
rom[14063] = 12'hfff;
rom[14064] = 12'hfff;
rom[14065] = 12'hfff;
rom[14066] = 12'hfff;
rom[14067] = 12'hfff;
rom[14068] = 12'hfff;
rom[14069] = 12'hfff;
rom[14070] = 12'hfff;
rom[14071] = 12'hfff;
rom[14072] = 12'hfff;
rom[14073] = 12'hfff;
rom[14074] = 12'hfff;
rom[14075] = 12'hfff;
rom[14076] = 12'hfff;
rom[14077] = 12'hfff;
rom[14078] = 12'hfff;
rom[14079] = 12'hfff;
rom[14080] = 12'hfff;
rom[14081] = 12'hfff;
rom[14082] = 12'hfff;
rom[14083] = 12'hfff;
rom[14084] = 12'hfff;
rom[14085] = 12'hfff;
rom[14086] = 12'hfff;
rom[14087] = 12'hfff;
rom[14088] = 12'hfff;
rom[14089] = 12'hfff;
rom[14090] = 12'hfff;
rom[14091] = 12'hfff;
rom[14092] = 12'hfff;
rom[14093] = 12'hfff;
rom[14094] = 12'hfff;
rom[14095] = 12'hfff;
rom[14096] = 12'hfff;
rom[14097] = 12'hfff;
rom[14098] = 12'hfff;
rom[14099] = 12'hfff;
rom[14100] = 12'hfff;
rom[14101] = 12'hfff;
rom[14102] = 12'hfff;
rom[14103] = 12'hfff;
rom[14104] = 12'hfff;
rom[14105] = 12'hfff;
rom[14106] = 12'hfff;
rom[14107] = 12'hfff;
rom[14108] = 12'hfff;
rom[14109] = 12'hfff;
rom[14110] = 12'hfff;
rom[14111] = 12'hfff;
rom[14112] = 12'hfff;
rom[14113] = 12'hfff;
rom[14114] = 12'hfff;
rom[14115] = 12'hfff;
rom[14116] = 12'hfff;
rom[14117] = 12'hfff;
rom[14118] = 12'hfff;
rom[14119] = 12'hfff;
rom[14120] = 12'hfff;
rom[14121] = 12'hfff;
rom[14122] = 12'hfff;
rom[14123] = 12'hfff;
rom[14124] = 12'hfff;
rom[14125] = 12'hfff;
rom[14126] = 12'hfff;
rom[14127] = 12'hfff;
rom[14128] = 12'hfff;
rom[14129] = 12'hfff;
rom[14130] = 12'hfff;
rom[14131] = 12'hfff;
rom[14132] = 12'hfff;
rom[14133] = 12'hfff;
rom[14134] = 12'hfff;
rom[14135] = 12'hfff;
rom[14136] = 12'hfff;
rom[14137] = 12'hfff;
rom[14138] = 12'hfff;
rom[14139] = 12'hfff;
rom[14140] = 12'hfff;
rom[14141] = 12'hfff;
rom[14142] = 12'hfff;
rom[14143] = 12'hfff;
rom[14144] = 12'hfff;
rom[14145] = 12'hfff;
rom[14146] = 12'hfff;
rom[14147] = 12'hfff;
rom[14148] = 12'hfff;
rom[14149] = 12'hfff;
rom[14150] = 12'hfff;
rom[14151] = 12'hfff;
rom[14152] = 12'hfff;
rom[14153] = 12'hfff;
rom[14154] = 12'hfff;
rom[14155] = 12'hfff;
rom[14156] = 12'hfff;
rom[14157] = 12'hfff;
rom[14158] = 12'hfff;
rom[14159] = 12'hfff;
rom[14160] = 12'hfff;
rom[14161] = 12'hfff;
rom[14162] = 12'hfff;
rom[14163] = 12'hfff;
rom[14164] = 12'hfff;
rom[14165] = 12'hfff;
rom[14166] = 12'hfff;
rom[14167] = 12'hfff;
rom[14168] = 12'hfff;
rom[14169] = 12'hfff;
rom[14170] = 12'hfff;
rom[14171] = 12'hfff;
rom[14172] = 12'hfff;
rom[14173] = 12'hfff;
rom[14174] = 12'hfff;
rom[14175] = 12'hfff;
rom[14176] = 12'hfff;
rom[14177] = 12'hfff;
rom[14178] = 12'hfff;
rom[14179] = 12'hfff;
rom[14180] = 12'hfff;
rom[14181] = 12'hfff;
rom[14182] = 12'hfff;
rom[14183] = 12'hfff;
rom[14184] = 12'hfff;
rom[14185] = 12'hfff;
rom[14186] = 12'hfff;
rom[14187] = 12'hfff;
rom[14188] = 12'hfff;
rom[14189] = 12'hfff;
rom[14190] = 12'hfff;
rom[14191] = 12'hfff;
rom[14192] = 12'hfff;
rom[14193] = 12'hfff;
rom[14194] = 12'hfff;
rom[14195] = 12'hfff;
rom[14196] = 12'hfff;
rom[14197] = 12'hfff;
rom[14198] = 12'hfff;
rom[14199] = 12'hfff;
rom[14200] = 12'hfff;
rom[14201] = 12'hfff;
rom[14202] = 12'hfff;
rom[14203] = 12'hfff;
rom[14204] = 12'hfff;
rom[14205] = 12'hfff;
rom[14206] = 12'hfff;
rom[14207] = 12'hfff;
rom[14208] = 12'hfff;
rom[14209] = 12'hfff;
rom[14210] = 12'hfff;
rom[14211] = 12'hfff;
rom[14212] = 12'hfff;
rom[14213] = 12'hfff;
rom[14214] = 12'hfff;
rom[14215] = 12'hfff;
rom[14216] = 12'hfff;
rom[14217] = 12'hfff;
rom[14218] = 12'hfff;
rom[14219] = 12'hfff;
rom[14220] = 12'hfff;
rom[14221] = 12'hfff;
rom[14222] = 12'hfff;
rom[14223] = 12'hfff;
rom[14224] = 12'hfff;
rom[14225] = 12'hfff;
rom[14226] = 12'hfff;
rom[14227] = 12'hfff;
rom[14228] = 12'hfff;
rom[14229] = 12'hfff;
rom[14230] = 12'hfff;
rom[14231] = 12'hfff;
rom[14232] = 12'hfff;
rom[14233] = 12'hfff;
rom[14234] = 12'hfff;
rom[14235] = 12'hfff;
rom[14236] = 12'hfff;
rom[14237] = 12'hfff;
rom[14238] = 12'hfff;
rom[14239] = 12'hfff;
rom[14240] = 12'hfff;
rom[14241] = 12'hfff;
rom[14242] = 12'hfff;
rom[14243] = 12'hfff;
rom[14244] = 12'hfff;
rom[14245] = 12'hfff;
rom[14246] = 12'hfff;
rom[14247] = 12'hfff;
rom[14248] = 12'hfff;
rom[14249] = 12'hfff;
rom[14250] = 12'hfff;
rom[14251] = 12'hfff;
rom[14252] = 12'hfff;
rom[14253] = 12'hfff;
rom[14254] = 12'hfff;
rom[14255] = 12'hfff;
rom[14256] = 12'hfff;
rom[14257] = 12'hfff;
rom[14258] = 12'hfff;
rom[14259] = 12'hfff;
rom[14260] = 12'hfff;
rom[14261] = 12'hfff;
rom[14262] = 12'hfff;
rom[14263] = 12'hfff;
rom[14264] = 12'hfff;
rom[14265] = 12'hfff;
rom[14266] = 12'hfff;
rom[14267] = 12'hfff;
rom[14268] = 12'hfff;
rom[14269] = 12'hfff;
rom[14270] = 12'hfff;
rom[14271] = 12'hfff;
rom[14272] = 12'hfff;
rom[14273] = 12'hfff;
rom[14274] = 12'hfff;
rom[14275] = 12'hfff;
rom[14276] = 12'hfff;
rom[14277] = 12'hfff;
rom[14278] = 12'hfff;
rom[14279] = 12'hfff;
rom[14280] = 12'hfff;
rom[14281] = 12'hfff;
rom[14282] = 12'hfff;
rom[14283] = 12'hfff;
rom[14284] = 12'hfff;
rom[14285] = 12'hfff;
rom[14286] = 12'hfff;
rom[14287] = 12'hfff;
rom[14288] = 12'hfff;
rom[14289] = 12'hfff;
rom[14290] = 12'hfff;
rom[14291] = 12'hfff;
rom[14292] = 12'hfff;
rom[14293] = 12'hfff;
rom[14294] = 12'hfff;
rom[14295] = 12'hfff;
rom[14296] = 12'hfff;
rom[14297] = 12'hfff;
rom[14298] = 12'hfff;
rom[14299] = 12'hfff;
rom[14300] = 12'hfff;
rom[14301] = 12'hfff;
rom[14302] = 12'hfff;
rom[14303] = 12'hfff;
rom[14304] = 12'hfff;
rom[14305] = 12'hfff;
rom[14306] = 12'hfff;
rom[14307] = 12'hfff;
rom[14308] = 12'hfff;
rom[14309] = 12'hfff;
rom[14310] = 12'hfff;
rom[14311] = 12'hfff;
rom[14312] = 12'hfff;
rom[14313] = 12'hfff;
rom[14314] = 12'hfff;
rom[14315] = 12'hfff;
rom[14316] = 12'hfff;
rom[14317] = 12'hfff;
rom[14318] = 12'hfff;
rom[14319] = 12'hfff;
rom[14320] = 12'hfff;
rom[14321] = 12'hfff;
rom[14322] = 12'hfff;
rom[14323] = 12'hfff;
rom[14324] = 12'hfff;
rom[14325] = 12'hfff;
rom[14326] = 12'hfff;
rom[14327] = 12'hfff;
rom[14328] = 12'hfff;
rom[14329] = 12'hfff;
rom[14330] = 12'hfff;
rom[14331] = 12'hfff;
rom[14332] = 12'hfff;
rom[14333] = 12'hfff;
rom[14334] = 12'hfff;
rom[14335] = 12'hfff;
rom[14336] = 12'hfff;
rom[14337] = 12'hfff;
rom[14338] = 12'hfff;
rom[14339] = 12'hfff;
rom[14340] = 12'hfff;
rom[14341] = 12'hfff;
rom[14342] = 12'hfff;
rom[14343] = 12'hfff;
rom[14344] = 12'hfff;
rom[14345] = 12'hfff;
rom[14346] = 12'hfff;
rom[14347] = 12'hfff;
rom[14348] = 12'hfff;
rom[14349] = 12'hfff;
rom[14350] = 12'hfff;
rom[14351] = 12'hfff;
rom[14352] = 12'hfff;
rom[14353] = 12'hfff;
rom[14354] = 12'hfff;
rom[14355] = 12'hfff;
rom[14356] = 12'hfff;
rom[14357] = 12'hfff;
rom[14358] = 12'hfff;
rom[14359] = 12'hfff;
rom[14360] = 12'hfff;
rom[14361] = 12'hfff;
rom[14362] = 12'hfff;
rom[14363] = 12'hfff;
rom[14364] = 12'hfff;
rom[14365] = 12'hfff;
rom[14366] = 12'hfff;
rom[14367] = 12'hfff;
rom[14368] = 12'hfff;
rom[14369] = 12'hfff;
rom[14370] = 12'hfff;
rom[14371] = 12'hfff;
rom[14372] = 12'hfff;
rom[14373] = 12'hfff;
rom[14374] = 12'hfff;
rom[14375] = 12'hfff;
rom[14376] = 12'hfff;
rom[14377] = 12'hfff;
rom[14378] = 12'hfff;
rom[14379] = 12'hfff;
rom[14380] = 12'hfff;
rom[14381] = 12'hfff;
rom[14382] = 12'hfff;
rom[14383] = 12'hfff;
rom[14384] = 12'hfff;
rom[14385] = 12'hfff;
rom[14386] = 12'hfff;
rom[14387] = 12'hfff;
rom[14388] = 12'hfff;
rom[14389] = 12'hfff;
rom[14390] = 12'hfff;
rom[14391] = 12'hfff;
rom[14392] = 12'hfff;
rom[14393] = 12'hfff;
rom[14394] = 12'hfff;
rom[14395] = 12'hfff;
rom[14396] = 12'hfff;
rom[14397] = 12'hfff;
rom[14398] = 12'hfff;
rom[14399] = 12'hfff;
rom[14400] = 12'hfff;
rom[14401] = 12'hfff;
rom[14402] = 12'hfff;
rom[14403] = 12'hfff;
rom[14404] = 12'hfff;
rom[14405] = 12'hfff;
rom[14406] = 12'hfff;
rom[14407] = 12'hfff;
rom[14408] = 12'hfff;
rom[14409] = 12'hfff;
rom[14410] = 12'hfff;
rom[14411] = 12'hfff;
rom[14412] = 12'hfff;
rom[14413] = 12'hfff;
rom[14414] = 12'hfff;
rom[14415] = 12'hfff;
rom[14416] = 12'hfff;
rom[14417] = 12'hfff;
rom[14418] = 12'hfff;
rom[14419] = 12'hfff;
rom[14420] = 12'hfff;
rom[14421] = 12'hfff;
rom[14422] = 12'hfff;
rom[14423] = 12'hfff;
rom[14424] = 12'hfff;
rom[14425] = 12'hfff;
rom[14426] = 12'hfff;
rom[14427] = 12'hfff;
rom[14428] = 12'hfff;
rom[14429] = 12'hfff;
rom[14430] = 12'hfff;
rom[14431] = 12'hfff;
rom[14432] = 12'hfff;
rom[14433] = 12'hfff;
rom[14434] = 12'hfff;
rom[14435] = 12'hfff;
rom[14436] = 12'hfff;
rom[14437] = 12'hfff;
rom[14438] = 12'hfff;
rom[14439] = 12'hfff;
rom[14440] = 12'hfff;
rom[14441] = 12'hfff;
rom[14442] = 12'hfff;
rom[14443] = 12'hfff;
rom[14444] = 12'hfff;
rom[14445] = 12'hfff;
rom[14446] = 12'hfff;
rom[14447] = 12'hfff;
rom[14448] = 12'hfff;
rom[14449] = 12'hfff;
rom[14450] = 12'hfff;
rom[14451] = 12'hfff;
rom[14452] = 12'hfff;
rom[14453] = 12'hfff;
rom[14454] = 12'hfff;
rom[14455] = 12'hfff;
rom[14456] = 12'hfff;
rom[14457] = 12'hfff;
rom[14458] = 12'hfff;
rom[14459] = 12'hfff;
rom[14460] = 12'hfff;
rom[14461] = 12'hfff;
rom[14462] = 12'hfff;
rom[14463] = 12'hfff;
rom[14464] = 12'hfff;
rom[14465] = 12'hfff;
rom[14466] = 12'hfff;
rom[14467] = 12'hfff;
rom[14468] = 12'hfff;
rom[14469] = 12'hfff;
rom[14470] = 12'hfff;
rom[14471] = 12'hfff;
rom[14472] = 12'hfff;
rom[14473] = 12'hfff;
rom[14474] = 12'hfff;
rom[14475] = 12'hfff;
rom[14476] = 12'hfff;
rom[14477] = 12'hfff;
rom[14478] = 12'hfff;
rom[14479] = 12'hfff;
rom[14480] = 12'hfff;
rom[14481] = 12'hfff;
rom[14482] = 12'hfff;
rom[14483] = 12'hfff;
rom[14484] = 12'hfff;
rom[14485] = 12'hfff;
rom[14486] = 12'hfff;
rom[14487] = 12'hfff;
rom[14488] = 12'hfff;
rom[14489] = 12'hfff;
rom[14490] = 12'hfff;
rom[14491] = 12'hfff;
rom[14492] = 12'hfff;
rom[14493] = 12'hfff;
rom[14494] = 12'hfff;
rom[14495] = 12'hfff;
rom[14496] = 12'hfff;
rom[14497] = 12'hfff;
rom[14498] = 12'hfff;
rom[14499] = 12'hfff;
rom[14500] = 12'hfff;
rom[14501] = 12'hfff;
rom[14502] = 12'hfff;
rom[14503] = 12'hfff;
rom[14504] = 12'hfff;
rom[14505] = 12'hfff;
rom[14506] = 12'hfff;
rom[14507] = 12'hfff;
rom[14508] = 12'hfff;
rom[14509] = 12'hfff;
rom[14510] = 12'hfff;
rom[14511] = 12'hfff;
rom[14512] = 12'hfff;
rom[14513] = 12'hfff;
rom[14514] = 12'hfff;
rom[14515] = 12'hfff;
rom[14516] = 12'hfff;
rom[14517] = 12'hfff;
rom[14518] = 12'hfff;
rom[14519] = 12'hfff;
rom[14520] = 12'hfff;
rom[14521] = 12'hfff;
rom[14522] = 12'hfff;
rom[14523] = 12'hfff;
rom[14524] = 12'hfff;
rom[14525] = 12'hfff;
rom[14526] = 12'hfff;
rom[14527] = 12'hfff;
rom[14528] = 12'hfff;
rom[14529] = 12'hfff;
rom[14530] = 12'hfff;
rom[14531] = 12'hfff;
rom[14532] = 12'hfff;
rom[14533] = 12'hfff;
rom[14534] = 12'hfff;
rom[14535] = 12'hfff;
rom[14536] = 12'hfff;
rom[14537] = 12'hfff;
rom[14538] = 12'hfff;
rom[14539] = 12'hfff;
rom[14540] = 12'hfff;
rom[14541] = 12'hfff;
rom[14542] = 12'hfff;
rom[14543] = 12'hfff;
rom[14544] = 12'hfff;
rom[14545] = 12'hfff;
rom[14546] = 12'hfff;
rom[14547] = 12'hfff;
rom[14548] = 12'hfff;
rom[14549] = 12'hfff;
rom[14550] = 12'hfff;
rom[14551] = 12'hfff;
rom[14552] = 12'hfff;
rom[14553] = 12'hfff;
rom[14554] = 12'hfff;
rom[14555] = 12'hfff;
rom[14556] = 12'hfff;
rom[14557] = 12'hfff;
rom[14558] = 12'hfff;
rom[14559] = 12'hfff;
rom[14560] = 12'hfff;
rom[14561] = 12'hfff;
rom[14562] = 12'hfff;
rom[14563] = 12'hfff;
rom[14564] = 12'hfff;
rom[14565] = 12'hfff;
rom[14566] = 12'hfff;
rom[14567] = 12'hfff;
rom[14568] = 12'hfff;
rom[14569] = 12'hfff;
rom[14570] = 12'hfff;
rom[14571] = 12'hfff;
rom[14572] = 12'hfff;
rom[14573] = 12'hfff;
rom[14574] = 12'hfff;
rom[14575] = 12'hfff;
rom[14576] = 12'hfff;
rom[14577] = 12'hfff;
rom[14578] = 12'hfff;
rom[14579] = 12'hfff;
rom[14580] = 12'hfff;
rom[14581] = 12'hfff;
rom[14582] = 12'hfff;
rom[14583] = 12'hfff;
rom[14584] = 12'hfff;
rom[14585] = 12'hfff;
rom[14586] = 12'hfff;
rom[14587] = 12'hfff;
rom[14588] = 12'hfff;
rom[14589] = 12'hfff;
rom[14590] = 12'hfff;
rom[14591] = 12'hfff;
rom[14592] = 12'hfff;
rom[14593] = 12'hfff;
rom[14594] = 12'hfff;
rom[14595] = 12'hfff;
rom[14596] = 12'hfff;
rom[14597] = 12'hfff;
rom[14598] = 12'hfff;
rom[14599] = 12'hfff;
rom[14600] = 12'hfff;
rom[14601] = 12'hfff;
rom[14602] = 12'hfff;
rom[14603] = 12'hfff;
rom[14604] = 12'hfff;
rom[14605] = 12'hfff;
rom[14606] = 12'hfff;
rom[14607] = 12'hfff;
rom[14608] = 12'hfff;
rom[14609] = 12'hfff;
rom[14610] = 12'hfff;
rom[14611] = 12'hfff;
rom[14612] = 12'hfff;
rom[14613] = 12'hfff;
rom[14614] = 12'hfff;
rom[14615] = 12'hfff;
rom[14616] = 12'hfff;
rom[14617] = 12'hfff;
rom[14618] = 12'hfff;
rom[14619] = 12'hfff;
rom[14620] = 12'hfff;
rom[14621] = 12'hfff;
rom[14622] = 12'hfff;
rom[14623] = 12'hfff;
rom[14624] = 12'hfff;
rom[14625] = 12'hfff;
rom[14626] = 12'hfff;
rom[14627] = 12'hfff;
rom[14628] = 12'hfff;
rom[14629] = 12'hfff;
rom[14630] = 12'hfff;
rom[14631] = 12'hfff;
rom[14632] = 12'hfff;
rom[14633] = 12'hfff;
rom[14634] = 12'hfff;
rom[14635] = 12'hfff;
rom[14636] = 12'hfff;
rom[14637] = 12'hfff;
rom[14638] = 12'hfff;
rom[14639] = 12'hfff;
rom[14640] = 12'hfff;
rom[14641] = 12'hfff;
rom[14642] = 12'hfff;
rom[14643] = 12'hfff;
rom[14644] = 12'hfff;
rom[14645] = 12'hfff;
rom[14646] = 12'hfff;
rom[14647] = 12'hfff;
rom[14648] = 12'hfff;
rom[14649] = 12'hfff;
rom[14650] = 12'hfff;
rom[14651] = 12'hfff;
rom[14652] = 12'hfff;
rom[14653] = 12'hfff;
rom[14654] = 12'hfff;
rom[14655] = 12'hfff;
rom[14656] = 12'hfff;
rom[14657] = 12'hfff;
rom[14658] = 12'hfff;
rom[14659] = 12'hfff;
rom[14660] = 12'hfff;
rom[14661] = 12'hfff;
rom[14662] = 12'hfff;
rom[14663] = 12'hfff;
rom[14664] = 12'hfff;
rom[14665] = 12'hfff;
rom[14666] = 12'hfff;
rom[14667] = 12'hfff;
rom[14668] = 12'hfff;
rom[14669] = 12'hfff;
rom[14670] = 12'hfff;
rom[14671] = 12'hfff;
rom[14672] = 12'hfff;
rom[14673] = 12'hfff;
rom[14674] = 12'hfff;
rom[14675] = 12'hfff;
rom[14676] = 12'hfff;
rom[14677] = 12'hfff;
rom[14678] = 12'hfff;
rom[14679] = 12'hfff;
rom[14680] = 12'hfff;
rom[14681] = 12'hfff;
rom[14682] = 12'hfff;
rom[14683] = 12'hfff;
rom[14684] = 12'hfff;
rom[14685] = 12'hfff;
rom[14686] = 12'hfff;
rom[14687] = 12'hfff;
rom[14688] = 12'hfff;
rom[14689] = 12'hfff;
rom[14690] = 12'hfff;
rom[14691] = 12'hfff;
rom[14692] = 12'hfff;
rom[14693] = 12'hfff;
rom[14694] = 12'hfff;
rom[14695] = 12'hfff;
rom[14696] = 12'hfff;
rom[14697] = 12'hfff;
rom[14698] = 12'hfff;
rom[14699] = 12'hfff;
rom[14700] = 12'hfff;
rom[14701] = 12'hfff;
rom[14702] = 12'hfff;
rom[14703] = 12'hfff;
rom[14704] = 12'hfff;
rom[14705] = 12'hfff;
rom[14706] = 12'hfff;
rom[14707] = 12'hfff;
rom[14708] = 12'hfff;
rom[14709] = 12'hfff;
rom[14710] = 12'hfff;
rom[14711] = 12'hfff;
rom[14712] = 12'hfff;
rom[14713] = 12'hfff;
rom[14714] = 12'hfff;
rom[14715] = 12'hfff;
rom[14716] = 12'hfff;
rom[14717] = 12'hfff;
rom[14718] = 12'hfff;
rom[14719] = 12'hfff;
rom[14720] = 12'hfff;
rom[14721] = 12'hfff;
rom[14722] = 12'hfff;
rom[14723] = 12'hfff;
rom[14724] = 12'hfff;
rom[14725] = 12'hfff;
rom[14726] = 12'hfff;
rom[14727] = 12'hfff;
rom[14728] = 12'hfff;
rom[14729] = 12'hfff;
rom[14730] = 12'hfff;
rom[14731] = 12'hfff;
rom[14732] = 12'hfff;
rom[14733] = 12'hfff;
rom[14734] = 12'hfff;
rom[14735] = 12'hfff;
rom[14736] = 12'hfff;
rom[14737] = 12'hfff;
rom[14738] = 12'hfff;
rom[14739] = 12'hfff;
rom[14740] = 12'hfff;
rom[14741] = 12'hfff;
rom[14742] = 12'hfff;
rom[14743] = 12'hfff;
rom[14744] = 12'hfff;
rom[14745] = 12'hfff;
rom[14746] = 12'hfff;
rom[14747] = 12'hfff;
rom[14748] = 12'hfff;
rom[14749] = 12'hfff;
rom[14750] = 12'hfff;
rom[14751] = 12'hfff;
rom[14752] = 12'hfff;
rom[14753] = 12'hfff;
rom[14754] = 12'hfff;
rom[14755] = 12'hfff;
rom[14756] = 12'hfff;
rom[14757] = 12'hfff;
rom[14758] = 12'hfff;
rom[14759] = 12'hfff;
rom[14760] = 12'hfff;
rom[14761] = 12'hfff;
rom[14762] = 12'hfff;
rom[14763] = 12'hfff;
rom[14764] = 12'hfff;
rom[14765] = 12'hfff;
rom[14766] = 12'hfff;
rom[14767] = 12'hfff;
rom[14768] = 12'hfff;
rom[14769] = 12'hfff;
rom[14770] = 12'hfff;
rom[14771] = 12'hfff;
rom[14772] = 12'hfff;
rom[14773] = 12'hfff;
rom[14774] = 12'hfff;
rom[14775] = 12'hfff;
rom[14776] = 12'hfff;
rom[14777] = 12'hfff;
rom[14778] = 12'hfff;
rom[14779] = 12'hfff;
rom[14780] = 12'hfff;
rom[14781] = 12'hfff;
rom[14782] = 12'hfff;
rom[14783] = 12'hfff;
rom[14784] = 12'hfff;
rom[14785] = 12'hfff;
rom[14786] = 12'hfff;
rom[14787] = 12'hfff;
rom[14788] = 12'hfff;
rom[14789] = 12'hfff;
rom[14790] = 12'hfff;
rom[14791] = 12'hfff;
rom[14792] = 12'hfff;
rom[14793] = 12'hfff;
rom[14794] = 12'hfff;
rom[14795] = 12'hfff;
rom[14796] = 12'hfff;
rom[14797] = 12'hfff;
rom[14798] = 12'hfff;
rom[14799] = 12'hfff;
rom[14800] = 12'hfff;
rom[14801] = 12'hfff;
rom[14802] = 12'hfff;
rom[14803] = 12'hfff;
rom[14804] = 12'hfff;
rom[14805] = 12'hfff;
rom[14806] = 12'hfff;
rom[14807] = 12'hfff;
rom[14808] = 12'hfff;
rom[14809] = 12'hfff;
rom[14810] = 12'hfff;
rom[14811] = 12'hfff;
rom[14812] = 12'hfff;
rom[14813] = 12'hfff;
rom[14814] = 12'hfff;
rom[14815] = 12'hfff;
rom[14816] = 12'hfff;
rom[14817] = 12'hfff;
rom[14818] = 12'hfff;
rom[14819] = 12'hfff;
rom[14820] = 12'hfff;
rom[14821] = 12'hfff;
rom[14822] = 12'hfff;
rom[14823] = 12'hfff;
rom[14824] = 12'hfff;
rom[14825] = 12'hfff;
rom[14826] = 12'hfff;
rom[14827] = 12'hfff;
rom[14828] = 12'hfff;
rom[14829] = 12'hfff;
rom[14830] = 12'hfff;
rom[14831] = 12'hfff;
rom[14832] = 12'hfff;
rom[14833] = 12'hfff;
rom[14834] = 12'hfff;
rom[14835] = 12'hfff;
rom[14836] = 12'hfff;
rom[14837] = 12'hfff;
rom[14838] = 12'hfff;
rom[14839] = 12'hfff;
rom[14840] = 12'hfff;
rom[14841] = 12'hfff;
rom[14842] = 12'hfff;
rom[14843] = 12'hfff;
rom[14844] = 12'hfff;
rom[14845] = 12'hfff;
rom[14846] = 12'hfff;
rom[14847] = 12'hfff;
rom[14848] = 12'hfff;
rom[14849] = 12'hfff;
rom[14850] = 12'hfff;
rom[14851] = 12'hfff;
rom[14852] = 12'hfff;
rom[14853] = 12'hfff;
rom[14854] = 12'hfff;
rom[14855] = 12'hfff;
rom[14856] = 12'hfff;
rom[14857] = 12'hfff;
rom[14858] = 12'hfff;
rom[14859] = 12'hfff;
rom[14860] = 12'hfff;
rom[14861] = 12'hfff;
rom[14862] = 12'hfff;
rom[14863] = 12'hfff;
rom[14864] = 12'hfff;
rom[14865] = 12'hfff;
rom[14866] = 12'hfff;
rom[14867] = 12'hfff;
rom[14868] = 12'hfff;
rom[14869] = 12'hfff;
rom[14870] = 12'hfff;
rom[14871] = 12'hfff;
rom[14872] = 12'hfff;
rom[14873] = 12'hfff;
rom[14874] = 12'hfff;
rom[14875] = 12'hfff;
rom[14876] = 12'hfff;
rom[14877] = 12'hfff;
rom[14878] = 12'hfff;
rom[14879] = 12'hfff;
rom[14880] = 12'hfff;
rom[14881] = 12'hfff;
rom[14882] = 12'hfff;
rom[14883] = 12'hfff;
rom[14884] = 12'hfff;
rom[14885] = 12'hfff;
rom[14886] = 12'hfff;
rom[14887] = 12'hfff;
rom[14888] = 12'hfff;
rom[14889] = 12'hfff;
rom[14890] = 12'hfff;
rom[14891] = 12'hfff;
rom[14892] = 12'hfff;
rom[14893] = 12'hfff;
rom[14894] = 12'hfff;
rom[14895] = 12'hfff;
rom[14896] = 12'hfff;
rom[14897] = 12'hfff;
rom[14898] = 12'hfff;
rom[14899] = 12'hfff;
rom[14900] = 12'hfff;
rom[14901] = 12'hfff;
rom[14902] = 12'hfff;
rom[14903] = 12'hfff;
rom[14904] = 12'hfff;
rom[14905] = 12'hfff;
rom[14906] = 12'hfff;
rom[14907] = 12'hfff;
rom[14908] = 12'hfff;
rom[14909] = 12'hfff;
rom[14910] = 12'hfff;
rom[14911] = 12'hfff;
rom[14912] = 12'hfff;
rom[14913] = 12'hfff;
rom[14914] = 12'hfff;
rom[14915] = 12'hfff;
rom[14916] = 12'hfff;
rom[14917] = 12'hfff;
rom[14918] = 12'hfff;
rom[14919] = 12'hfff;
rom[14920] = 12'hfff;
rom[14921] = 12'hfff;
rom[14922] = 12'hfff;
rom[14923] = 12'hfff;
rom[14924] = 12'hfff;
rom[14925] = 12'hfff;
rom[14926] = 12'hfff;
rom[14927] = 12'hfff;
rom[14928] = 12'hfff;
rom[14929] = 12'hfff;
rom[14930] = 12'hfff;
rom[14931] = 12'hfff;
rom[14932] = 12'hfff;
rom[14933] = 12'hfff;
rom[14934] = 12'hfff;
rom[14935] = 12'hfff;
rom[14936] = 12'hfff;
rom[14937] = 12'hfff;
rom[14938] = 12'hfff;
rom[14939] = 12'hfff;
rom[14940] = 12'hfff;
rom[14941] = 12'hfff;
rom[14942] = 12'hfff;
rom[14943] = 12'hfff;
rom[14944] = 12'hfff;
rom[14945] = 12'hfff;
rom[14946] = 12'hfff;
rom[14947] = 12'hfff;
rom[14948] = 12'hfff;
rom[14949] = 12'hfff;
rom[14950] = 12'hfff;
rom[14951] = 12'hfff;
rom[14952] = 12'hfff;
rom[14953] = 12'hfff;
rom[14954] = 12'hfff;
rom[14955] = 12'hfff;
rom[14956] = 12'hfff;
rom[14957] = 12'hfff;
rom[14958] = 12'hfff;
rom[14959] = 12'hfff;
rom[14960] = 12'hfff;
rom[14961] = 12'hfff;
rom[14962] = 12'hfff;
rom[14963] = 12'hfff;
rom[14964] = 12'hfff;
rom[14965] = 12'hfff;
rom[14966] = 12'hfff;
rom[14967] = 12'hfff;
rom[14968] = 12'hfff;
rom[14969] = 12'hfff;
rom[14970] = 12'hfff;
rom[14971] = 12'hfff;
rom[14972] = 12'hfff;
rom[14973] = 12'hfff;
rom[14974] = 12'hfff;
rom[14975] = 12'hfff;
rom[14976] = 12'hfff;
rom[14977] = 12'hfff;
rom[14978] = 12'hfff;
rom[14979] = 12'hfff;
rom[14980] = 12'hfff;
rom[14981] = 12'hfff;
rom[14982] = 12'hfff;
rom[14983] = 12'hfff;
rom[14984] = 12'hfff;
rom[14985] = 12'hfff;
rom[14986] = 12'hfff;
rom[14987] = 12'hfff;
rom[14988] = 12'hfff;
rom[14989] = 12'hfff;
rom[14990] = 12'hfff;
rom[14991] = 12'hfff;
rom[14992] = 12'hfff;
rom[14993] = 12'hfff;
rom[14994] = 12'hfff;
rom[14995] = 12'hfff;
rom[14996] = 12'hfff;
rom[14997] = 12'hfff;
rom[14998] = 12'hfff;
rom[14999] = 12'hfff;
rom[15000] = 12'hfff;
rom[15001] = 12'hfff;
rom[15002] = 12'hfff;
rom[15003] = 12'hfff;
rom[15004] = 12'hfff;
rom[15005] = 12'hfff;
rom[15006] = 12'hfff;
rom[15007] = 12'hfff;
rom[15008] = 12'hfff;
rom[15009] = 12'hfff;
rom[15010] = 12'hfff;
rom[15011] = 12'hfff;
rom[15012] = 12'hfff;
rom[15013] = 12'hfff;
rom[15014] = 12'hfff;
rom[15015] = 12'hfff;
rom[15016] = 12'hfff;
rom[15017] = 12'hfff;
rom[15018] = 12'hfff;
rom[15019] = 12'hfff;
rom[15020] = 12'hfff;
rom[15021] = 12'hfff;
rom[15022] = 12'hfff;
rom[15023] = 12'hfff;
rom[15024] = 12'hfff;
rom[15025] = 12'hfff;
rom[15026] = 12'hfff;
rom[15027] = 12'hfff;
rom[15028] = 12'hfff;
rom[15029] = 12'hfff;
rom[15030] = 12'hfff;
rom[15031] = 12'hfff;
rom[15032] = 12'hfff;
rom[15033] = 12'hfff;
rom[15034] = 12'hfff;
rom[15035] = 12'hfff;
rom[15036] = 12'hfff;
rom[15037] = 12'hfff;
rom[15038] = 12'hfff;
rom[15039] = 12'hfff;
rom[15040] = 12'hfff;
rom[15041] = 12'hfff;
rom[15042] = 12'hfff;
rom[15043] = 12'hfff;
rom[15044] = 12'hfff;
rom[15045] = 12'hfff;
rom[15046] = 12'hfff;
rom[15047] = 12'hfff;
rom[15048] = 12'hfff;
rom[15049] = 12'hfff;
rom[15050] = 12'hfff;
rom[15051] = 12'hfff;
rom[15052] = 12'hfff;
rom[15053] = 12'hfff;
rom[15054] = 12'hfff;
rom[15055] = 12'hfff;
rom[15056] = 12'hfff;
rom[15057] = 12'hfff;
rom[15058] = 12'hfff;
rom[15059] = 12'hfff;
rom[15060] = 12'hfff;
rom[15061] = 12'hfff;
rom[15062] = 12'hfff;
rom[15063] = 12'hfff;
rom[15064] = 12'hfff;
rom[15065] = 12'hfff;
rom[15066] = 12'hfff;
rom[15067] = 12'hfff;
rom[15068] = 12'hfff;
rom[15069] = 12'hfff;
rom[15070] = 12'hfff;
rom[15071] = 12'hfff;
rom[15072] = 12'hfff;
rom[15073] = 12'hfff;
rom[15074] = 12'hfff;
rom[15075] = 12'hfff;
rom[15076] = 12'hfff;
rom[15077] = 12'hfff;
rom[15078] = 12'hfff;
rom[15079] = 12'hfff;
rom[15080] = 12'hfff;
rom[15081] = 12'hfff;
rom[15082] = 12'hfff;
rom[15083] = 12'hfff;
rom[15084] = 12'hfff;
rom[15085] = 12'hfff;
rom[15086] = 12'hfff;
rom[15087] = 12'hfff;
rom[15088] = 12'hfff;
rom[15089] = 12'hfff;
rom[15090] = 12'hfff;
rom[15091] = 12'hfff;
rom[15092] = 12'hfff;
rom[15093] = 12'hfff;
rom[15094] = 12'hfff;
rom[15095] = 12'hfff;
rom[15096] = 12'hfff;
rom[15097] = 12'hfff;
rom[15098] = 12'hfff;
rom[15099] = 12'hfff;
rom[15100] = 12'hfff;
rom[15101] = 12'hfff;
rom[15102] = 12'hfff;
rom[15103] = 12'hfff;
rom[15104] = 12'hfff;
rom[15105] = 12'hfff;
rom[15106] = 12'hfff;
rom[15107] = 12'hfff;
rom[15108] = 12'hfff;
rom[15109] = 12'hfff;
rom[15110] = 12'hfff;
rom[15111] = 12'hfff;
rom[15112] = 12'hfff;
rom[15113] = 12'hfff;
rom[15114] = 12'hfff;
rom[15115] = 12'hfff;
rom[15116] = 12'hfff;
rom[15117] = 12'hfff;
rom[15118] = 12'hfff;
rom[15119] = 12'hfff;
rom[15120] = 12'hfff;
rom[15121] = 12'hfff;
rom[15122] = 12'hfff;
rom[15123] = 12'hfff;
rom[15124] = 12'hfff;
rom[15125] = 12'hfff;
rom[15126] = 12'hfff;
rom[15127] = 12'hfff;
rom[15128] = 12'hfff;
rom[15129] = 12'hfff;
rom[15130] = 12'hfff;
rom[15131] = 12'hfff;
rom[15132] = 12'hfff;
rom[15133] = 12'hfff;
rom[15134] = 12'hfff;
rom[15135] = 12'hfff;
rom[15136] = 12'hfff;
rom[15137] = 12'hfff;
rom[15138] = 12'hfff;
rom[15139] = 12'hfff;
rom[15140] = 12'hfff;
rom[15141] = 12'hfff;
rom[15142] = 12'hfff;
rom[15143] = 12'hfff;
rom[15144] = 12'hfff;
rom[15145] = 12'hfff;
rom[15146] = 12'hfff;
rom[15147] = 12'hfff;
rom[15148] = 12'hfff;
rom[15149] = 12'hfff;
rom[15150] = 12'hfff;
rom[15151] = 12'hfff;
rom[15152] = 12'hfff;
rom[15153] = 12'hfff;
rom[15154] = 12'hfff;
rom[15155] = 12'hfff;
rom[15156] = 12'hfff;
rom[15157] = 12'hfff;
rom[15158] = 12'hfff;
rom[15159] = 12'hfff;
rom[15160] = 12'hfff;
rom[15161] = 12'hfff;
rom[15162] = 12'hfff;
rom[15163] = 12'hfff;
rom[15164] = 12'hfff;
rom[15165] = 12'hfff;
rom[15166] = 12'hfff;
rom[15167] = 12'hfff;
rom[15168] = 12'hfff;
rom[15169] = 12'hfff;
rom[15170] = 12'hfff;
rom[15171] = 12'hfff;
rom[15172] = 12'hfff;
rom[15173] = 12'hfff;
rom[15174] = 12'hfff;
rom[15175] = 12'hfff;
rom[15176] = 12'hfff;
rom[15177] = 12'hfff;
rom[15178] = 12'hfff;
rom[15179] = 12'hfff;
rom[15180] = 12'hfff;
rom[15181] = 12'hfff;
rom[15182] = 12'hfff;
rom[15183] = 12'hfff;
rom[15184] = 12'hfff;
rom[15185] = 12'hfff;
rom[15186] = 12'hfff;
rom[15187] = 12'hfff;
rom[15188] = 12'hfff;
rom[15189] = 12'hfff;
rom[15190] = 12'hfff;
rom[15191] = 12'hfff;
rom[15192] = 12'hfff;
rom[15193] = 12'hfff;
rom[15194] = 12'hfff;
rom[15195] = 12'hfff;
rom[15196] = 12'hfff;
rom[15197] = 12'hfff;
rom[15198] = 12'hfff;
rom[15199] = 12'hfff;
rom[15200] = 12'hfff;
rom[15201] = 12'hfff;
rom[15202] = 12'hfff;
rom[15203] = 12'hfff;
rom[15204] = 12'hfff;
rom[15205] = 12'hfff;
rom[15206] = 12'hfff;
rom[15207] = 12'hfff;
rom[15208] = 12'hfff;
rom[15209] = 12'hfff;
rom[15210] = 12'hfff;
rom[15211] = 12'hfff;
rom[15212] = 12'hfff;
rom[15213] = 12'hfff;
rom[15214] = 12'hfff;
rom[15215] = 12'hfff;
rom[15216] = 12'hfff;
rom[15217] = 12'hfff;
rom[15218] = 12'hfff;
rom[15219] = 12'hfff;
rom[15220] = 12'hfff;
rom[15221] = 12'hfff;
rom[15222] = 12'hfff;
rom[15223] = 12'hfff;
rom[15224] = 12'hfff;
rom[15225] = 12'hfff;
rom[15226] = 12'hfff;
rom[15227] = 12'hfff;
rom[15228] = 12'hfff;
rom[15229] = 12'hfff;
rom[15230] = 12'hfff;
rom[15231] = 12'hfff;
rom[15232] = 12'hfff;
rom[15233] = 12'hfff;
rom[15234] = 12'hfff;
rom[15235] = 12'hfff;
rom[15236] = 12'hfff;
rom[15237] = 12'hfff;
rom[15238] = 12'hfff;
rom[15239] = 12'hfff;
rom[15240] = 12'hfff;
rom[15241] = 12'hfff;
rom[15242] = 12'hfff;
rom[15243] = 12'hfff;
rom[15244] = 12'hfff;
rom[15245] = 12'hfff;
rom[15246] = 12'hfff;
rom[15247] = 12'hfff;
rom[15248] = 12'hfff;
rom[15249] = 12'hfff;
rom[15250] = 12'hfff;
rom[15251] = 12'hfff;
rom[15252] = 12'hfff;
rom[15253] = 12'hfff;
rom[15254] = 12'hfff;
rom[15255] = 12'hfff;
rom[15256] = 12'hfff;
rom[15257] = 12'hfff;
rom[15258] = 12'hfff;
rom[15259] = 12'hfff;
rom[15260] = 12'hfff;
rom[15261] = 12'hfff;
rom[15262] = 12'hfff;
rom[15263] = 12'hfff;
rom[15264] = 12'hfff;
rom[15265] = 12'hfff;
rom[15266] = 12'hfff;
rom[15267] = 12'hfff;
rom[15268] = 12'hfff;
rom[15269] = 12'hfff;
rom[15270] = 12'hfff;
rom[15271] = 12'hfff;
rom[15272] = 12'hfff;
rom[15273] = 12'hfff;
rom[15274] = 12'hfff;
rom[15275] = 12'hfff;
rom[15276] = 12'hfff;
rom[15277] = 12'hfff;
rom[15278] = 12'hfff;
rom[15279] = 12'hfff;
rom[15280] = 12'hfff;
rom[15281] = 12'hfff;
rom[15282] = 12'hfff;
rom[15283] = 12'hfff;
rom[15284] = 12'hfff;
rom[15285] = 12'hfff;
rom[15286] = 12'hfff;
rom[15287] = 12'hfff;
rom[15288] = 12'hfff;
rom[15289] = 12'hfff;
rom[15290] = 12'hfff;
rom[15291] = 12'hfff;
rom[15292] = 12'hfff;
rom[15293] = 12'hfff;
rom[15294] = 12'hfff;
rom[15295] = 12'hfff;
rom[15296] = 12'hfff;
rom[15297] = 12'hfff;
rom[15298] = 12'hfff;
rom[15299] = 12'hfff;
rom[15300] = 12'hfff;
rom[15301] = 12'hfff;
rom[15302] = 12'hfff;
rom[15303] = 12'hfff;
rom[15304] = 12'hfff;
rom[15305] = 12'hfff;
rom[15306] = 12'hfff;
rom[15307] = 12'hfff;
rom[15308] = 12'hfff;
rom[15309] = 12'hfff;
rom[15310] = 12'hfff;
rom[15311] = 12'hfff;
rom[15312] = 12'hfff;
rom[15313] = 12'hfff;
rom[15314] = 12'hfff;
rom[15315] = 12'hfff;
rom[15316] = 12'hfff;
rom[15317] = 12'hfff;
rom[15318] = 12'hfff;
rom[15319] = 12'hfff;
rom[15320] = 12'hfff;
rom[15321] = 12'hfff;
rom[15322] = 12'hfff;
rom[15323] = 12'hfff;
rom[15324] = 12'hfff;
rom[15325] = 12'hfff;
rom[15326] = 12'hfff;
rom[15327] = 12'hfff;
rom[15328] = 12'hfff;
rom[15329] = 12'hfff;
rom[15330] = 12'hfff;
rom[15331] = 12'hfff;
rom[15332] = 12'hfff;
rom[15333] = 12'hfff;
rom[15334] = 12'hfff;
rom[15335] = 12'hfff;
rom[15336] = 12'hfff;
rom[15337] = 12'hfff;
rom[15338] = 12'hfff;
rom[15339] = 12'hfff;
rom[15340] = 12'hfff;
rom[15341] = 12'hfff;
rom[15342] = 12'hfff;
rom[15343] = 12'hfff;
rom[15344] = 12'hfff;
rom[15345] = 12'hfff;
rom[15346] = 12'hfff;
rom[15347] = 12'hfff;
rom[15348] = 12'hfff;
rom[15349] = 12'hfff;
rom[15350] = 12'hfff;
rom[15351] = 12'hfff;
rom[15352] = 12'hfff;
rom[15353] = 12'hfff;
rom[15354] = 12'hfff;
rom[15355] = 12'hfff;
rom[15356] = 12'hfff;
rom[15357] = 12'hfff;
rom[15358] = 12'hfff;
rom[15359] = 12'hfff;
rom[15360] = 12'hfff;
rom[15361] = 12'hfff;
rom[15362] = 12'hfff;
rom[15363] = 12'hfff;
rom[15364] = 12'hfff;
rom[15365] = 12'hfff;
rom[15366] = 12'hfff;
rom[15367] = 12'hfff;
rom[15368] = 12'hfff;
rom[15369] = 12'hfff;
rom[15370] = 12'hfff;
rom[15371] = 12'hfff;
rom[15372] = 12'hfff;
rom[15373] = 12'hfff;
rom[15374] = 12'hfff;
rom[15375] = 12'hfff;
rom[15376] = 12'hfff;
rom[15377] = 12'hfff;
rom[15378] = 12'hfff;
rom[15379] = 12'hfff;
rom[15380] = 12'hfff;
rom[15381] = 12'hfff;
rom[15382] = 12'hfff;
rom[15383] = 12'hfff;
rom[15384] = 12'hfff;
rom[15385] = 12'hfff;
rom[15386] = 12'hfff;
rom[15387] = 12'hfff;
rom[15388] = 12'hfff;
rom[15389] = 12'hfff;
rom[15390] = 12'hfff;
rom[15391] = 12'hfff;
rom[15392] = 12'hfff;
rom[15393] = 12'hfff;
rom[15394] = 12'hfff;
rom[15395] = 12'hfff;
rom[15396] = 12'hfff;
rom[15397] = 12'hfff;
rom[15398] = 12'hfff;
rom[15399] = 12'hfff;
rom[15400] = 12'hfff;
rom[15401] = 12'hfff;
rom[15402] = 12'hfff;
rom[15403] = 12'hfff;
rom[15404] = 12'hfff;
rom[15405] = 12'hfff;
rom[15406] = 12'hfff;
rom[15407] = 12'hfff;
rom[15408] = 12'hfff;
rom[15409] = 12'hfff;
rom[15410] = 12'hfff;
rom[15411] = 12'hfff;
rom[15412] = 12'hfff;
rom[15413] = 12'hfff;
rom[15414] = 12'hfff;
rom[15415] = 12'hfff;
rom[15416] = 12'hfff;
rom[15417] = 12'hfff;
rom[15418] = 12'hfff;
rom[15419] = 12'hfff;
rom[15420] = 12'hfff;
rom[15421] = 12'hfff;
rom[15422] = 12'hfff;
rom[15423] = 12'hfff;
rom[15424] = 12'hfff;
rom[15425] = 12'hfff;
rom[15426] = 12'hfff;
rom[15427] = 12'hfff;
rom[15428] = 12'hfff;
rom[15429] = 12'hfff;
rom[15430] = 12'hfff;
rom[15431] = 12'hfff;
rom[15432] = 12'hfff;
rom[15433] = 12'hfff;
rom[15434] = 12'hfff;
rom[15435] = 12'hfff;
rom[15436] = 12'hfff;
rom[15437] = 12'hfff;
rom[15438] = 12'hfff;
rom[15439] = 12'hfff;
rom[15440] = 12'hfff;
rom[15441] = 12'hfff;
rom[15442] = 12'hfff;
rom[15443] = 12'hfff;
rom[15444] = 12'hfff;
rom[15445] = 12'hfff;
rom[15446] = 12'hfff;
rom[15447] = 12'hfff;
rom[15448] = 12'hfff;
rom[15449] = 12'hfff;
rom[15450] = 12'hfff;
rom[15451] = 12'hfff;
rom[15452] = 12'hfff;
rom[15453] = 12'hfff;
rom[15454] = 12'hfff;
rom[15455] = 12'hfff;
rom[15456] = 12'hfff;
rom[15457] = 12'hfff;
rom[15458] = 12'hfff;
rom[15459] = 12'hfff;
rom[15460] = 12'hfff;
rom[15461] = 12'hfff;
rom[15462] = 12'hfff;
rom[15463] = 12'hfff;
rom[15464] = 12'hfff;
rom[15465] = 12'hfff;
rom[15466] = 12'hfff;
rom[15467] = 12'hfff;
rom[15468] = 12'hfff;
rom[15469] = 12'hfff;
rom[15470] = 12'hfff;
rom[15471] = 12'hfff;
rom[15472] = 12'hfff;
rom[15473] = 12'hfff;
rom[15474] = 12'hfff;
rom[15475] = 12'hfff;
rom[15476] = 12'hfff;
rom[15477] = 12'hfff;
rom[15478] = 12'hfff;
rom[15479] = 12'hfff;
rom[15480] = 12'hfff;
rom[15481] = 12'hfff;
rom[15482] = 12'hfff;
rom[15483] = 12'hfff;
rom[15484] = 12'hfff;
rom[15485] = 12'hfff;
rom[15486] = 12'hfff;
rom[15487] = 12'hfff;
rom[15488] = 12'hfff;
rom[15489] = 12'hfff;
rom[15490] = 12'hfff;
rom[15491] = 12'hfff;
rom[15492] = 12'hfff;
rom[15493] = 12'hfff;
rom[15494] = 12'hfff;
rom[15495] = 12'hfff;
rom[15496] = 12'hfff;
rom[15497] = 12'hfff;
rom[15498] = 12'hfff;
rom[15499] = 12'hfff;
rom[15500] = 12'hfff;
rom[15501] = 12'hfff;
rom[15502] = 12'hfff;
rom[15503] = 12'hfff;
rom[15504] = 12'hfff;
rom[15505] = 12'hfff;
rom[15506] = 12'hfff;
rom[15507] = 12'hfff;
rom[15508] = 12'hfff;
rom[15509] = 12'hfff;
rom[15510] = 12'hfff;
rom[15511] = 12'hfff;
rom[15512] = 12'hfff;
rom[15513] = 12'hfff;
rom[15514] = 12'hfff;
rom[15515] = 12'hfff;
rom[15516] = 12'hfff;
rom[15517] = 12'hfff;
rom[15518] = 12'hfff;
rom[15519] = 12'hfff;
rom[15520] = 12'hfff;
rom[15521] = 12'hfff;
rom[15522] = 12'hfff;
rom[15523] = 12'hfff;
rom[15524] = 12'hfff;
rom[15525] = 12'hfff;
rom[15526] = 12'hfff;
rom[15527] = 12'hfff;
rom[15528] = 12'hfff;
rom[15529] = 12'hfff;
rom[15530] = 12'hfff;
rom[15531] = 12'hfff;
rom[15532] = 12'hfff;
rom[15533] = 12'hfff;
rom[15534] = 12'hfff;
rom[15535] = 12'hfff;
rom[15536] = 12'hfff;
rom[15537] = 12'hfff;
rom[15538] = 12'hfff;
rom[15539] = 12'hfff;
rom[15540] = 12'hfff;
rom[15541] = 12'hfff;
rom[15542] = 12'hfff;
rom[15543] = 12'hfff;
rom[15544] = 12'hfff;
rom[15545] = 12'hfff;
rom[15546] = 12'hfff;
rom[15547] = 12'hfff;
rom[15548] = 12'hfff;
rom[15549] = 12'hfff;
rom[15550] = 12'hfff;
rom[15551] = 12'hfff;
rom[15552] = 12'hfff;
rom[15553] = 12'hfff;
rom[15554] = 12'hfff;
rom[15555] = 12'hfff;
rom[15556] = 12'hfff;
rom[15557] = 12'hfff;
rom[15558] = 12'hfff;
rom[15559] = 12'hfff;
rom[15560] = 12'hfff;
rom[15561] = 12'hfff;
rom[15562] = 12'hfff;
rom[15563] = 12'hfff;
rom[15564] = 12'hfff;
rom[15565] = 12'hfff;
rom[15566] = 12'hfff;
rom[15567] = 12'hfff;
rom[15568] = 12'hfff;
rom[15569] = 12'hfff;
rom[15570] = 12'hfff;
rom[15571] = 12'hfff;
rom[15572] = 12'hfff;
rom[15573] = 12'hfff;
rom[15574] = 12'hfff;
rom[15575] = 12'hfff;
rom[15576] = 12'hfff;
rom[15577] = 12'hfff;
rom[15578] = 12'hfff;
rom[15579] = 12'hfff;
rom[15580] = 12'hfff;
rom[15581] = 12'hfff;
rom[15582] = 12'hfff;
rom[15583] = 12'hfff;
rom[15584] = 12'hfff;
rom[15585] = 12'hfff;
rom[15586] = 12'hfff;
rom[15587] = 12'hfff;
rom[15588] = 12'hfff;
rom[15589] = 12'hfff;
rom[15590] = 12'hfff;
rom[15591] = 12'hfff;
rom[15592] = 12'hfff;
rom[15593] = 12'hfff;
rom[15594] = 12'hfff;
rom[15595] = 12'hfff;
rom[15596] = 12'hfff;
rom[15597] = 12'hfff;
rom[15598] = 12'hfff;
rom[15599] = 12'hfff;
rom[15600] = 12'hfff;
rom[15601] = 12'hfff;
rom[15602] = 12'hfff;
rom[15603] = 12'hfff;
rom[15604] = 12'hfff;
rom[15605] = 12'hfff;
rom[15606] = 12'hfff;
rom[15607] = 12'hfff;
rom[15608] = 12'hfff;
rom[15609] = 12'hfff;
rom[15610] = 12'hfff;
rom[15611] = 12'hfff;
rom[15612] = 12'hfff;
rom[15613] = 12'hfff;
rom[15614] = 12'hfff;
rom[15615] = 12'hfff;
rom[15616] = 12'hfff;
rom[15617] = 12'hfff;
rom[15618] = 12'hfff;
rom[15619] = 12'hfff;
rom[15620] = 12'hfff;
rom[15621] = 12'hfff;
rom[15622] = 12'hfff;
rom[15623] = 12'hfff;
rom[15624] = 12'hfff;
rom[15625] = 12'hfff;
rom[15626] = 12'hfff;
rom[15627] = 12'hfff;
rom[15628] = 12'hfff;
rom[15629] = 12'hfff;
rom[15630] = 12'hfff;
rom[15631] = 12'hfff;
rom[15632] = 12'hfff;
rom[15633] = 12'hfff;
rom[15634] = 12'hfff;
rom[15635] = 12'hfff;
rom[15636] = 12'hfff;
rom[15637] = 12'hfff;
rom[15638] = 12'hfff;
rom[15639] = 12'hfff;
rom[15640] = 12'hfff;
rom[15641] = 12'hfff;
rom[15642] = 12'hfff;
rom[15643] = 12'hfff;
rom[15644] = 12'hfff;
rom[15645] = 12'hfff;
rom[15646] = 12'hfff;
rom[15647] = 12'hfff;
rom[15648] = 12'hfff;
rom[15649] = 12'hfff;
rom[15650] = 12'hfff;
rom[15651] = 12'hfff;
rom[15652] = 12'hfff;
rom[15653] = 12'hfff;
rom[15654] = 12'hfff;
rom[15655] = 12'hfff;
rom[15656] = 12'hfff;
rom[15657] = 12'hfff;
rom[15658] = 12'hfff;
rom[15659] = 12'hfff;
rom[15660] = 12'hfff;
rom[15661] = 12'hfff;
rom[15662] = 12'hfff;
rom[15663] = 12'hfff;
rom[15664] = 12'hfff;
rom[15665] = 12'hfff;
rom[15666] = 12'hfff;
rom[15667] = 12'hfff;
rom[15668] = 12'hfff;
rom[15669] = 12'hfff;
rom[15670] = 12'hfff;
rom[15671] = 12'hfff;
rom[15672] = 12'hfff;
rom[15673] = 12'hfff;
rom[15674] = 12'hfff;
rom[15675] = 12'hfff;
rom[15676] = 12'hfff;
rom[15677] = 12'hfff;
rom[15678] = 12'hfff;
rom[15679] = 12'hfff;
rom[15680] = 12'hfff;
rom[15681] = 12'hfff;
rom[15682] = 12'hfff;
rom[15683] = 12'hfff;
rom[15684] = 12'hfff;
rom[15685] = 12'hfff;
rom[15686] = 12'hfff;
rom[15687] = 12'hfff;
rom[15688] = 12'hfff;
rom[15689] = 12'hfff;
rom[15690] = 12'hfff;
rom[15691] = 12'hfff;
rom[15692] = 12'hfff;
rom[15693] = 12'hfff;
rom[15694] = 12'hfff;
rom[15695] = 12'hfff;
rom[15696] = 12'hfff;
rom[15697] = 12'hfff;
rom[15698] = 12'hfff;
rom[15699] = 12'hfff;
rom[15700] = 12'hfff;
rom[15701] = 12'hfff;
rom[15702] = 12'hfff;
rom[15703] = 12'hfff;
rom[15704] = 12'hfff;
rom[15705] = 12'hfff;
rom[15706] = 12'hfff;
rom[15707] = 12'hfff;
rom[15708] = 12'hfff;
rom[15709] = 12'hfff;
rom[15710] = 12'hfff;
rom[15711] = 12'hfff;
rom[15712] = 12'hfff;
rom[15713] = 12'hfff;
rom[15714] = 12'hfff;
rom[15715] = 12'hfff;
rom[15716] = 12'hfff;
rom[15717] = 12'hfff;
rom[15718] = 12'hfff;
rom[15719] = 12'hfff;
rom[15720] = 12'hfff;
rom[15721] = 12'hfff;
rom[15722] = 12'hfff;
rom[15723] = 12'hfff;
rom[15724] = 12'hfff;
rom[15725] = 12'hfff;
rom[15726] = 12'hfff;
rom[15727] = 12'hfff;
rom[15728] = 12'hfff;
rom[15729] = 12'hfff;
rom[15730] = 12'hfff;
rom[15731] = 12'hfff;
rom[15732] = 12'hfff;
rom[15733] = 12'hfff;
rom[15734] = 12'hfff;
rom[15735] = 12'hfff;
rom[15736] = 12'hfff;
rom[15737] = 12'hfff;
rom[15738] = 12'hfff;
rom[15739] = 12'hfff;
rom[15740] = 12'hfff;
rom[15741] = 12'hfff;
rom[15742] = 12'hfff;
rom[15743] = 12'hfff;
rom[15744] = 12'hfff;
rom[15745] = 12'hfff;
rom[15746] = 12'hfff;
rom[15747] = 12'hfff;
rom[15748] = 12'hfff;
rom[15749] = 12'hfff;
rom[15750] = 12'hfff;
rom[15751] = 12'hfff;
rom[15752] = 12'hfff;
rom[15753] = 12'hfff;
rom[15754] = 12'hfff;
rom[15755] = 12'hfff;
rom[15756] = 12'hfff;
rom[15757] = 12'hfff;
rom[15758] = 12'hfff;
rom[15759] = 12'hfff;
rom[15760] = 12'hfff;
rom[15761] = 12'hfff;
rom[15762] = 12'hfff;
rom[15763] = 12'hfff;
rom[15764] = 12'hfff;
rom[15765] = 12'hfff;
rom[15766] = 12'hfff;
rom[15767] = 12'hfff;
rom[15768] = 12'hfff;
rom[15769] = 12'hfff;
rom[15770] = 12'hfff;
rom[15771] = 12'hfff;
rom[15772] = 12'hfff;
rom[15773] = 12'hfff;
rom[15774] = 12'hfff;
rom[15775] = 12'hfff;
rom[15776] = 12'hfff;
rom[15777] = 12'hfff;
rom[15778] = 12'hfff;
rom[15779] = 12'hfff;
rom[15780] = 12'hfff;
rom[15781] = 12'hfff;
rom[15782] = 12'hfff;
rom[15783] = 12'hfff;
rom[15784] = 12'hfff;
rom[15785] = 12'hfff;
rom[15786] = 12'hfff;
rom[15787] = 12'hfff;
rom[15788] = 12'hfff;
rom[15789] = 12'hfff;
rom[15790] = 12'hfff;
rom[15791] = 12'hfff;
rom[15792] = 12'hfff;
rom[15793] = 12'hfff;
rom[15794] = 12'hfff;
rom[15795] = 12'hfff;
rom[15796] = 12'hfff;
rom[15797] = 12'hfff;
rom[15798] = 12'hfff;
rom[15799] = 12'hfff;
rom[15800] = 12'hfff;
rom[15801] = 12'hfff;
rom[15802] = 12'hfff;
rom[15803] = 12'hfff;
rom[15804] = 12'hfff;
rom[15805] = 12'hfff;
rom[15806] = 12'hfff;
rom[15807] = 12'hfff;
rom[15808] = 12'hfff;
rom[15809] = 12'hfff;
rom[15810] = 12'hfff;
rom[15811] = 12'hfff;
rom[15812] = 12'hfff;
rom[15813] = 12'hfff;
rom[15814] = 12'hfff;
rom[15815] = 12'hfff;
rom[15816] = 12'hfff;
rom[15817] = 12'hfff;
rom[15818] = 12'hfff;
rom[15819] = 12'hfff;
rom[15820] = 12'hfff;
rom[15821] = 12'hfff;
rom[15822] = 12'hfff;
rom[15823] = 12'hfff;
rom[15824] = 12'hfff;
rom[15825] = 12'hfff;
rom[15826] = 12'hfff;
rom[15827] = 12'hfff;
rom[15828] = 12'hfff;
rom[15829] = 12'hfff;
rom[15830] = 12'hfff;
rom[15831] = 12'hfff;
rom[15832] = 12'hfff;
rom[15833] = 12'hfff;
rom[15834] = 12'hfff;
rom[15835] = 12'hfff;
rom[15836] = 12'hfff;
rom[15837] = 12'hfff;
rom[15838] = 12'hfff;
rom[15839] = 12'hfff;
rom[15840] = 12'hfff;
rom[15841] = 12'hfff;
rom[15842] = 12'hfff;
rom[15843] = 12'hfff;
rom[15844] = 12'hfff;
rom[15845] = 12'hfff;
rom[15846] = 12'hfff;
rom[15847] = 12'hfff;
rom[15848] = 12'hfff;
rom[15849] = 12'hfff;
rom[15850] = 12'hfff;
rom[15851] = 12'hfff;
rom[15852] = 12'hfff;
rom[15853] = 12'hfff;
rom[15854] = 12'hfff;
rom[15855] = 12'hfff;
rom[15856] = 12'hfff;
rom[15857] = 12'hfff;
rom[15858] = 12'hfff;
rom[15859] = 12'hfff;
rom[15860] = 12'hfff;
rom[15861] = 12'hfff;
rom[15862] = 12'hfff;
rom[15863] = 12'hfff;
rom[15864] = 12'hfff;
rom[15865] = 12'hfff;
rom[15866] = 12'hfff;
rom[15867] = 12'hfff;
rom[15868] = 12'hfff;
rom[15869] = 12'hfff;
rom[15870] = 12'hfff;
rom[15871] = 12'hfff;
rom[15872] = 12'hfff;
rom[15873] = 12'hfff;
rom[15874] = 12'hfff;
rom[15875] = 12'hfff;
rom[15876] = 12'hfff;
rom[15877] = 12'hfff;
rom[15878] = 12'hfff;
rom[15879] = 12'hfff;
rom[15880] = 12'hfff;
rom[15881] = 12'hfff;
rom[15882] = 12'hfff;
rom[15883] = 12'hfff;
rom[15884] = 12'hfff;
rom[15885] = 12'hfff;
rom[15886] = 12'hfff;
rom[15887] = 12'hfff;
rom[15888] = 12'hfff;
rom[15889] = 12'hfff;
rom[15890] = 12'hfff;
rom[15891] = 12'hfff;
rom[15892] = 12'hfff;
rom[15893] = 12'hfff;
rom[15894] = 12'hfff;
rom[15895] = 12'hfff;
rom[15896] = 12'hfff;
rom[15897] = 12'hfff;
rom[15898] = 12'hfff;
rom[15899] = 12'hfff;
rom[15900] = 12'hfff;
rom[15901] = 12'hfff;
rom[15902] = 12'hfff;
rom[15903] = 12'hfff;
rom[15904] = 12'hfff;
rom[15905] = 12'hfff;
rom[15906] = 12'hfff;
rom[15907] = 12'hfff;
rom[15908] = 12'hfff;
rom[15909] = 12'hfff;
rom[15910] = 12'hfff;
rom[15911] = 12'hfff;
rom[15912] = 12'hfff;
rom[15913] = 12'hfff;
rom[15914] = 12'hfff;
rom[15915] = 12'hfff;
rom[15916] = 12'hfff;
rom[15917] = 12'hfff;
rom[15918] = 12'hfff;
rom[15919] = 12'hfff;
rom[15920] = 12'hfff;
rom[15921] = 12'hfff;
rom[15922] = 12'hfff;
rom[15923] = 12'hfff;
rom[15924] = 12'hfff;
rom[15925] = 12'hfff;
rom[15926] = 12'hfff;
rom[15927] = 12'hfff;
rom[15928] = 12'hfff;
rom[15929] = 12'hfff;
rom[15930] = 12'hfff;
rom[15931] = 12'hfff;
rom[15932] = 12'hfff;
rom[15933] = 12'hfff;
rom[15934] = 12'hfff;
rom[15935] = 12'hfff;
rom[15936] = 12'hfff;
rom[15937] = 12'hfff;
rom[15938] = 12'hfff;
rom[15939] = 12'hfff;
rom[15940] = 12'hfff;
rom[15941] = 12'hfff;
rom[15942] = 12'hfff;
rom[15943] = 12'hfff;
rom[15944] = 12'hfff;
rom[15945] = 12'hfff;
rom[15946] = 12'hfff;
rom[15947] = 12'hfff;
rom[15948] = 12'hfff;
rom[15949] = 12'hfff;
rom[15950] = 12'hfff;
rom[15951] = 12'hfff;
rom[15952] = 12'hfff;
rom[15953] = 12'hfff;
rom[15954] = 12'hfff;
rom[15955] = 12'hfff;
rom[15956] = 12'hfff;
rom[15957] = 12'hfff;
rom[15958] = 12'hfff;
rom[15959] = 12'hfff;
rom[15960] = 12'hfff;
rom[15961] = 12'hfff;
rom[15962] = 12'hfff;
rom[15963] = 12'hfff;
rom[15964] = 12'hfff;
rom[15965] = 12'hfff;
rom[15966] = 12'hfff;
rom[15967] = 12'hfff;
rom[15968] = 12'hfff;
rom[15969] = 12'hfff;
rom[15970] = 12'hfff;
rom[15971] = 12'hfff;
rom[15972] = 12'hfff;
rom[15973] = 12'hfff;
rom[15974] = 12'hfff;
rom[15975] = 12'hfff;
rom[15976] = 12'hfff;
rom[15977] = 12'hfff;
rom[15978] = 12'hfff;
rom[15979] = 12'hfff;
rom[15980] = 12'hfff;
rom[15981] = 12'hfff;
rom[15982] = 12'hfff;
rom[15983] = 12'hfff;
rom[15984] = 12'hfff;
rom[15985] = 12'hfff;
rom[15986] = 12'hfff;
rom[15987] = 12'hfff;
rom[15988] = 12'hfff;
rom[15989] = 12'hfff;
rom[15990] = 12'hfff;
rom[15991] = 12'hfff;
rom[15992] = 12'hfff;
rom[15993] = 12'hfff;
rom[15994] = 12'hfff;
rom[15995] = 12'hfff;
rom[15996] = 12'hfff;
rom[15997] = 12'hfff;
rom[15998] = 12'hfff;
rom[15999] = 12'hfff;
rom[16000] = 12'hfff;
rom[16001] = 12'hfff;
rom[16002] = 12'hfff;
rom[16003] = 12'hfff;
rom[16004] = 12'hfff;
rom[16005] = 12'hfff;
rom[16006] = 12'hfff;
rom[16007] = 12'hfff;
rom[16008] = 12'hfff;
rom[16009] = 12'hfff;
rom[16010] = 12'hfff;
rom[16011] = 12'hfff;
rom[16012] = 12'hfff;
rom[16013] = 12'hfff;
rom[16014] = 12'hfff;
rom[16015] = 12'hfff;
rom[16016] = 12'hfff;
rom[16017] = 12'hfff;
rom[16018] = 12'hfff;
rom[16019] = 12'hfff;
rom[16020] = 12'hfff;
rom[16021] = 12'hfff;
rom[16022] = 12'hfff;
rom[16023] = 12'hfff;
rom[16024] = 12'hfff;
rom[16025] = 12'hfff;
rom[16026] = 12'hfff;
rom[16027] = 12'hfff;
rom[16028] = 12'hfff;
rom[16029] = 12'hfff;
rom[16030] = 12'hfff;
rom[16031] = 12'hfff;
rom[16032] = 12'hfff;
rom[16033] = 12'hfff;
rom[16034] = 12'hfff;
rom[16035] = 12'hfff;
rom[16036] = 12'hfff;
rom[16037] = 12'hfff;
rom[16038] = 12'hfff;
rom[16039] = 12'hfff;
rom[16040] = 12'hfff;
rom[16041] = 12'hfff;
rom[16042] = 12'hfff;
rom[16043] = 12'hfff;
rom[16044] = 12'hfff;
rom[16045] = 12'hfff;
rom[16046] = 12'hfff;
rom[16047] = 12'hfff;
rom[16048] = 12'hfff;
rom[16049] = 12'hfff;
rom[16050] = 12'hfff;
rom[16051] = 12'hfff;
rom[16052] = 12'hfff;
rom[16053] = 12'hfff;
rom[16054] = 12'hfff;
rom[16055] = 12'hfff;
rom[16056] = 12'hfff;
rom[16057] = 12'hfff;
rom[16058] = 12'hfff;
rom[16059] = 12'hfff;
rom[16060] = 12'hfff;
rom[16061] = 12'hfff;
rom[16062] = 12'hfff;
rom[16063] = 12'hfff;
rom[16064] = 12'hfff;
rom[16065] = 12'hfff;
rom[16066] = 12'hfff;
rom[16067] = 12'hfff;
rom[16068] = 12'hfff;
rom[16069] = 12'hfff;
rom[16070] = 12'hfff;
rom[16071] = 12'hfff;
rom[16072] = 12'hfff;
rom[16073] = 12'hfff;
rom[16074] = 12'hfff;
rom[16075] = 12'hfff;
rom[16076] = 12'hfff;
rom[16077] = 12'hfff;
rom[16078] = 12'hfff;
rom[16079] = 12'hfff;
rom[16080] = 12'hfff;
rom[16081] = 12'hfff;
rom[16082] = 12'hfff;
rom[16083] = 12'hfff;
rom[16084] = 12'hfff;
rom[16085] = 12'hfff;
rom[16086] = 12'hfff;
rom[16087] = 12'hfff;
rom[16088] = 12'hfff;
rom[16089] = 12'hfff;
rom[16090] = 12'hfff;
rom[16091] = 12'hfff;
rom[16092] = 12'hfff;
rom[16093] = 12'hfff;
rom[16094] = 12'hfff;
rom[16095] = 12'hfff;
rom[16096] = 12'hfff;
rom[16097] = 12'hfff;
rom[16098] = 12'hfff;
rom[16099] = 12'hfff;
rom[16100] = 12'hfff;
rom[16101] = 12'hfff;
rom[16102] = 12'hfff;
rom[16103] = 12'hfff;
rom[16104] = 12'hfff;
rom[16105] = 12'hfff;
rom[16106] = 12'hfff;
rom[16107] = 12'hfff;
rom[16108] = 12'hfff;
rom[16109] = 12'hfff;
rom[16110] = 12'hfff;
rom[16111] = 12'hfff;
rom[16112] = 12'hfff;
rom[16113] = 12'hfff;
rom[16114] = 12'hfff;
rom[16115] = 12'hfff;
rom[16116] = 12'hfff;
rom[16117] = 12'hfff;
rom[16118] = 12'hfff;
rom[16119] = 12'hfff;
rom[16120] = 12'hfff;
rom[16121] = 12'hfff;
rom[16122] = 12'hfff;
rom[16123] = 12'hfff;
rom[16124] = 12'hfff;
rom[16125] = 12'hfff;
rom[16126] = 12'hfff;
rom[16127] = 12'hfff;
rom[16128] = 12'hfff;
rom[16129] = 12'hfff;
rom[16130] = 12'hfff;
rom[16131] = 12'hfff;
rom[16132] = 12'hfff;
rom[16133] = 12'hfff;
rom[16134] = 12'hfff;
rom[16135] = 12'hfff;
rom[16136] = 12'hfff;
rom[16137] = 12'hfff;
rom[16138] = 12'hfff;
rom[16139] = 12'hfff;
rom[16140] = 12'hfff;
rom[16141] = 12'hfff;
rom[16142] = 12'hfff;
rom[16143] = 12'hfff;
rom[16144] = 12'hfff;
rom[16145] = 12'hfff;
rom[16146] = 12'hfff;
rom[16147] = 12'hfff;
rom[16148] = 12'hfff;
rom[16149] = 12'hfff;
rom[16150] = 12'hfff;
rom[16151] = 12'hfff;
rom[16152] = 12'hfff;
rom[16153] = 12'hfff;
rom[16154] = 12'hfff;
rom[16155] = 12'hfff;
rom[16156] = 12'hfff;
rom[16157] = 12'hfff;
rom[16158] = 12'hfff;
rom[16159] = 12'hfff;
rom[16160] = 12'hfff;
rom[16161] = 12'hfff;
rom[16162] = 12'hfff;
rom[16163] = 12'hfff;
rom[16164] = 12'hfff;
rom[16165] = 12'hfff;
rom[16166] = 12'hfff;
rom[16167] = 12'hfff;
rom[16168] = 12'hfff;
rom[16169] = 12'hfff;
rom[16170] = 12'hfff;
rom[16171] = 12'hfff;
rom[16172] = 12'hfff;
rom[16173] = 12'hfff;
rom[16174] = 12'hfff;
rom[16175] = 12'hfff;
rom[16176] = 12'hfff;
rom[16177] = 12'hfff;
rom[16178] = 12'hfff;
rom[16179] = 12'hfff;
rom[16180] = 12'hfff;
rom[16181] = 12'hfff;
rom[16182] = 12'hfff;
rom[16183] = 12'hfff;
rom[16184] = 12'hfff;
rom[16185] = 12'hfff;
rom[16186] = 12'hfff;
rom[16187] = 12'hfff;
rom[16188] = 12'hfff;
rom[16189] = 12'hfff;
rom[16190] = 12'hfff;
rom[16191] = 12'hfff;
rom[16192] = 12'hfff;
rom[16193] = 12'hfff;
rom[16194] = 12'hfff;
rom[16195] = 12'hfff;
rom[16196] = 12'hfff;
rom[16197] = 12'hfff;
rom[16198] = 12'hfff;
rom[16199] = 12'hfff;
rom[16200] = 12'hfff;
rom[16201] = 12'hfff;
rom[16202] = 12'hfff;
rom[16203] = 12'hfff;
rom[16204] = 12'hfff;
rom[16205] = 12'hfff;
rom[16206] = 12'hfff;
rom[16207] = 12'hfff;
rom[16208] = 12'hfff;
rom[16209] = 12'hfff;
rom[16210] = 12'hfff;
rom[16211] = 12'hfff;
rom[16212] = 12'hfff;
rom[16213] = 12'hfff;
rom[16214] = 12'hfff;
rom[16215] = 12'hfff;
rom[16216] = 12'hfff;
rom[16217] = 12'hfff;
rom[16218] = 12'hfff;
rom[16219] = 12'hfff;
rom[16220] = 12'hfff;
rom[16221] = 12'hfff;
rom[16222] = 12'hfff;
rom[16223] = 12'hfff;
rom[16224] = 12'hfff;
rom[16225] = 12'hfff;
rom[16226] = 12'hfff;
rom[16227] = 12'hfff;
rom[16228] = 12'hfff;
rom[16229] = 12'hfff;
rom[16230] = 12'hfff;
rom[16231] = 12'hfff;
rom[16232] = 12'hfff;
rom[16233] = 12'hfff;
rom[16234] = 12'hfff;
rom[16235] = 12'hfff;
rom[16236] = 12'hfff;
rom[16237] = 12'hfff;
rom[16238] = 12'hfff;
rom[16239] = 12'hfff;
rom[16240] = 12'hfff;
rom[16241] = 12'hfff;
rom[16242] = 12'hfff;
rom[16243] = 12'hfff;
rom[16244] = 12'hfff;
rom[16245] = 12'hfff;
rom[16246] = 12'hfff;
rom[16247] = 12'hfff;
rom[16248] = 12'hfff;
rom[16249] = 12'hfff;
rom[16250] = 12'hfff;
rom[16251] = 12'hfff;
rom[16252] = 12'hfff;
rom[16253] = 12'hfff;
rom[16254] = 12'hfff;
rom[16255] = 12'hfff;
rom[16256] = 12'hfff;
rom[16257] = 12'hfff;
rom[16258] = 12'hfff;
rom[16259] = 12'hfff;
rom[16260] = 12'hfff;
rom[16261] = 12'hfff;
rom[16262] = 12'hfff;
rom[16263] = 12'hfff;
rom[16264] = 12'hfff;
rom[16265] = 12'hfff;
rom[16266] = 12'hfff;
rom[16267] = 12'hfff;
rom[16268] = 12'hfff;
rom[16269] = 12'hfff;
rom[16270] = 12'hfff;
rom[16271] = 12'hfff;
rom[16272] = 12'hfff;
rom[16273] = 12'hfff;
rom[16274] = 12'hfff;
rom[16275] = 12'hfff;
rom[16276] = 12'hfff;
rom[16277] = 12'hfff;
rom[16278] = 12'hfff;
rom[16279] = 12'hfff;
rom[16280] = 12'hfff;
rom[16281] = 12'hfff;
rom[16282] = 12'hfff;
rom[16283] = 12'hfff;
rom[16284] = 12'hfff;
rom[16285] = 12'hfff;
rom[16286] = 12'hfff;
rom[16287] = 12'hfff;
rom[16288] = 12'hfff;
rom[16289] = 12'hfff;
rom[16290] = 12'hfff;
rom[16291] = 12'hfff;
rom[16292] = 12'hfff;
rom[16293] = 12'hfff;
rom[16294] = 12'hfff;
rom[16295] = 12'hfff;
rom[16296] = 12'hfff;
rom[16297] = 12'hfff;
rom[16298] = 12'hfff;
rom[16299] = 12'hfff;
rom[16300] = 12'hfff;
rom[16301] = 12'hfff;
rom[16302] = 12'hfff;
rom[16303] = 12'hfff;
rom[16304] = 12'hfff;
rom[16305] = 12'hfff;
rom[16306] = 12'hfff;
rom[16307] = 12'hfff;
rom[16308] = 12'hfff;
rom[16309] = 12'hfff;
rom[16310] = 12'hfff;
rom[16311] = 12'hfff;
rom[16312] = 12'hfff;
rom[16313] = 12'hfff;
rom[16314] = 12'hfff;
rom[16315] = 12'hfff;
rom[16316] = 12'hfff;
rom[16317] = 12'hfff;
rom[16318] = 12'hfff;
rom[16319] = 12'hfff;
rom[16320] = 12'hfff;
rom[16321] = 12'hfff;
rom[16322] = 12'hfff;
rom[16323] = 12'hfff;
rom[16324] = 12'hfff;
rom[16325] = 12'hfff;
rom[16326] = 12'hfff;
rom[16327] = 12'hfff;
rom[16328] = 12'hfff;
rom[16329] = 12'hfff;
rom[16330] = 12'hfff;
rom[16331] = 12'hfff;
rom[16332] = 12'hfff;
rom[16333] = 12'hfff;
rom[16334] = 12'hfff;
rom[16335] = 12'hfff;
rom[16336] = 12'hfff;
rom[16337] = 12'hfff;
rom[16338] = 12'hfff;
rom[16339] = 12'hfff;
rom[16340] = 12'hfff;
rom[16341] = 12'hfff;
rom[16342] = 12'hfff;
rom[16343] = 12'hfff;
rom[16344] = 12'hfff;
rom[16345] = 12'hfff;
rom[16346] = 12'hfff;
rom[16347] = 12'hfff;
rom[16348] = 12'hfff;
rom[16349] = 12'hfff;
rom[16350] = 12'hfff;
rom[16351] = 12'hfff;
rom[16352] = 12'hfff;
rom[16353] = 12'hfff;
rom[16354] = 12'hfff;
rom[16355] = 12'hfff;
rom[16356] = 12'hfff;
rom[16357] = 12'hfff;
rom[16358] = 12'hfff;
rom[16359] = 12'hfff;
rom[16360] = 12'hfff;
rom[16361] = 12'hfff;
rom[16362] = 12'hfff;
rom[16363] = 12'hfff;
rom[16364] = 12'hfff;
rom[16365] = 12'hfff;
rom[16366] = 12'hfff;
rom[16367] = 12'hfff;
rom[16368] = 12'hfff;
rom[16369] = 12'hfff;
rom[16370] = 12'hfff;
rom[16371] = 12'hfff;
rom[16372] = 12'hfff;
rom[16373] = 12'hfff;
rom[16374] = 12'hfff;
rom[16375] = 12'hfff;
rom[16376] = 12'hfff;
rom[16377] = 12'hfff;
rom[16378] = 12'hfff;
rom[16379] = 12'hfff;
rom[16380] = 12'hfff;
rom[16381] = 12'hfff;
rom[16382] = 12'hfff;
rom[16383] = 12'hfff;
;end
endmodule
